`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
YyNmaNBFWFkoMr4+SC+IzSvEvuhU+08RTp6DmZab8WwCf2Itvs2IBd8QIIy2qq/EaCZSt5XDwA8+
wCS7I5qEWA==

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
FyhTuiXNspB6XnGauxASeTCNdgPX7G/s/XRKNQzKPhbVxDGHkZXEey2/R34AqKdASX6h2hOKACo+
fRCJ3LdJibtZ2X301AMleEGlLDc5L7dc0+7jPAdc4nxmshxo4MC5S/iqo55N5I8O7ROMvZUMVXG1
aPpyrzKzFx58EBiMtBY=

`protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
uUGQnnGhB4iDJ0s9LQfu/DBBT/StsiTG2arvDSUkKip73HY8HBXf01BdR5mlLLlRlcoXgfAuE5G3
rD01cFA2ouPF3Mmeredw7oQYoKrXUeQPdxnPie6MeR2XjIKHQAlofs3A53Jf2ecZIJ7Q/yZTtnco
um5aVRiRcfRwQy0Mecm5M9aEwZgjyj6RPtj39BeryW43MUOv4C/1XYpQtE8pkEOriTrpJLSE73de
ri14JMKE5fCds0kLelPZ3FJlPD62D/cYzvZ//qttIOIKdf+WXVQEg+JXNPo6/go3Sl5cfhvkIAq4
8Dh8Xk9acbmWep6pgCFVZQnGA7IXpuv2UdGj4g==

`protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
iLZZY8kP8FSLOFJCSj25Q6pbUXihEa/skxzaa/fEEnujOdFxf65O2nOGlI4UmFj9g52KRL+7sP4G
KaKiOpVC2BnHda3+d9bkRTQ/X3UXPGxsQFAsrpJwUeI4qjGm4KXt5DutGyZdKde89OjGm4fwaBCn
FbR+lUjB4X/SD4VxNbXEaFkC9x6wcSYocqNQ/S/t1QPowXE1URDFDkzw/k404LmOxG+2pVL2k2FU
mXziN9yaN3MOgJkoJOy3iWbN+5PVVRZJkBQ1FqQVRm6dTU3jcZTiYtVWEpnroQw87jYsWB3DAZwK
uq5JjK/mJ2v8SIlADi1OXJqzDFVVJqjdycxh8w==

`protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2019_02", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Z9DaMdD0zQtUHK0rq9bor6QHPoz+guzhftIcONOobwP/qIHkbtqb47bY3r9jv+BwMm/d+kZ9YP1O
jRNLbxYZzxtpouKLK0iI1vD89nQRoIXo6sbiAcFHwhi720rH0tNGcH6Iq9iIeRAw0o2GRWqgq/aC
9BRkKWm8okT/3DkutdGcD/pdBRUp3rRg2CBo3wtXQ9UeJNpq+SMMkP7PIu1cqRskY64p1zKcceH6
zYhavLqpXEL2dwsXNKhcyylG4U6PqLLfwPJcepkXa7rOlENkNCnwyL9ERbG/+90Me12Wk9+l7aSA
N0Bu69cN5FpLEOOffLrAtM7/NvmefWwGFyE8EA==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
ty9iuk6xp6f78B3IERkvNFAKzdw4/yzk5pAUCNVQizmj2JR/W5s5UWzZejCBkSEk3iGAbuu0petS
Tifz6lGdI6HYTvwnBHNketTyBKePrlHTvEtymeb3u90r1AuuvZBNyiMmFSw0585n4IuNJ5bmXMrA
XNmJ7cSntQphWVU1mO8=

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Z5VJ4fLO374Nt+T4JP3M0ARICFXixwpF1orTTQzmu0DwCEWJQ7eNx/pTp8bBbFj5ZhLks1DS06qh
s8o56ZWMF3h2G0RscYhDbeNVeK8e232mulQJdI0Y8ou9abYT7O6B5vk3hwA0zPSxUMipbgby7MSl
uec8iuO6O3YFPJ9/Nn6Vq/A6H3w8wgKMVybjUkl4RICiPnt/cOL/27UQDP7BKhJ+Vs0rqIjA798r
o77qdiOOcG3u2BV7mWNaJRLw4GO4dpt4xoBCa3x0g7GairuRc3rXBwbrDjg+0L/QkhjxyCyrpsGb
TKyep1pMdA1fEFSakOvwaDQ3RqWNery0K/ciew==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 1817168)
`protect data_block
+xcLu9trrMQ+ut75+ynM5mVWaW9TN+HvKW2x/pGdupMeuqSHPq2cy9RgWjLIbGmikieHJ74hdKVr
RU0DOG+LubRplbFI+2ZImdLnsNII3oDgGwAL5s4axR5Qhdmj5mVZRSxCPQJWFUNZG0YYxhBXAIcn
Bym5mPcEb9yyOA6yosOj6oJnUcpHk31SmNKx49tyncTbpKiXviEzh9dhbRvwOCoNWN36LKdlYwdL
mrrTmoca3dsT6e52jkZXFN5B8o3jT5GYrgf9MR16f1R5PlvGGEFPAxDDZb+jLCxXsBJGgqWsMrAe
TZW5kAEpHnKNuASPovibTHiXkgonO1iboZ9fqaJteP9VniCPKeqGTSHj+scyNJuDnrG++AAAXTaq
dICGofEeyP/T60gySGuu4wKzxEAq/CWVbJmnb1H+VsRJj+OLXy1qqvWfY69zWKA0H+OIFh3Qnzd4
y65FQ1USfX6FpyXSY3fDAiTCgENBgBR1744Ifz2QAGjbQIAMYA4uNDaf1eNuERuEbXgo+0mht4J4
JnZsxcobm6rHGwRd+FWfNxXt43INtdmTFHB/Od3u0aJWLnPcQEA++sr86i1LGSti/wWojFoZjzJj
DeCA7vUqKXuOiLu0x7bH+MDQ4Mt0pFdXYGOJYXJGzf+vSyHsUwNyyOiJtH2LMYv2rI3lJ54/NGIG
ubXLnnJZIqGXaVVVDe6xwraAuXrI7zy8spRt1E5m/ZMu9bmhjxNPSzrVyFktjwFrCD7o+9VGZURw
EDmq4TMATA0cmHhDtRYI52sISbN09l0ML0xGkXchERNA/JQEbndSqRlUsUZvtMX8WgfrWqaIm9wk
YNcafRAT6U1XhfWAwukMWrT88gx/c/vjOthLmIKNnCzNdaSpnh+AlS2xFRBMnVkR9jgaBzMMhg7V
5iVSR6IDToDZkWMtpxWs0EcLZLfyqhAH14Z6z0zsAfcTKgIZdSRJnsvQhPSQDBSFKb5g3xTdbE2P
AChvVhD1JCB1z7nrEF175Vnh2bq2CtkH+xJXn4LdXuWOE7FzEBrjd7F2fiIec/yEuSVNEhlgD+Dk
wJ2KT4/sTWBeEi3jnUnPXk7rlde6nWZPJ8X8X2HYs/THtpaXM/ME5PokiB76mHIC3ZZnEmDXYPy1
WKyUnipRc+r598xcqPTF2oqDXJWecCczVbaPXhH+NPRsqj+OVfj4uBF83Ojyt8X5t1BSUfFkDJhh
XdOSintljb2OxYjL8ny7psfRs5BWWf8sF+BXukFUgXgqOXkIHo8dIkrD/78I9t3uRRqn6TC9p1Sd
jw7KYpWf/X1SjDQC5dAYpKEIESnfPchVPZIL76gkwD5jnEDr4S16oxxfFiuSqaiA3asXw/w41hns
2E8FL7fwh3M9KaEnVWAp140FuCczjzkV1clOcVGgNCpjz5i7z7TBg8XtACNP3mlnsldrHuODw5yU
1pu6h64gXsuV1iWMZ2GfwDC+kg6nxkJR0PlKucPWMfKUZhzcFlGv0Zwa8iR+YZIx1HzpFpi7ni3A
86iNn+Q42xp9j8tlvCw4bZm37nJVht0sAu1oSsHglyfs3GC3VzDoBkYEEuGBvze3u3LHv1Vl806t
vr8w5f9SIW1ZgyZXPn8yT2aS5yA49VbDo2qb3b338iVGj4j+fkYCOCPRjzMbMfiQQDLHHTloIfiT
RwTGWgyf0vrgz7stCQIUj3KTm1fXKdJlPzMCWp5TQ+da4GQjv/GQcLvyi0lPCDvF9TTLVKEXLroB
QDu30/lFgQMjj/MTh/+Ix4Ea891oNiN2YgdPVFMZJ4bf29trzbTKXT6szLLOUzz6YtnsOjzDsVN8
mEiHyEG+wR+2HFcYtwLdeE/4obaodVxwbPx6tbMHdS1CNDoHb14+wQsz2Lw1C9e9Le9ph1OPcmdZ
/djwLEMJGjNZRZI872MuKkrF+pXPLJB24eHQSEiViGvbtsoBQHp26ZJ9aEv9Db1qeYep8seU66XP
N8kR3fgORHsGa5hz5kCN92ZlL1SszgDSODv6IX2Ts+zfNTidrfx+6mVRw5O1Rqy4oRLwAEwZCDw3
9Nlk4U0/Vqh3Jn1nlhAIrbpNG0i4eX3qEmlyUwvXgPUT7OxVvvMr0VDSnF9nG9i5o0JatoeajOxC
Mab5umzHUXaocwgRRzQChaz10ripAt8VFpNutKXKdyrYYoilHNzdIpFTpytClbV6UawP2ylkiX0u
nvZuRJjmoqGWhQpcE7cZlCJmti/9pM/wQ1eXXtuxPEC6d6k+wkjTK8xhsmDEdXMX1KhZEXLO1ehI
XBAfOkmZPH2n2G3jncdx4UEgV0GvcIs6XAznI942t0N7M8peMR48LUpUK3Gg21mZUPg5xJBUkGNo
dxClIFG+hpUtLLUu8MJsb8Oj3kVdvN47E2YMSlq1cfQjVGlnqGmZM2sLVJ35002CSuy+BnZHkN0Q
x7SaSqeKkXFg1r6E44nTAWJ54usTdFTMnTHab2Gz1H8s36oBXkZlbKwlkgdvatuRqt/4IWmodQ9K
taM1zDgZShGvzY2AbaXx8UtPBrIry6chmwqSzD4b8NpDAmqW+s1gc5GdU+V+Ka1zXBojDeBAx38f
fjVfvNR/87alaSkNVKTDioi8BUyzI8KiekMQK285OOdl7uMdiojIA6U22nX7JqZvSEH8UGRWl35C
Jm9vMucu5QRO/PiC68mI5bjQN+5Dwhv1weJGgCkMjcelKne+9Nr0G7fqQYSorxLlgq5AhTZyYm8m
g3bONDmNhqgrQ+S19vORMQBmIouyGWM4A+UglSxX0SZPoRouPlfPP3pgy5mtCnZ9AXfm9iFq+RxS
+dfIEl60qF5pwkq2dDX22G6rn0g62JdXR5FHoNr5QI82hUYHWWu79lFa6YekW9rNpy3Y9uAQV+R8
2KzFdYRIDycyY3pftlQNP6PGv4q1c6tW82FOPW9icucDLkE2tedjFGXk/ZW9w+sgR72bfR3iJ/OV
4tCSvG7cB8aJwfHI4XJJF3vljDLMIgi3Q6cFodfshb5Q0jQjmszei0ihVYO2/TOXa0JF/YXz7inR
CmGpo4tqkVHtgM6lVnqQ+eRBsC5ovgpExFSOQ3s7bZMxcX5UQxW4wb8infn0C2sIs/lbEhhGrqJ4
TCa09bNuX/nag4GwoJVzw/Q6ONYVUqIPucvpFOkVz++LuHlhKLkbJMe2E1LN4y7+1FuMpImOlVqE
6To5R42VtbqgQSsR9gpQaRuAQ7fIketRkjLKjsqxqvor1M9nflG8TFlhL1ZtShenCp5ljJ1+Wvln
61JQTxoIMi3FlSNqAGPDWEPMTxLBUljQ3m7Qr8avj+57UOwfO57NwllS7/9dm+QYOI23x+xnae4R
tfRO1z6vvmQV+1jt33ZwRJuY+uF2nB7lz/EW8qoM7ZwF6K3oJqU4SiljVgonh1UMLYYaQS7PEzi+
TGoGTBCDUgqr9pXnjlmL2TXYM6gwxDM7UA3iu0DNyyKqdX5Mi0GvQiYj+cpSdpBuBf9ieAPCJ/Yr
b0u1SqkMQ1MRSdzJe4pAjo2KFmdjVx+2/XtEucswkLXvKLnp6joupuuMBvVjpvmL/N8RFWsau0xJ
SmbDBgS5CZCtRpxEkyS0SE+zACYL1Fnq7YDisyuT1F+q8OVs9tLKMf8OEPMQlBV/ahWigmm6jshv
6Pt9Ki5mYKb064PKbLPlmU42THFQ08GqGSWtdPiipn+JeN7Zo22A7icROgiUbKuUI+gPsujovRTe
AsHcxqa9evwWxuGsk6P+eiNbdm23yaprtl0lk0maMLioIPsqmk2cUGjw3i0G20eU0hUDpmffzYsd
TjTWKR1GU9Ko+0WuQ4JpRf5lLQ1+h7GMh2czPEE2jHiyQNHmxcr7bl94KYyc0EaLKLO/TfXON9e1
7gZCp/M19aDvNeyXgTVk+bDtUqlUmmoY6quX/ZDCkLoHdH3h3kj5Shr2z/Jd9ZrVPvCxXwU1/+KS
WY01z43+QlFtw96yxPMSb2fVAbhKoYCQY4sq531TDl1/QHg8lsnOMGvl3CnlSc8hBkIqmnEqFn8P
BLlwBo/dGhRkfg8iKunmwp6+uc8XXNF0WynddQuMHhqL0+/HlYV7gmNU7qXk81oRs9uzclC0qhcK
BeB3HR1nAsnexicxV3IPKHQC/DN4HATWh8Pshp0dxnpAO9B7mQowive2iPtaG5yBkSlOCcug26K0
E1YmNpq4cq3Orsx/eJwqfj606LJ07W2yHsqwhkdlcvntLHE2Vrt4qTRGEFX3m+rGaphQUxvnhpZB
uHB6wa54+LB2AdihSBylWNdC2G2zsII1f19xEcNEW3fCF9jZ61o/HKEW4GWzqh0imj0QLjN6N64Y
O+/r9zRKA+rv1702Gcsi3B6lDRAyW8+WlSrHf9ZsLK9U8tUvHj1PLIMhFagwFhZ0ukMiVUNaaFTr
RZIRCYyGJHMn5GPHvJkhVH5+ArOVpb8efLqCVq5sm2C/DFceOmOFbdrMhEyS+/F0wp1iy1UiqUFj
0i4PBEpkj6aVGyqi4V21uyHHs2M9k+DDoGz4D4MzOXKxU6C+GI/uQK4fexYrOzRrebtnwPOtq65m
7oEsXSTN5YRCIt0wQWXsnug8JDD4Ud1Ut+mtdyJRfhGoj/zQkdkJ5rra1mxknBUzFF3c5QlGX0t0
8/tL7YQ4co89uZjVw2NB3gp9kzVMOb+sreKsvnHU3i1byYiQW2oePeZiN53b7mzuUjq7Z9oXD1ed
mPY43loNEU1vXg+AlPuONoOtNImnUxJMeNrmFsTVjK66BGdWAvyAniXVZalRnsi2mVP2FNYCL7B9
BOJ7Ow9z0hL3WJgjFr4P3AYy4mRGH5Ow3asJBb1i0TP3zGpscDFLiCBZzN+w8EJvIi2C4bSxfK2n
1lugBJNSpNqlsTK4hDo3UUYfsBcUVkr6chdNmkWmBUcb9T7OxgxST8mQSNESKt8dP8O3VrhKxrkr
qxfgD3/gG4N1efB/6Zp0wO3XZguLLmd56WREYVuGWMqu0iqmQx+fsF7FQ+FBMkLw5P5mhf94j6AS
EQ6LWRxD1XXU9IzyficQWlbcKA+ineOPiOYaXy+9R0PNE8eriSMSz3RBhYF3VOtjYBTZ8NsMoyG5
wS0mkUICU2k9mphNdhOuDyA2gDHY+JhT9/1WiwPhmvTasfUFsd8n56awD3eH2yECeS8+Onj7n9b5
26aa2vLUrVG6Tq79ajzyJIN0rjeRee9748i5sGXj/EAyKVTAA5QIToJs9ER0jFunvMT2qloijmuM
kANRz/1aYw/jqiLD4E7DZW4sjO8PCLJHNfO4loKub527UCe6Di9QoQC/OEL/FYXTxTviLPpSAMwI
G9do0GUU5rgC00z4yLhiI1PV42whyNPFVdiQrXBzPbFdBpoPkdmwa3qxzTiXLpfTL8PDsc1N+9xy
XdY0roW91RkHYj/Acg8HsTaKxwNoU1rndyDBQiJGbQz4ryjP2G7D0R2SbebWBEW3gS55c1/kwpod
1q1gQ2iIvTc0KuXrsKP+HjzdTmNE+ZC1MfiZ56Z1Jf5xYwgk0JQCmWzCcmByC77lGj745j8KYWZA
qCOvd0EnCmSfWQZJDihhSxc7FlD996VqcqC0AKY0fnoVm0iuRPSS9x2m6MNLCI9/JzT9U7TbzaHW
GHUNM7djveohJnO8bimWZ/52oko90E9hCHzSOvunEdhlxZZRP07VAeOHvmcEBEytpApeAuTgKOil
ctra/WJkRtImuh1/T/SVERyj9M02yS1gMeEthUJN8Le24Lv/sNth308SWVHeG+lijRrhXwAw38Cl
ySKJ5jCTdY7WMjynFo6JAleRza2iPFrgp0mbt5u+C9qK/GXu4kxrb5s59sUOFSvJ484sOGVl/+/i
Qqaa4dT6YaeGZ00jsSWAczCxRQ7nJvmbuRRkwNh71IPjaUn7Aunlh8i/QzjN4hECw8PWpI/LL5BB
JDH99SgeToArxfLi2K75RX8EvlnQ3GnrMc1JWPKrHcxkS2REB0+KgJY/pZ0BDLgM5TpDTx0pF3Zk
Or4sGuiZPIn3JZv0WqbS0kZniRYbynCbwfkeiaQjTDFUNsj+EgcCr/U1GhaNnvjNjVCZbc9fwvnr
ugcQnPqZhvCmYSgaPjNdPTBfK6YrXysR5s3P8wjqa5T7powlnIA4mIpMhyAJCjGfuUDzRAaSBkWp
65wytZwsoM/Uy9cyeN7znAzwmZS8mz4nbu+1K1+0OwgMXlNQOXXoWu1SMgYQMheYM4Wi/QA2yKSQ
ak+yLTqHqvhFy8rB8DGY+odmfJq3IgKuKMUalCPvLGXeeauQXm+gHMfPcWyvAdSAIJWmWbzG20Ra
l8rQ8umDNaPpgpusB3jurDfcI+B2IqIiC/AEecR8sWu2Az5DsTOfJ6v+xRfeUAFZidrYg3HM2GKJ
2uOc6DHtCL7+I6aUMOHTYryWzo1ySx18V9NpFJUh2I+qHELGAmsmY9iHq+D8bYim6EOvIhQz58Oy
AhHtXWFAS9LNvvZOhr/Sj6I3X+gwT0xmQSokuN8b+DBK4x1jaaewHzgenEdFIUoMaFDiehnGZNWa
olpJjR6q3w8nANEjfcAsBJ9+xIZPdEnjlh6DE7LBFDTCv9h7a2PDF/9ValvyUCo04UtrettEzmYK
hBIgRXKCsIvf1RT7qWEii8N13SSBJHikZykdhMq5N+U2RcbiosaLOgDrIe/OpmQF9aeptmsYx0zD
e1Vsgyf3kovYAei65WV1UgVSk/Y1fp2hKKBjU2D8ofpUEruaUAsF/j7G6gts78sgXa4aTs4sU+rl
iD8hRBM45GRuAOiP1G7VLNF4mheHWBO8lOGbYdzlFJtheSL58jXjia3uD1vDKQDfwcYZvBWYmTvn
eIvCkTDZdQn1iLz3wzx4zC/ZwaN5dqLome9nLpqUlCdBc1LZEsx+RtJYu52VFTQ8jOLhTxFIFT2X
hmMOrHDQfx6CIHA/h6yln2f8NehjmpuUcIEju9PWSjVa6JtQa9RkebtG1GtwqKsLWF7Eh2M20pAA
jAMVG7z/z+Hon3ELsXbIZ9v1iri8OObfWAswRYwgEcSrVI1vuadMs37zLeZbdPJqaXilYLlKMng6
wNFk3gm0y7r2c+H4CAcuFye2pGxHPJJ174CCvl0VYZlfUITQxA3H+L5kNvkgFIv2VCY06S5YRWUE
F1EdNG7R+pARJLHNk59zOwfiVYBhZFF1D0xNaBzz3PP8s8ZUvMkSHCDLvUtGyqo097fWQDsmyTJY
/aFQybMvT7i+NaG5w0IwTWvQw16p3O2X02cjzwon0l0lcFuI8FGrOv2beksowFQElhUbYfi7AFG+
yjKu88duI6suU9sktl2yvPGeO8+7EdItOhtUdTJOI2+FB3ApiwtRTxy/CFAtzyRSAq/0SDk3OJ+y
H+V6fxHIAGG1H6Ou3INIBB+8xwxx3qCE0OF8mEG1k953+h5S9OK0ZV1dhB58t6n0mvjCAW01bkyO
WyUhLj8Z8X5CickMGg1N7v1H4tV8OB9i7ww5cWrHXbxggrAR9NRP+po82qhTKl9liZpqnp081u8D
xdBVUpBcp8EpecNaFN6JpJ6txSbeyyEW9dPwQxyjEZ+Y46R7nyPb69vclbqeE+avqbrqRrpj/Bpe
tvhGsK53y0YjgEVmir4FEEzVjALNGxtWtAdvpZXbdyKqzJ+d3u4gbR9++YxCnaHRJ9G+6ZN1dty2
qmDCacTRi8LcrE6I6g++1LQMADD6FGBbizFvgyabthFnIOWohdAW83k2cp0CGWkYRIcWvkkzVqM1
s+QUt1EzOspfkEorkJS9H1lHssRjrjsBxMvdEa57DW8tb0VkNtJWhb1bPNKjP0CoAvDNLObyIlgs
TFzlSL6M98uOdRc1mU9XhoRftZyg9/cZPsp9ekK6enfVBWOR9BLZnHMiAeEFz8dObxTwmmm/QMJV
t5fwg42qQHznMMCnKo6Vb58EByNXphVIZgVtHjpav0lJc6AypAE+3GujVB+xlxfHhXgPUh11y0YH
jz7htS6Q2Y/Twf0NzFDDt1QcemZf181VVuPgXeVuFTbo90fvKWyjsjRInL0A4r0n5EBJtqo9Itbu
IPjNjofaX2BZRiV57FKkPB5XT7VZX92SdqskINe8Sic4chE4ehxl3oF9a72aqVCmMz/aKOGOylYF
TKuMrxNBUzYzUpVdeti/bV/CeZMpMtckSaynpaQl8tPunQAYVxU0HLWXAY15OstWLNYkSU/13hlW
wEeAsCyrEUQrED7wadePpemH+VX/okyd87vEc89QI9nE4pg5Louy2R9sxBxbtkvd86dbl0LjNsWm
G46LeiNmAQvWZ7IJaS27/5AQuMmgxAAFw8ylwWtsH6Hzh3CRJXFzYrG58/6M12QyyydQgwlas1im
/cEKImXnS/TvoH8O6uX3l/DQOzExhDlrPAElVpHwoSnyr5XNK1gt6A+RaZ/AwfUhGzDHezU/w+MZ
ms8m1aj+ig0OHW3MRVfQar3hdm3b6PBZ0a0ftzWvBtSkY66Nu1E2yzB6uQuirQyjJ7IQ83FRSMVx
QR5uPf5BKgQoXIAVylBHd9zYrqk97ogMBpBAHim5PpHPdzFmH6Aruviu+yOtsCewTfxpO/urYS5y
WTLaj0c6GRGhppZ0zFxul3NqoetXMfxViC6uAHeqqWzhomlCBwq5srL40A421lVdh1HkIJ1HMYVW
my1DgxbY5Qzbw4Ol+h47OOL6v8o07ZoBAWSdgJqkauWQpvpp2TDgil32k7hcVK7VLXtmZkQv7pQT
G6tiCtIGGDiuGVPVVIcEejS3qYa/7i1lMLdWzWWlIsqqPHYDRn/4BDJ0dZ39ScyamrmiEP5iOuF9
/yux8gqnOmu/mujVmAzg32kKppBi9kVqc8EOlzYFzvVChGASLsy1iA7uqve674yf+0OY222ru9fP
+JjhenrRhgDDTacqcaJSk0+cHRfvUYYzzqDr+oga6li49LE2uJMu8RIUub+oItcUnGmgfzFxB130
T9kCuAWfFrTvyyUS5NZHVorD1V/slqbIoVfGax+fVGMA5XaaS/c/XnrfckOif/OCDWNcVEaJKNqF
yqM9ZMRYEAmXdQrq+0RzDa86zOq+5SaH2kXVRqnHm1/H1MncLMDhLTBv4MtMnV6kqeAysjpuVaxR
n11q+ohv1QGujawkzFcE2KUQqlUxNKqaXc4c1qAnZ66dM7ZHxIeQlazjBEk8lIMU6ZmZPlij2era
R8Xcjuk6Xr+jWhjSjurzlHCPaXhfw5s22+Vs28a23uCfghslAnn2FDab0ILx5jIM4LtaapyRQVy8
RuHfl/xQLbmKwe9B4jlCfsDgt0b2+ZWcCroimeh9BH6CP5sBmGRmwdRAE7GT5zBU7eSEKOCNr8QB
LR37LLbzwrztlGxHn76wZ7K2/D2WgLkRdYLCK4t28g6zY1GoGscsPF22A7TC+88ZO8dtn5VXYme+
EiNwZwwHTXIaeJ+UyN6xsanWk2d40vM6wFNWycxEFVuMmtSmM8TkYGBnOaT3IkY+pFzH+3Jn+3qw
1m1L/ZcLr/VQ5ccyxoAiwkXZ6u50KQ333O8xWJM+sZ+SER5MrCplyr7xdJKubh5rJBtzDZvq07Ae
Ad1a1o6qSVUqyRrtAm3+iWbtllYDw04Rv2myIKftrpTCshSBeDal79SyMeyV7eQLwoJkw0v/f6oq
0km189+PfNra/l0Oj7XCvOvdU366zRibfWKLsDDFnrp1sQDzUQvJH+Kn9dl3BiP+S9A0jhsxWRAs
ZfRJsWw+38JpMVu95WM/Z/yXzHY8HvtlTZMUnv+jijbK/h7lNEzNNoYQgdLF4q+vUOVLIkFXwbhj
AgjYCgrF18WSBWpbH2AgoKMhjXV4acvZ+Ak+uJ1qqkSiI2Y93zNHzOYBJ/l75UXpne21xiwH1lcp
1iSPWfJDv+68Oj0j0+X9GMW70zOYDEPzjpnZ8w70gh9uPbUBbgRTzJzAguDQluLuQljoFHkNY0BV
WQfEMHeHEcR65uJnt5D0zr4tCeIlDEQWFpK3F8jgIk9PBnFuKvMJBKTQ+F2ZxDG0WNCXTQy50ITh
KgjLOIrtHEBPmwvcl9KtWYlTkCnB0neoCrMhvv5EyPhd9CWlCc7My89BFpNxwUi2S5eY9nSFWzvH
2nB1V1+folRNZtlp7tYWlzaNNY57Lq8qbaBmtrWAUqCIySqmoALqnrstQRDGDvR77hMFCBsad4rD
RCpkQam/S/cvKGlEb4FzpANUDg9aJzc1KdV5IKMJMDU7sVlg0fjPhQzSAYcO4yg4X3n1MwV2TbdH
XfJ2Co2cwMtQK0r4WfDnYFwPk9fMp1G3k03WyMd/VOt460G5mnVxLdMM4A8deKAGOCNvc6R51pF/
gARAGI+kenW5jGbBvE4CJIDU8Pc5SgLUHRY5GZe0/AarLWx88D/ozktIgo983CaoF4v28dFCuRlS
R5XzKYJn60mI+cakQBKMlDTYBrDIOATEaxUDkJNrNRwV/JuXnG7jMtHrOX8xYQV/dQppGRLdaxDZ
nj0hdeUhy3eL0Ssv+6JWg4uOA94DOGpvga7c4NLm+WUsf76zSPyNtJYXMIh8yHss3Xn2FqsyhJBD
ucPOluWecm25yxn7EJSn2FMw1QsLobIRel1mbJeJvrv4sRriR+cTD9nGEM10Y21B8gcm8OyIcGYY
8C3nhCBgW5bGC8duCz2VV0/x59Tle1Ts7WqYFYlt2EcIEgGUU6gOYEDkgbz/Eu8v2R24qcYU5Tci
cuaV7NauWfd3vnA5Ukboe93pLOBbwzd9y48M//t1+OsAZ+4+u6p97ku1nRUC7xqjM7jWAuINEck8
AuvixgUbk0riCxPfJ8+11TnRs/e7NJ4NAWdlZeQ5GMmfo3gSTMEdMvUY4yJFB6lLyfDA9H2bsm7B
FldP5eqJk3/YK3oI49bMx8f3N2dgZ1k5PhpwSI5eoegzd4BW7eVdwQ6XVjtMCUOJUEBL74u28op/
e+m5fJfCiyLGSaIqGIb0f5H3+xThJXYTBrbBS601pSTxBfYCNpYkcIiQTl7/vKwXnDFTnL15zYSM
wcNGJkcPoU08+BN0x/L0HEDL6w1X2H3g5tvraa3cARZGe8YcR/+F07z0FuYVK3Tjf35WjWaV+p/9
0OgZup/wtgtXphzze6Dhocjx0XALkzqDA5oiLXA/aHVbP8mAPhCzvO4LnXzWkHn+ZMUOHTUGQv64
VndUJe5UjD7r8RIQSx1UwmG1oi3YFJQMujWQc31f7xfiankg8rAK218tXB33B4Co6NhaobhU6Kbb
q5Gq/LoomVEfPR5DGS5xtIa8M0duSttbMfX+Z0m682tO89waM2N2xtHCEIvrDxFjpa4QU+kXl4dx
5+dGu9UaHTjPVbcK9KLtVP7iD/4G2X391Xg7NLlTCWtm5y3CaUwfSS96dYt2Nl3btnWp65ExEWuH
/H89nXna0ygU4fDnzYzqx75746C5p9hzcxF2810xUOrPf9mFY9y908+qnzptTIy3mL2+ywrUSI9q
GYKcPcmTqWsLBrZB16ck3L75O63Jk8SRMegdhE9In+TeM5meUf6sN2JkLID9HNapX8kCkOR+UA5z
llBDpE9pKSWsB2TciUi5C5mGJlkW1YB2VNkv4s/2ffq9pmsOe0HHHZfjIfctdncFM5lqZrLzWQJv
pyFBCy3xNZjFWTREKtr7H6kPlsihd1S0aZOyK7ATfzXyjnXmzWit5kzCUIaFaRxsPohfvp0g/3fU
HspBfPcsDPrAGnCTfGTxtuolUTK7QNCMiLtuGT8yWcfLK1m8s7X7GckDLJymgMV7+fhSxiSG7cXX
Tm+wEw6gw+QmNVj4iiMEJc5mAvR0P2+Nj0I1tgpseUIVikTuNrJxbP4g85DGh3JCH/Qavvq0pj9I
Xd4hfHpdFaJn9jhKmN8KikjmSWy2cTrjhvf4VeuVdvy2DCNDkqF+5i2bFnXF0Oh2OtmV+ufJ8lDE
Vw0j2tOjujeqw9rGHk8fff7Eaimsx7INvYwxN4jZogcr2FfdYThBO4JZXIL3RzXN7DzTo3OIgvN7
XVAHPlCS9nY4tm99C7nPXWDiVWzlxuZXdh+pHae/ke1eSlS/O4N4QAc1vkRXJGqTOD0Dbvf7Ic29
63SQaWoun3XiXFOr4SVGJ+To8iJdcady/dQgq7A76cvd7/ZKNujqSGUean5g0E9KiSP61HbzA2Ew
jVcyWqOyf0wWnfVQZQ9R1UF4levPj1wR1B7eBj0GXEWK49OAN9M6X01UQp2B+Y0ePX4FfZ+1PZ3F
JtJwJDH2/Bnq0cZdcEYVVnXoDIIv4ofl/8QFWTzoo7SjUKTVySdpfa5WGyr54dkhNWdHn+sESSyL
DLORUzs0+vSAlEJY+nhiaeTHtVXsDiPq34aaWXgqcHLv8w60ZXG+btSNUjo9s9ofV/pUDKehvAus
LptbLTLzi8+BPFUQ6YUdYecDVilqVX6upnPc5nswSuXud8h3XWboCzwodZpFpKsnrtAP4gMzCVeN
wdRWurJlvMtturuHKC06k8dFQJxW8O6N/bkCCCX7VnuzWUrO71FcF4K+YTNNqmb/QAXLwV1wViKP
A1QCcrQI9u9T33iZu/aoJ3xBZrZLGX28YlETAGf6FMg3EsUwcjEsDmjRGxRlcsvZaIiPCVZPvhYi
ZFNzE5jWliwP+Z7Wd74g2CRnQGhbIJpCkjuR4mAtR5f73yadx7CPAWB8s+P/zKuiYF5nk68lIEm+
eqifmmXR6DIetl1oTwUION+bOxlAXqfkwnCOuCAXleNrPmPbenp6hfidID/8KpwHxruyQu4Q3ddI
0F3FpKMIem2d5AcPA6lGue/JavZws/D00GACrT+GEWiyXzV72LKjS/lj0wO8cgtTkEF15YVclxVt
xt75R+sjm8TcOxZAVQvSNgK56ses3z9eXw+DoKr7D8EIxjTY6I8O1RP6oq42vcIqiBePoJ3muS/W
gnol5vL1stPjQcn91iWn1rQcBhgtlDgQkeD0Ozrn1fubiAEohUnaCXggSVB721NNG6OHonFBvRfr
1NE8mtDeIr0e1NSzKMD72iUlWKRSH51tYKDYwZWP34tvPhwpQds2Pr7Fj9QGXMTLey+VSyODlBJX
KaSlKQocQHO0f6zbw7Dwq5l1u5QwiyW9CIzSUqL7LuXuq1xNnE8lxk4ZgoF3cFwbwRIqCIGW5Jno
JVQF91cyIJGbBJU+mZmD7WAgPDxpeTByW8+mNJMq9AFLL+K7m66dZzyL8whUuS7QsFWVbm5PunDR
bWV/biGZmynnOQVEVIbOUQzsPB0bsfDIdptnXS1+RJ3C98yA48NmPQEJzp1KstatMN3FCqRlBZ0Q
9HYWiq0o/w3KDsLD4s7VwGW40dk7h64YYFniSB5wcQAuLOKHcdvupRjMC6Ab2UqNsvUHl4CSOLj/
o9VNfEpNXzUaMsuGvgXunpjlZTAhNzeKOP6KgnOy/wkqKqa8meh7OTtYssmJqr3xFwqr7NWqUO+K
cW1pPe+jlqqZZIgEL913MUFoGLW/eApSMdirYANKany+V0M0Ac9MKg6oxb1tcNzptlto3OzsU1P5
ciNXMZJMaPLBmaLRml01dCxOtRj1c62NnFt4zg+AI2bM8AyVceyy7S/hDqhQa2Ub43a0XHY5VafD
BOdO5s2BUxpOU+PLPrNXTmLvers08sNYlyLzUi0oqxpjNVPcnmBQFUrpfbI6pbQChzrRdFcz20os
bp9kXbaYyYJjCFGRB+G7K2XOoNjk9/9z3Un/K0qEFSLD6gFQxvL3hFEAFdtBLUp4BzdqM9Q4jS1A
pXqRXJnErx5VqJfCj8HQc/mbtpDY8Rp6gTOmB4FeYuE8oUeErmKC8m5HW68lmSyCwYdNvcpFLcFt
kOGxr56dZT+cybn0WJt3qHmkMBx0C9o46fFGIDP/SlTyZM8tJxBtguY/9/RNIaRJ+SlLrPSnkCMa
KmTF2Lc+XcRLly6X+jITpMfvrcQ2oDc8CvhAkAHXjaFBRHgiFw4s0+/eQEE5rJJ2JesIIGKGJDHW
iLilSFuL3QOoRioo21sq0qqDOfJ85ArB5ibbdbuD9qWw4wNqCVHq7r1RQYD5d1IXfMI+Dazu1IA7
ol1Mo2ypLd7YZCLteC22GPDQf7S5/Wb00RFM58XIyFLq2FgnUWYzcUO2b91vqGklbV6cSLWAW00u
IRbXQ8nlyaOXwKVm65UBf5YeGrIqfe24i5eKg++VkhPlEca0qbL+au5TsXdrpajD6iL2DlI0Cw3r
rsxdaWbo21aYccklVKSZszspAho9dPUA0IXfV1mZ3P7vwX07AErQCpaB+BwLnUs3t9CNeimeyzIW
RKQloaftsSZOtWCD4YsVNst1nl2rxFEiT93HlNupfT9+TUHVNh8d/lgNH9x0hpvuvvSLFbRSq0sm
ctM1RgEHH5tVfBfHp1LPx9FyMidoF6Ovgva1msRvCcPUAw6BpExjinuOW8xAL9rLFEHq1v7FuUuH
767cfbPrR1/ONyzZ1nHmFIZt0ayGd9jnQvaIaVQZttADNjxIkbeYIYYKmaFZLA/9FMow853A6nk7
C8tJ+Ywoy9iKmNJaPpvKUOz2XYRsm/sPlZexZm1J2oTjfdkQltWBR1mSsPKtRibx0ttKYRWjkBOH
tbyyimSPHYTG+l5kh/95GBrZ4pfJ65cmq6UQgpg19X9SATcNrDLgB2cE0/VodfrsQLVVQMjRlA6k
LQ/1voVi32Q5QipcmUoZGQw03Dm6Ro1aF42A/opBmbBmdEhjp4ol6jKuaujpVFYoZnA3Yexlpk/r
JXgpTnRDeudB2hXRoxB+DnWxNaorodAQ6PilUndtEuPu8nj/PqHOIxNERGTugqodR5Bt4cTAwQXd
CmYb4zEcRgiemc3lOKYecNQ7UKDGwK11CKU8U6AcvrLkUjyaOFmXLzS1s0oYQlzfm/2PiXphJ//J
4qlkJEGD/w2r8VRio/vZ6ZEey/kYCqecjJFuvKzPrcpu6EzysJp1MA/6Ll1FzZop9SvXknL4fUQN
12E3TM6TWW8L1yCiccl/8kf6Dj4hJgapasLKQAA3NsZ1rkArtyFM3zF3LYXCppLCRZuYOc2XKdXc
gRH3vXN2ozwsAKoNNzHFxf3odPbLDz+146U+Q5+VLYigZtIQCuWk3WXYawG/JgacWc/BEPPC2jJj
8I8bTYyTKlta43vBr/m9GcLIWTiajoSENGwsodtHzqK9F5liz/8SnUIa7U09d0liRmzDmqp/hsf0
W7mNbCH093xGyCT80rebAH7txS9vGwKVLCnsB4UhsctWMVZUMa8kpb8jcnySpKGPaDc82aLy3mKx
LWOsLgo4lgwh173lwHvpD70isYxfpVFpM3Q0QjRX8fkCkOAuavYXJLFqaqe+fLDqykcNe6FOJBx0
zAvSmgQPtOrnYTU7DRU7PA4xtnhq3Pivk76rB6PmxsdgwtLrKus3/UqY9fzZXktZtCaXavTiiuNS
lhRjhwPPFwjJex6Tfy0MRVcQHe/L0BNJX5WP2m8zAgsQUMRmk4LrJ+E4vJgguUuM9B3ivU1KTnFE
Ukg8nn/Aks66KQY++lJURZxzmt5K8GDZ5J761hV42fIcMiH+nrhOUjzcDK8SbjV/bHtFV3Je5KTo
zNa/jxRUNabXU/yf0DUQiy4rLZWe73dyhXZmvrGOx3rYW0NxKXZvo9oqq1FSftvFuclJqsX4aa2v
eHViI8K91UwuL42qxfSQssaslNWj/4x2fWMrzowsfXGWwNJ7/CkU+0gDagpx0W7bXI5mlmCM70rh
DRwT7GFUgJm1d+krXfDkJh46PPJOk9z5ysMb08alCizBTHX8RA7zAUdNkBXMkSu+Mff/b2bGiNpa
V6uVTkNbnRGu+7J+dY7LkkOrEgsCQMHUdLRGmAzyADeF8r/5exoArYhWZqX0E4MCVymA/7pYcBky
NWH13yX35KnI+XHrCH1QqXmy8HlCVZBT8otxOPuq/IC8xi7FFFDOPSpQ8ZhS5acJl/SfcLXMfnmd
4namu/Ph1nFYRx3m4EMcpPKZFQcPx9T5AW6E8PI5WmnSnfymeadjR9My0r5XB53TRvqinQz5WKKf
CB67iDdwBycCcpkDP/nIativYEDVEFE7TPFvRbq/ubkWe5tcJhueB9eLUtoAmVg0OunE7mllU84F
5jl3sspeA8j47vFdYyYEOVm4rwUHaw7pJtgzLJedLc9AGUFLTO5QBN6lYjw4D3aFG3kh/o5bP1tc
Yh04ZRi8J/nNkjXZYalWzmzGseWrhdfGBlL+sgIzrCZidTLXQrNfa/AT44Qm5n3l49M/lbgWSGcZ
n53uyxA0z2EqbYzLPDFuf0rgna+TDcIu7d0lPwMru/ryifMUx6EgZoy8gP0Kbmxq9hf+97PXxf2J
VG17ulXPgIp+r2jbl0Vvux19CccabrlVo72MneZU+Hktjkr7uieE0OwK9JyURSmyZyzMs3/Bm+Hl
ssawAJYu/ZP9k7jGX/HK3N6yfiOGDYIwvJetr5uhapNsWlEQbeycLQeQJ21Ab2m43j1/R2n2C7LA
84mfWszqBFwDDaSBoN1VHnUHMQLVxitF/FtaVdiA1ivaaB8x3Wb9Gfzr6g+/Jo5epk8038y/Ddd1
EiQcD1FQoaPtFOZVZL/DNB9g0zN5Iz+tx+Ael752oDH7tm76qk97+NAYnLSe9lYgUWc03TWKa7hJ
HS0cCPtrhOF8ymtIUXOsiMtZYHwba98dkeRGPNrgakvPvxkHZhUmNOBzJnVzapmbNCd7pX5E91s9
7cYlkFBXEVmGzuHSdb/q8Ml5rsRz7+B6f3zKj1kBwGwMRv8CR7bT2I44hF9CiM1ABsq3gEOxqnjY
7dk1bdBlUpl7t6b0nT/KjkuwHP0DWqdrTMwF3JBuccD7AKNpzjTnKpvOXP3pVGO/gtgOIRpu1ag4
sAeyALqBXFbOeMU5rOyp0sEL6ivXCIt/xQemUz+cg3oNksUo4HFJeoq3RhY9bG4qWDhE6OeJcm7Y
cH++M1u0xpnoLb9If9pVbgmlNYX/PNU7IgNSvc4bBZedP4O6mLHCOgrtl7yCqciSfQ/QJfn/25yq
/JdZSWqL++1HlAYTXKr7rEcdeim41cjVzRP3Qtl9qDvE0IWWs1mR25yIj8w8ZgS2VoDwjD1HW2RE
iuOeDCh0CV7MNpDV2BzkXhHg5h+k68CHvX/p7vdK9nt1+HxNkoJHJCx7KaHqPx4mEbSIblvNt9PZ
DNFh2yYMi8SdvJdVjeqBqFcXaaS+67qHr/9mIRGNagRDqUzQd+RRV5xGXWshhjM6CjHj/XrWaHWc
Z9hW74Fjq7rHKqwqVnoymdRkAT3JL5fK9uPmdt7pHEQu5GyRn6sJwKOPdiWSO+JTG4ERxIgzHcZ8
H1oZ+sX3f35gnIZIKzU8F18jraVCYVNnC18l/99slG+9TscOKyejFNl4IPJZ5Ioq0VdPwexOa0oG
2EG/xqW34pmfMEyS5SmAUnT1p+Ki4uN6jHQib0LTDE+nrq57oseIm1It9DZ1CNV4rMRlweKANnRG
VThYYWNgsnJyGYMEK+3/NWFhICL/+kjiNIW1IsfcrVwBgILBpxdJV3uQTU0uveT48367yzuD76us
V+O2gQg2KR8pNbxIHQ9VdHXIJeOTFhkGQMgVQ+yfkAao5WH7ctbeTTS/23IRaIh+wz9FvstrMbmV
VqHh03wsRzBSIsS96fdqv1wZdXfBrEbqGwjMy0M4XdDQ6WbcX2FokMRVHUr6iiwUYv7reRc7Wjo0
vNzObL1nbuJ6tkWhhDahBx2iGTuzk0BFDpe3qU9mYxJX9A1xVtbtkuRmblcWuAu09d02na0rOqtq
KFlkPZBR80Y7Pl5KhZ331Q8frB3lC6pyfeHgjLWDIKGoeit2GdM3jMDR+1eZm/alpJImoBc2a/fy
Xnfcvo4vj+fallhGBrlbTJUBVoZJDQd9PXT5iIx69CJQ0iCNu5ShzgLtxv6MdQjnveP7Vrboq+Eu
z3WSTNCyAaHib8zwqaD75Ud9/0PrmmbTLBGUK6SaNGL2kQnMfoRnsNDQat2kgus4e1Xkac5LyV9P
FuCVxctWb23/cfgh2R2QwqNu9C/cNSJVb54tfqZCE28t+km+ag9JmPLFVYyWP7EVv+y34wvwcNTW
aWIFaAsL69MQ1fYn8nU9yooXBm5anHuOAjeOPtpwWvvTdHtPqDM5C4huQ3FyJTuISAD7CcbsY2Sr
SyqV/BlVHsQOTHNu1zsUxEWOf1v5CqXvxl8TUILH6LCXpqAUpD76TxZLzc9YXISttmnqueR0y6aF
b14zhza7w4LXrF/sPYQmteZWZhMSgSjvYZiemSliiBkwB5QHIIdIliroPmO28VU53VmhihweTBBK
f3rhup3xkNB5RBjEGwbUohTdKpA8HJ2nv72Ic/hzS/DWYIJ+ZIxqVzAftZ6rnUbInCC5NdCjCPoM
KR9bar2Lznep7Yp0tiO7gq2XxokqiGQarvPA/XKGDX1o9jQ1lxrue0vODaIX4S6MX93rQ8wGlcOV
4Wdi7KpCTb3J72jqG3nqy87xIDniGjdqqZfvKSjTBVYSPiOTVKM7xlwx6kkgy3UtMQCLfzN7Q3RW
4sfkD0IQBqUl/Or+H+NWpIfUTn4a9rQLr9SnrXKR9hd2td7AjN5xE8dPG/Kz1DwJwMe/TwIPZYSI
qUJA7AGvtzHBt0s8d4fq3BrcX4sJEDrZrwwnVdQf2NOo8xSIdaaAkYj+/BGnH/JHGmB7ahueY+IM
WPB7kJ+lHS+kVAXWrkbJRQql2lVPPx0vQMwO3kIBrlv+AaXf9rXUs+dcB6n2+VqVB9b0UjxBGopo
devZcdDn0HsfkC6tdXu9Xys9Zfi8/ipCuubdQtpNXZYTnLiDMBnLD3prFDkxhLT0dj5aY3Gx96NN
aiFHawGnYdkWYfTOa+Tnzyk3yVPec7V0vnHIS5Pg8Zl68rTd2xbWJgr7VAKD3rhcI6s2+fRQTNf7
B7lik8mg2RaqSgGkX7t4ZeJSwC2qcCJ6Q5ff6hNryW+d80f9EtRwEUnv7V8KGgi1GTvdNrAPp/Ef
KtsQe6lI868jsZQJbg0+64Sx62P0VBOZ5fgFeyoUDr+7gJVm3hIpzCzQU6uZwA6CZcNySTHyZOxl
iRBgfqbDv2GBhuDGtHcra8J9lLbQg8++bfPLBPWrwqtTj3Cz+V1CkrL/Z3aI+z8r0TQs+wTjnXXp
h0nKfiOPsiUmTIU5ekcDyDht6/bxV2DBOBxlAbEfsPY/YcE+epRuurKbl2EnpS31WICBKgWmI4is
fe5gWQl5HxWsQQsqXuB5F6OHpKJxLtTugL6gyutNBW3iCdaXMmh/HGzmOn/k7peo74WuXNjNg81u
YsSQ2xRBMUc0Zj8Zqv6w+thQXfmjt4PSoEXiwtdMM3AbvgwRJGQuskrY8RaTMxqIQnRRy6tgwpnZ
S1//JFm2pmHiLm26fWwH2wLAwNprdJUkqk+cWchWIESvyVcH3Qsu5tdTjLJet01KkjuH2DcRRyKP
cykvinmqDw25vXDfcYHQkN6fbWWzNoKieP4nlgGQHzPn0FuaiRrF20/yLNXpMivMSmuk6l98hBPW
U7f0ISXu+79C4BMjsXW+1pVzqII2LTacbXXtkJXBcOkZtFN6Omjex2uOyuU61UjodG//hqHP+pG/
9PPq5i/zzAEsJG7406gWWrhUpaKYAHnJQCAgqlzjYOKTNJOsPWZ1r/Srf+J4NOHzJL9TqVJmD7LV
snEkRO+N5vM5BR2R/3cUdflhzGSIYXtbLezjt6tXO8zN/CL/lLtASGjwsKnT654M1pq3U/LKHJBK
IIZdVhMi3PCGnXkyBBx5oqt3/V3fP2mD8elGOQwDbde/iDtp/LDk/SNeqw5MwSKQarH4GlA5mw9h
CuqiZk76WuQ3cPHwDL9fRqRpoaIt8LUgS16J5LE6V0uu8MOPs+AGQtCC/uufFcYNJ/OKBPlfEqhp
+QwciGzzCEhHC6Tck3iSnzcSyVj6d8ikbjoe6j3vvUhH9MFd/ybolJtwTE5qAGoLROCFQiYPhmsO
dNfVkJjbaj7rXx5Dh8vTxA52gERX27qM19A9HmqUNMKWEdDeWMB7WZTHTeuufViwh8lyh0Dix+6Z
pdyEgaqveLKcsKJTopNtYTNr2QGi4hzzBekWkdrcT209NlIvIJq4If6YwaLiyssj5PKsxI0xeQVn
bSiQGyPWQkk+9qR5OXKaeBix/ysibzv1VO6ZGyoAT8GVibxrWzXaVdJO+b+04A/TOXYVbAq2KF+a
7Zl4UaPMbSMB8fIHtee7twDeGNUxrqT6dYOwfh6cDHw3bl2d64xXsfM44x3D3LOh1oVQVozxFKgA
e5bWB5cokzPRdUm4dNnarXre+HIVLZwDVS7rKErs/EviWmGY6AX3oYpYtYSpVipFeKlnV5/Tu/Lh
RygjV7WVzV7UQQHa2AkIY6uV7uz6a0TaXIvbh4A23CwrUVtD+QN/bN4EMlshfxjhg2kKBKO9M9St
6SIEddkkUjoUdUEHhl2wGlhPCVWfJXWcNdzZkZkwXpleRWNPGeR1wRDxxX8TfPkXLUv0odcUgI6l
r9Z1U4gZYWzis19HGbZgV2BtaUhhkDy5hTH1I/2d9n5N+uUTd9S1idIPZrlMBoqpNSE8/uBhRMz9
UKo/5A/ZiKjk3oenOVfp1N304+V/Yu0ipn3x5xDA0ysHnjiAoBd4CPNZxJNbwnotvSdYG6PiwAfo
qYtWCf2uFRMjYG0ABEnSN7rjJUR+oa75VotBLAXDASc3JGiqC5c4lKNrWiFgpm2M0pGgX9Y+4lNo
y8NP8oYe77HX/+YF6SSH9gWWn5OdQNPw4iyKb48w2M00rctxPC/DpgIYnuaCy+N9sb2CMPiuj/NG
h0+bBnhSGBg5VngpLpdnM2zgu5Py2Pqw6ILznNP20ZaOYhh0Z8x2TEbSBZfNX6Zx9g1PFVNDC6L2
+vxLa2kc8CpUIP6zLWFwTLnladw7HgtwVb8XyKMs2pHG9jUhszHAVdybiNbMUA88XoYFy3/S/CUa
3yjmRlOXIwNoC9URtjK3bzpC8/gWUxmhnP5MSztD3/PupnKG0YuDlV+egv97qmOKZP3HEWdkl74t
F1AOWmE+3VZ3GMomTuVsNWclLqO/4rHTRIWHe9ENSZnl9RjSB+YR5YBn4uEbQALvjIXxFLZfyY5Y
qGHW8JZFbLNkzrfYSqwh5UPR+xQmMA5wxWW8M7/Bqgylb6AftlP+4yO5o/Ah5YKNhOVj4ziMsnrn
ChKpF/+qLTaI2NA8oiqFDQgr68SCt0XHIFNs58JKtrVscasWk+tN803bTQznl1tT2xbap/GYHTa+
L74vm2xT8grK0I5xwOhshZNJvbtA2wOFj7Eox6/iZ548A20yi8c570mFuzXqXEF1VlMa2eJJTzdv
+Y85NZ1cWUm+C2mQTB1oN7iTgZQOTEbGnWYHnddvvjAaYB+MgNTrl6yXuic34nLWJPXadEw7zwzb
VI2O4SpjvS3rpckQrXnK8/qEivqfb+HsmMeAqYPCSHfzGc9pWVUFlwAPXRUF5o+ci83xKPSQ3zbQ
C9YgoQXFUHRMdduSgfTeR/JpPsxuMXvPRj9wAUFFrfl9dp8iROvG+8whsx3keGJxUefvGHKi9wxU
IqYvo/SlGUoZ3ikM0PCO8/0VDph1ezbxhEa+wmJOjuTzxIAarLLAHzIsi6VAP8C/nekylOpvkIwr
4IJVgL3upTcdgyPT5SMC9u33dCTpupAfXc1vtOrvYqX2VrVHoQz3zJ0eLzA+kUt6QBaqyKl/4PCq
Gjhq6VL9Jr8CCSgmdZnbm61/iFggyFlcJqxYorwFhSZswAdohu5i0YFP7NBhUnRqcThOSaEpiSrp
JdSfY29fhCu8WRgbpIIVYvjkuDhIxXlgYZi4bwLvopBwH++s4jMGqvyXaDztWBDxHc5uHY6Xryf9
tWeG8UwOpq23gRR3PrrCeWRg91Va8ZjU+6jua5Yzn6ULwmA72QNgcULlyXlg7VxgZhAPNtUhQgY/
n63C/ftLfogauQ936KYxZyjzs9QadqSkmOgrK00+0Mpwhfg57kqGV/pYzz5ZLUy4agkHlcbOMYvJ
yyqRHW1rLxHCUPiX93cHgmIDKgN6c2OIbuz/jirOgaWEk5T2gNOhWjsYdMa4JCgFAYuWqBh8qSaz
Ezd2/jZWJdcYFhd47pfCrAxGZAcQp6X9uTxwWxblm21dsgmLJFl9j4FJ99FLLO4ry0z05NW1hxFp
Q9lvJcyMLYqi+AgJ8WQDmIb1ztNpQB+HO3q1RocBYRcOy3v+Xmg9qWRtWzbFL++rshrZBlYabHHL
pXFppLj78V8pCV0/Mms1Qff3VnvFoxCxOJyYMGRobVJzG/32VBPE7CxQ77Q19lA5nIDzkV16gGTD
7OgXFQ6EEUDaIucO3JIwads0djlX1vO89qWXCiuO7Twu+nNzZs35etY8zC5kOzlLi6EwFpXBbTVQ
urPDnlwg7pzYTcWCxBZaT7EOFBBkl0G6bppMVOtPApH8GmN0ZXf/WIEURSwyRpbfPvhhSFyrGJzz
5g+RB+PoE2ScRZ5BmLMY3I9O27CHEyYu6MXcGj2MX6WJuam6n+91lZaPIl2OesHp3RJIdat0Oit0
UCa5tp8HEuB6KxlHUNH6DN0rAEgQqwAKeiZwKf9sdXrpJ91ZwMnS4UDH5BON2kDx01oZdDs8CkMT
elBTwp1FCLMZZ63OzoFGkgzmrl2XdapIBiPyEICYsIAXeQMykIlt7jcJoK1hbNhzJBprXoAqOHmY
w5ez+p5gglTjcWZEfvfYYmqcOobhMXShm4oOH24GAeERGltAhMNISlGUXdpQ9hg8LIJJTXxQ+wLu
9O6gim5/ZDx30cgptneOMJjSABVJGlc6PioBtNhzq5e+l8+xXl+UlKmNCwbimgRLCSHk53oeIxXC
Ej3KMKJgSPRIEAwn638TOLrIb+8W0W3CbdmxhhM0pe3M7bBf/Dtmy8iU1sRFMeySDQ+1Uc87+qBu
8uDVlFUzmzBsBjdC9UlO/5ZeJJc4Y56DKDt72knQyQijm4QrWy3g6ay2ph+ztImzAmqumiW424wP
9sXH1/Pg9MySZMoBZHJuna1c8UeEA1Ehzrv+WazVR/jrsXPYG9Op4rfzP6pRsabLEUlzdRvpKthe
chp+nqq2ntuLeKLj0I3VrwIH5LZ15T1KQFAlTFPYtf9j47XO5sUAAG+OKE9ZwyoMCPajikKhO4qJ
XsIvOFJKx3VggWfF2alW7KWMMMhSYOPICSh5W2j3aB8po9QET9vfr1bhmO0oEMU8Tn9yPqdUxBxH
iKxb92H+kFAuoOonL0F4Jx9XOI0vGHKW+7XEMHzctSm+fHi7dDiCrSaVSS7KDhqLDmrUz8PoMc8F
n3ktQ76gxu7BzNyUwny4WK0rnWTJVd5ZlJNIAvH3JvSOmZC6f/GnT5KbjMlppGpeCzyiSsDix6Cx
y5AuzHNdU2g3EVZHNpGgeGIQoPAt2MntZcjwqwHiHdkCImqRwOr22De/iQ9v/aQC1hPd8+pBqenB
zJueKTAjOVwZMWQcsqRClzVUWE1KKY+ZPhAVP3gVZq21xqW2tjvAqCt8RRMzSDlLZyFKTSuoNt/E
0QTE2A7G+jStfNiLZGfTRIMd4u526tN8fu7UVB+PnlEtjC/x3ZuAPmv8YLJ5CEgA5Ok4MKNH5d9M
6+bX7sYQ+npSTn0vwDAiKA949NS7GJH91u01fQ9zXjqCgJcLLgyoI/M5IaGZIBtbIk3hzzJFKt7h
/P7opFdaucFabAhTnfO3xGVzDNVrNG8SKcdMo+nldlnFJ1fjY78lXt85R2afURYdX5kkCP8dDppZ
0lDH2kMt9PfsU1FyqsP/2up1++eXqsymVSnNITR66ylwe0ztGIDmGJZ3m3NQpZt1QQ5kojz5a771
WWUipXWeUAuHkcMMTyiIK66s03kh8CanxyS8g/yd/fGkTZIfDrWxlHpeX4ZqLr7AZlGBY12vZtIu
BOybHDDWhoSQ0L8gzpEG8ToiHWpTr2Xcsll4jRzAqQD72mYd29nfjSYXqbJZZn2nwPQIFNZia065
gRqUYLoL1HXay0ED1xs10PrQBKaOrocH1y2/HLVLDEmXfY8FUAGUaBsTW1EyvjH7gVhHZJpq3gBN
TaANd8yrGnlvfQc45dh7s7R0fYp2kb1n1fRgzyWLjCZnIQekTanQ/mBnMs3SYfqD/Ts98H/iJeyp
5GjVEX05AaQmmxiVtqPvM3RIXxGTTc3P9v8ugr0B/ZqErI3EqkJO2Qolv1qc0BVX9KLy8GaXCkR3
AfW89z/gJvkeg1JuAn8JPOuaY6Ss+kx6yuK5U/x17sjbXS7/9HS3MYFuznDkhRHnaCaja0qPf255
yu5uNkIRpZHrQYB7+keRR/yIxafSkoNI+cx6ftr66KZiLYGZS7dgFMXagjJr+cwkHwuZ7zXLKR7T
Jnrvq+gU+dGxcSvC+M4/K2N/AAcHRZYSYV1ORWjfB9evQ4Z3CHNiDPPvwjWjDCZgTfDEIz73diS+
HPc7CdrgqHcGPFraOeIs2ePmIgjcgJCExZ7t02yKQ8iwBIkTNy89yVrXgHNwt93sm2u/v55u1Krv
KVFgUHPiYWM73x665tpdIClk2dZXpkESM19wSztfubYvYicy2EhrSIzkM9biTvIFQn1rbkuN9xM8
sJU3gZpV0QHqXTMKcx9PwWoPIQAHd10f9n5JlcrwwzA6wZm3fQ4WwGqxxJaWMwZ+ZStY4vrmMUiL
wdbrM0sU4UMNWh7i5XHwlrrfrMK5G/jBN0+ZHXTadwmiwo79SeNbf5+GuWsWcWJv6vtZRl4QrwYn
RUwp5pDrQ+Hky+FOX8kcqgnS7Eh8AI5GTVQ2K/QYE9o82TsBZpMPvOhS4aoflLswetDLkYUnRXVl
Y+bB86bR++/k/CfVDBnnzheO6N5ShURWgJWxFAbpH9rXQYDR7m7Bndgcu8gwvynPF+aQIZ3A0ix3
nkUox5C80hosfMMQq+Mj4IkQMbY0u7P2HUEsztEc19gACu9qzDLlElpGEUA2yUTJpmQHYdS/HTZL
w1sSCHkxbu/Tagav4QLN0T4rXxW6gW1l4V840uarMnNQaJ4MFWvfLg0HC3BkSbySPv8dGJd4AHpM
m4sL7wlwDv+dR9L+NSN3FBqIK7dr7Hqza5CPmjcZTZFsHlbbcKiwbRSeFw92Esgz+BvUniQoxLlW
2c67qoDQ8yMBRsTiGhA2cvz/XGWtqKFwxa5yw5aviKpyxZ8SsBkI2ae6tbIfG6FbRTrx1YoI6N6K
F0oXM5o8/bYfHe8Y6OnJbSh2LwOHKxwfF/KlaIGI4e8d0MGn55faQJX0tgqFayzgS7EJiTTr34G4
tQx7iX/X6i0cgzA2Has0lbCwmFr0tdMVm14TPVbdmUoZTbVGa7Idqhw9WDS1Zpjirdu2J93jkI7t
kIyw3UG5RoPglwMonOox/cyzpqj7bH85A2Lf+VtrzEGuPWBHPI+JdrYmgl6pnJFVUC7WZzdqD+/A
yjh5YWakHSmHenediyVO3MFu7A+wUuSwZWkcJM8TS/0qOJ9HUUAy2D6PhWu2HEKzHiq5uaTsBBxz
cU6M6EcMQiCpWB/ckK5MF2BroLx2nxajt0woBgLJ4YCc1I1YFlMZU5pQDiNJOQwjEap7Ny+6Q6ur
G7iJYvW0BLP3v4znoUGSW1C5dq4MdSHwANfc9QRMZ+q+IT9iD8kZJ4roYMtCm8Dk/gXkL6dXBJVN
Z1JgrpKGmUYmQUU9uGIYteP9UdknCXE/FaLNQW2h3X3wf9z4xAsj4JIOmY5csMR6R4x2elu1ecG4
aCbjR9QT62XVxIpvSJos4pBLijot+QyA+jsdzQBNJ54xS7PRVYQdWm6q87HWSx8O8EBs+9PZgcN4
Q6CEH4ZBXYw2DrGvw2igFO4hVFH1TVGn207OqsnFtBzhGRaQ1LB6DAYQqFLAnYZIFu0aKmRau+7Q
A1JxNPMmQqCZoM1DdDivNrpMPTjOeQ9ZeTQSQkAQnzMPmOWr93JluKO6vsI3d0zF3aOFkFSAHE5A
GjtnlCt4Xubc8nHdMFdqp3zkfh8e24RMKODBX6I18Jp+cGlIYR/D2l5d9GWL58aYOb7opRmrRsPs
uBKNEiwXjEeDq32Kt91f1SwzlQQKLgCeaXM4FE5AZEHOhgrQXR0UF9IeC2EIdt2RbgcHEY8NGa+Q
jqZ0sNHZ7Q1dS8MOwEa7ddF512n5OCcUAXHPes5zozJ8bsVASiInZE7vE3JHyKwhs+KudpAN2JQv
DcMzvrylwAcRwv7SehLflde7n0rCdAv209ssGAxWvfktIf61XoOGqbJwguxwSc0kT4i21YAuFmkc
bHZoYwIsW05vyBGFQ5vM/Dt9/qRloH5t5Z5gKlObU/0A/1gK7eJHhb/BHM/tN/jJxXhIFYeRYzzz
37Eg1NVu97GcfFb5rWPErlNJjQ0nZjMFcXkiwwGqeakHugh3gD1tjRr2sM3IRxgY6cIY2R0V/NlG
6VwQ2JJL6ffiQ+0YzPv8ofGsTk2aeio1zaliwL4KGZjLZxm2KImNQefpnbzDcvr/wZ7synarR6nu
yEpNNbgnIkyXzsJHzQFh6YBSyjjoaHtcyEETWCukONqa+Fsb1nA6PQ1uTJ0zm5Vv8EVQMFFfVl2T
hQeOvZpeNn7CZ1e4/ryzIP0MLydvYBtow3VLtTtPBwp4Ji6CXno554xZTnb5di2ubDd+OidYA9GV
V77mz8E7AdS40CudBgCjo0vHbAk2nxOvF/DN/2RmSDO6GhgR1y/tXZKECf66Xa8aMDkyADMsE5RV
9lSfpMGCXlozhxX7IAsoVFV6vkJgk8AMbbBC+bb+0SWle4KmaVuk2ZyLIJytIKZDrpABzqX0Fk+d
IIr2PGhvtEGwwPjqh40DHODkF8UeK0qB8Wkij5OjJnDomrbefaOLxAeqrI40u1GpAfDJ3Pp4rjFN
hfwo63r6lrGBZgrF8aFQx55Y8XpzOyScgcgwKOfMAhiecbeduE8KOgLTO8TRTarpRudeYsfZvv6l
9qQpMq47prEoGGvOcsMhiLsmgOmXVscwyXR06rSf7K08rzOrfGT+8SQY2MTeyL90l4YqsDfW6bFj
NCZWXKRDIV3/dekDtcBrM6rjR1Xg5LhOpkuxmZX2V0eEWYnghKo2vDIbY9y819LS+w3GgVvYrQZd
7yygtk3C+hycSHPjrCcaWM2cPXIFPr5uXAKZiPvf4v5IKWY+4XJ7bXw+o5FPP9Px6AUsAyu4F0lA
8Hx7r81PSoRqrXKd46tSlWrP4Q0Wl+q7woVIWIkiuITFODZ7NWa+s2E4H/9s9ik2aEXk4FdnDrvK
vSMgZVLAz92rKG/06VB3CI8dMGnuqtsdu2uVsBTCqCTNfr5AVleoTXu7q9e9QwGQcoJyyBSqdpd2
wj9umdnVlhu9D5MC+0Q1Q/BLOLlJEUHoqQ3bUtWcjSogQRSZFbfopuANoZLQ8DqojuBbeeX0TLQn
kIn3JoxqQZDKuoGsCv8/Ewc5fIuOudCyK8novcPoMa9sGBzgj7gG6SMpgi2fTm1sh3Qx/On8WuXR
Nu55W7iVh5Hqwbr592STX8XlsV71Uz2k9Kp3n9SAGTcdAI/sgKni4/980heL/QPW9SXjw19CeNSE
x41E+vC2gXs5jb5/kdAL9QV6dE0FfqMJwt6d9SYwY6PKAlFBDft7X8lEvaCCL9u0S2TuAmbtIxAv
XDodAlBG1qN4Plm7VBtujc6LzDRCV+deahKYQGYWDzN6JNEz6Qtl0oKsIdSgE572HI4qUuLmdzH8
v3zlJVZbjuqpO++f5fwRLphE56impz+mTaSGBoc8lUJIPULvtJRXJ0+cKNwS4VlGJz4WFSUpbqwp
Wkxl5iJBwrWT8GDIB8Ff+b4IUfQJtpR1aYuwVRxtEHJ6SiZjY13WBu6+ma3O4CdDg6d0mEzvgzyL
7x/KrriV43MjKEP8i+qYUlczKSRmgoBn0Sm8wcE4n1nvwI/DXiH54N0nycTQrBuUgVzmdbFJymWY
XAwgzidKEmPruFuzIFhLDh0p+XARA47ZLYZkdyflNtQtjbyUdsxOOq2v7rpjD1eLonCTI3tdxdYJ
5UFb2NVZsqiLaZfilh1Uz3Ej6/DYdXatsvRNR0Ur1xwv/R4vF8Rh7QmFQFgTDnfi8bX27fJJF6bi
4pvfpvwZT0wfcgqiA4fd015+J5FT6U3Z2ael765IJMOJgYiU/JC1IeIdyYBezS0Rk0E9jeNIYYGL
9DBAad/OzndSkH67sOu0ljBSWcgI5vSkDaMo1dQebae/vKE8a7p4b7WfNyNbQYN/oXQr2uYL0LnJ
+tmDUlBrbdIbjOjhYVq7bwF+k3tCY7rcLXF2O82sGb2MaaiQlOM2YDrYMLzfunpIQwg4R+0mcT+x
cuCWKQh28MMonH18vNQdwq1Y0R/oo6gewLHOGFfR3swowxoBjzotiiM4LOEyHEBq1y1w6x3P7ezN
/2QU61IsUQQOnAXA9Rr3gP5n9/HKzVYz2pIMs8MRFW2TfqKsV8TH8wSGIF66hYW4TfOM3nU8MwfZ
n6YCHUmyUPJ0oHZ3n+uDxNovsRrxE1adDM1rl46XdNhyP8RLejxlAwplhTrCqR6UW7r/k4BXubfq
4GE4mQtLEqe+nWLhzG9U6LW6mMFT/bJZLKmhEh6WX+iSLurgIL4s9HFd4SbQL2MIMHxEUs5LDJue
eKAvcSp/9+Hg+kEPnAOlQtYMrG+fmdZ1xsP5j3nQn1vWRKy32MNH2d+m53rPGAqNKrTJw6oEQgfX
6Jp0ntK2D3Ax+ENevfXMX/sUkHC0jFS6s16oii/7dSTrULmygO0Inay06tDyzAKXADxeWSO7n8FU
wk3Mb9HAwUddWAT5m8q77coaxWaeeAxEb9DBLJBw02YCV6wwhuc04xqRKW+9bSuMu1ehCa9UJaSw
jnxBFQN9v0yrXyrQzbf6qi42wbf5/GKWV9i5Y81dfKVGG9+D597qi4eite+vEI2PWUBJIntaxtA3
fs0wiH1ldjg/e3ozPHUQsecHvG6zOdIELRjY295QdvhaYcNoZCbbwvUCIpJdar6+co2iu3HoAuWx
rzpyUW90YDJ+X4BF4/sdIJ1aInV/F1nWZCSj4TeJlESZuTVE80rI2zZur1l8bTUuU7wNdogdslk+
uqnlncy742IK6iBX2Gp7ZmB0/KZIuWBRcatgbBU6tL0wyb6xjhOXMHAyizMQgImLi389pEbyrnrw
DMV5Gi6WYBkWWTf3D5WZvW9P8dXZ1lmW/tFQ1OQYDXxgtWYNtNNeuNgkH6BgAevtxnND8toTVaRB
NlpL024l3OuGl9eNTgO1m4W7hfkFhzhZpVWMbw7JxPxdvL9A6belzvSQ0S1ONbXZx9hv4bTA8rpR
V0p+y3MzjcLw8ESyYYwa5xqRoqD0KYOpF/5C/lewtoYy/CWNGUwvAmTdFq1GZedlCDTeZ8fzPJUL
rs3zWh1cqvCa9fB+hF6UVuG06lmOOwFp7yGDLc2/pbZNGJtjk0y66n9gPgUMlLrEoP3IGgUByMCz
+LesQUa1gUW3tJ446ZraGooCHqSIgBQgLznHEnDG9JKLF6EGnT+pML70s2iP808vUbIuqIQM10bl
E5VYSudtGYK/AKbma/qyMjSfzHI+aej7LHK3PV7BMLcWUycNmLdTe5XB0gPzUswEcbZIfSw6UX6Z
Sbhu8qN1jWabMv0WLCkKR69i7ymWA5vr2OlCTF7H8JvcUxHRd04DGf1bh/0pDw6lMj6ZM2haEKfO
1/FknPkc80QUnyRZpdeqK3rgvzvaPCLcnUzVlEmVLueZmeFDz0C9RziN8gfSondCWMrWK5UFiBps
N4Pp5gjaHyjTSvw495QBEt6ixQNet4ICZEJ9wA0iRd5iyb2OGJwu9tf+t5GFaSKr/eGsheO/dMtZ
jzr93NfPiUO/UbmGsxlaZ/TUG9Z5Lw2FKkSFVIN215eOOp+usVHAQJhgCorXQk8Z+EG/c3Nnhr+R
ogFaOHc6j4TtpwR9NdBHFZn1Yqac8rkczPEjn4yuuJ/0lZXejeFpGlECWJ42BSXTj2SwR1ZEtvLs
ysyQWXVamLG+UbX9et4N1mCNNFJgoGs/b94xJpDhom+rxrQ6ScZw2xgxygNWfc2Ts7td1nlxZrSL
iNSRRpAnyGmKTuT8HxngOlRfh4iV1fRt0C+J2LNDsNRqyW2RsOLp8cmyCwOTdArQyvYWJZPJ22sg
YGsFd1ZEiumhxWsEAd4+cVAFbFTk3xnO7+98cbWHvtbGFWQZlLPqcIPlZV4CibIRBghNDIFUmcdD
sbHO2kDbawCqlZCf6gnrEcOwH9X+gWlLXHagFTFXrBOIwfvxSDaa20qYD4p6EkmfLDQ8QVUgoyuR
wDQvVF2Pm2GKpkZy4qWKEsOVe551+KfGjTP35RGPiSPc8hkaw5pYMr+sCQX8FpuCkZsc7aBYnCDi
Vv0ApDVrYer+/orVseoVsMh4X+R9QVikWZIIZW5Gs8TSwB2/kjHM7mhKaRBvmmBkc99QWF2kygJ0
+FLXJHCOBCEFijUlLoYmxEzkqHDEmJXEvbi395PRGyfSMGeqsnYp3ag2PHWPyQ7gHUm3wTdHkACa
nSRrzEjQZUFu4C9SVk6sY3oYGn2++xQaSbiMaSKuJFAoku+kl//yA2YFxbYyCYSGKglAUa0AYFT7
nBushCTyIX8D+2dsZQodpPuzE4LODU2+MuiqvBLkLlHKfImdqNRV/aNlMpqvfU1ZZaz/kThCsYrQ
SFofqzzTCYJfAupaDOXlBvQqMB77sRnF3U8RiFHN8OjioYK4lrstmLdXzaN3t48Ucxc5fW9fMA0y
11GCtq1GdWrJBhDIAmcyzs65d9b2ZfGfpvpLEtGJtLvvk2up0nNPa8xYy1MVyjOA41cXoKzDmojk
DXVWyyEt4jIWjYSNQ2KPo0x2COVUqmvMpGlW7aRYCCTD9R/nQ0riyeHNX7G0asqh04CVUJm76swi
r6FMWeRFo5St9mLv/3C3vq+SLa2vppTwxz9oitrhu619Q9SQRUP/12tzSs3EyuIKYgcklMOtK0mS
1QhjcPNmN7tRVg0KP/vS2QLXAqrNFDcTTu2UwbAdaEddNvZjcz9YgblyFB1aKLJb2YZEhKPBNB79
vgP8Y8QnxRsmAfbjBvVRzvHe01yjGt/BBSRacH67goe159jUMa0ss093HyLBR03HmAOQImXPpW++
FNVfid5NGU77Hjlxmfp4WmQ1wW7wPjbjLevSWephKqnTsKs2unG9hx1M3k6PhdcGDM7I2qD4B/Dg
NocNN6Ga0G+QxAFfehrg68UCHNeRXNslDItoJ1scXMjJhAxK9NBYCKwp+IWqc+6ut2PoId7zL0dM
lcrkgGipu4IMuoKHiwrxKxcCmCC5T9Ue9ZjCZx51nS3/pzHt4szf1uj1Y7bcvzCMLhDbvSJiWu9N
vNsnBgvN0L2N/1SaTy97o3GHiizF1ti+b9bgurMVcIC5Nvtf1ug1RFkb1p4Xmxs9imlHHgPhtih2
8fWcdhnSkyfO9Yy3H+3+QaHv+5QDSxk0DmXMXudKLlxcpKM7pLy6KPQvLqrLfofa7buTAvvwdYJ3
k/s9qahY1TKcCN2qGupNRMysoPqsvWKv+VD30iT36y+rq/t4QPq26yObtJ4JGRQQk7bVSfGcUMpN
d4oxpSYNRQec5WwqDnb/168NpAqEYa/t4AL7eOKSiZkPo9yNWTm9UWnnz/VKkhrZxmsX8yJjG4gK
W7sKVt3/CsOmOE1+/C96Q+NsMT/yXL8BDH0Q2Ajnn8HEji8JReWZS0b7KC1a+pC+StNU9Y2qCf3F
Z9YoliIW4RykScsjjcGWKer60fh18gNheMBuLgS0WuSIAYc7EGRcq/5XiyGywMWNDty5Z7ZBzl2h
voB4433c4IaxlfyqpFOmx1bsOdJEp6uIhFfnGbNNRTgygIPpRuEfMARn5YyF18x5qtVUNniNYCjm
J1bgoawn5uWXWWIRKkXjDC4+ZHa/HQFcjr4tVATXjur5GR+kskDYR23aUnaaSI5SB3I3E7BF+FM+
pfYlr+EswaiAb8qP2QMC9GcBNKduRq4ZybhtEmnwaIc5ZbgEeeQmWwKStMLus+GEWOnscRgY/O3P
F+vtFlOjLsut+9FMcsUsXW8ExS0mrwVhznfy5iF6x4cVOE/vQodH+pvjVESp5R5CHBUfaj7ZgMcQ
4zpSRtGaYCMUa+f39EgiTOJJiGq0HNPUVgt1Y9h2xuh4rWSlGLwFrfOqWPM6b+N1tSaenXj/+tIg
BK0ckABk4UzP35bi2HARvDnHoqqFsCnuWR61k8dhGiC60l3b34MeCWB0iFleRG1qHYcL1fdXKVih
KJEdMkixcjEhuiXamOHR+CA9WOGIixSl87H2DI3J0sGUNe6AveiVeoaf+qr9boXsTCDrLLn6NNWH
UUDa+BkCJiVLiFSG2WBvUYvWna7gCjYbwAEWxIQjgd19DL9ESDdLBSTkclyaRqKId0qp5vkWD+ed
qp/OWA1xKN4AB2kk5D2kpLWqobA6fF5/Hj14ZsdV73eCPx2zQD8QwgcqE17Nz9lhiKQ21QGl75tc
/hO5FF/jzrLOvcOIiLeUTE8iKY3qWdbItTL3SYwR/7Fy/HBeuaOtGocT2DjKxvbvLP3r8yX6mgTr
CLAh3qTCoSYtiTo/szSxouLPk4Ggiz0WkP88cywVjdUVex9fSWxpogMULIUTZDmdYoQrwAS1BeiT
qhQJBlXQauiDQupVfGNZLpLHmRrE21aGFI/xJPZY8CykOr9wJ4HTYCdaDg/nNwixrF+sbAEjm4qH
n5AdKSsewOtPF88esleFI7XgUJzafsuEJ/oK3elAoqAcjJooINYQIRqYP+q5WOeUb+bl4bJ3S6OO
TPUixaFU/3AlRXg5eyYTHtasWIxZ4hPt3j6ffLod+JYNMn4unXFoMK3X+rZdNV3DiGRz2ApyYcj6
ECcvvEcycvGa8mf1MitRsc2gHlsUgBizBRGoyxgaU3h7IofNNr3axvI1JNiONW6awlP1ybt17kby
L7eCtoMF7v5EGR+c9cb+Br3aJ4xyvp3GhhmC0CeVq929fUfeyYZoEqBqHSLup3Fhurymq5qp53ms
YoBF5s0MDGOnKndSHp+G3BY7jYKQyBDSP1FPZOsXPoKyAdrL44L/SP3ULYxVeViTQUKfDJfemiqY
UX0Bkdt62GSn6q2WZibhv5bqj+VKRBgKuZzuAe3xmoTu42Uo8aGilXpOKQCNvto8V9QyikZd8eqF
bgJDMwCa+fgMuHhQy8jnAnpyMpodb73JS3CdxSGmXAi4M5/k7rPPqcZyt/x62YXPcQv4hWVnGHbY
Lgz/KNp4JDni66Wewu8Yy6q32ouTcAUwcFmfNcexkYCqm5zFMwqNr8RBx5YJbl8oxX/MVlBtlix6
cxhlb9pIuO1tPWgPlD5c4uxw6hGc3AVXlnuBcfrQe4ZIeW1nyEc4KJcWCnr/m9+VQxzmSoJa48nO
P8qQssUZihz0l7wFFWmnzlX+3Vnd+NAn4yku4TB1IH4UunbGjwcWzvg3Z2CnDMdAeXZZ8wgQ4V4Y
TfB1A6Mb48EdsRYF/KDu+MVt8mcj1dxenFTkOHNfTUlMqoc+qQGc4gdsDETvmeXM/cwMuWn7g4if
FrJMDjFmztTujcDLee2/bnDrGCY4JT9G9Kv36YsKUvJ6TE/etIQxLxIIiWEBs/spOZa/LPY9xFIz
ClFNzMQ8VOh2hP2wbTOHesryTWHuN1/76O85d6ulBaHbDkNzXEhc/fNHovS+mQUqViVqUA0Z6b18
RislZlwjjWN9Cpfy5Rty0yTqLXMMjco0ooZWMkxPoQ++ZkcwL12+fLNTNphTdyZS3xZot/ZxoJ2r
nnjftB2/7TErbaDyvWrNh9WePNxvHIu00ob/87fpgIIFwwcZCLSLm7rFQYoXzDXhdF93rAddQrvA
v+0d1Oj4KZtUK3OpGKxsWCha/Y6zg7g48wB2JVsFQGA7/JHMsc0k4VeHmaajDSKCzmyvSJYy1Nn6
pxgqpnMXPLL1nIHo5keLinZ/eArA6WK30KOYwFCx2VxfMvWl1smhBrSJAahpPbbpSyEe9pFIogjS
ii8GaSCnZ9OwQ4RDOVWVEDXPLq7ji/3i0JG/GhU3Jzn6mMRolJ0VA9I+vLjXrT+vZhYl0smnTTD+
+Tgi2Ah7gOiPR1ZDL8OJXqjPMa36k8rzJnkqtG07bM/mKR/AE2HYcd+z4enyHphR8EzdLBQDPsuK
9U0+TqD6yBjnmurqiCn0rtpvnrwTReHITmXhnqQr3Ooayu1zXtxTJ2lSN/K2byU6HEL+kbK7G7e2
i+3FY25KCSaUXtVEg4YVEqgauSAX8NxlPHZ1CAY5ElQvtWVmL4vWjZ1ln9xJO9ctgXAi8/iyL4KB
fk0d6hxUbJ3G8Rkt6drjCmF6SffZ+IIZMFTbA3hPZQj9FrIe3vY4SJdoGLWcPRKweqvSuJEss6Ad
s/8+SiQpXAO2cmmaYSN83xnjwVxvVxxgmIAiJOern2VzExmYWZziRTaYZNdcCFF4R6G2c5oqI153
iTtIHMG+pHovRDCL60dc3O2aIYH6YUkg0dufO2swPF1OTqBUiYV5mqvajmd5UdTspjOzIlSpljhm
HSJM0/bEmHQ6P/0bc3PfYxc9kEL1R9Qi1RHXlewKn6+r5FodSho3rTltzzqGHXpHLwq6B9JvS3cV
Jr1QGUkh58VZLvomYAnU7FYc5RH2uA7AhPzFUWDr2lnuN7kvasKWHfW843txiBPYl8IEHIN3B7Lr
srI8hCvTj/1ys/d8OUgcG5iUMcQ9rz/XSzECBgbLfC4Fp4b9KK2vIsfwpgkCE0hl5ujHPaMrgAz0
kfQnn+jeaey4T+jkdi3gH/5PlTKBrbDQFhisYTuBZyVaEQljoCwPxBVvPnByQqmfZ5iPjmJEuCMQ
oQd5eFmpwQWCkLe9pKfEIcfaoHxfqXqsSGjTsGuMLtUsQJp7fS/JhAM2xJwz4iDiuv+4l2/L8Z4l
6vfVHnO0Ujw6cjUosS8fAydGSvJlnlZPqzRhPsC/Iu/EhiNpo+tn+0vT9vGXjhkXZ2SXHM4NdKt7
CZxdrfayfUOiJADTiDbI/BbJR00btUNXqQdRau7sISX9Ynt5yolCtGmk6bMEQsZUUAq6ym3kMJKF
5HyrPn+vW/AmuM9bKzW+PF4jFA67rEQWxqrL4WUCs5d1+7KqMn1DhvVSw2nidp1L+XESjyLSVCdu
NfA3czkitQJQdC3SaXjds+HNqHYS0wLrmk85RnC297ROy8sF59k/AaV45M6cg/7gAI2OegUqKWxr
/d+93o+Cv8ix8wWpzPCv/lV6pAKrLt0fYf8sWWjHqixK/DtBNcogabE9CJvULlpfjD2Ha+kRJ5kQ
N6DYM7OprycVSyaIBI2RBzw+wD0lWNaOmYpog/Se7FpNyJZ1hWfP/HtUafdxolQAN2J+YmOajhZ/
JX5EcEw1rmaOjalGNp9FU9zVOrwh59Cgvsm+/FUVP5Qbtp5wVckJMgj8C2dpTDM8T65GYAzno34n
cH0YN/VXpTLCEekJCqzTyHctWndQdjVdPu43gdV+F65w08Ugpsz7AhPY2a512x9aLj/jSf5gv3BB
WSgHWyp4wDuz91Fxw2Q1yNkkCROre+aXukIHHmcCLbLNub7TAB/jexIju3Qro6HoMESZcNjN9Kyu
tBrYyAx5owVQWQFiqeG6DJSNpdetJR/wr99DICaWOHl+cYbp8Tjtu0B980Vxio2gq+etd4CFUC6L
rNwWpUlM4M6qc1OImRruyP7DN6lpzHXhZQCzlSn+dK5s7e2khORnEzywXjq2PZnom9MMdso1HmqD
hGxDqvdEYX0eKf9jJgkkecVQgDK0WT+ED2CwR7BtPiZTbaAoah5Q1dNq+rD3Wk/VseDp31dFvg20
frz9yLVxnjHHUj8lw1501/DB67lgrngGO5sBkFr6CrWkHnTrzz8B3wyHFjzIDkeyFtyFqBaHyN84
Gv/Uc3jTXQNWhu6SULZj3HSQrrfsEJ0BBupgaqAhOCHLvUjZYGIH1NulbbePozC1116sTGrtANAr
gYROxMh09z4dQIoRkJIXdXEA9qzMNuuXO6fXujFuy7pR8o9G6i0xSmaQ1zZ6cuGc2fHcJzciinRU
Di42++QO68Q6+LVUMoOsOa0QqC04CXuB0Z6MQDK0fCrWd35GCBSvyRC5HssoFY2F5O64MeQJCPoJ
S7atLtK2rRFyyyfexkv6DmigTS3U8vyEDx/NVbzoaBaCinMS7nfvSofD+yzSCqXkoHQiGWoKTzzV
xTriU/+ravf+NR4aljs5TgO6hdoONsf0ei/xwJeeFYGT9o5snxR/fmFch0VW6MR8u8a2z/Vqxahp
DAnKAxeeM/JdddSHymR3fHbu21u8kPUodbU9JwRVHKg5NXbj+eIysRtHku30CVouZNeOBb2p1NxL
GRrb+XZTCRXoR0F5lbrQpIa6TvYVkA1NolOaCZUEkF5Ldz8xk+X14U63+vDjS+GT8Hmm+BZp/42l
83Eyxu8gHrh21XQEdLB1sbvEGxe9by0GEathKPFT9IpSooDAvYmpFeNClcCjLVyKrG5mdOrREO9q
tLcpp5lfNSOiKEijJzBCV6oFhjqLYbYdIcI1lqZ1oEABZlVr9ymmMRUpzzbgydQmuPZTpkYUrMyc
PFSN6V/HnBDXyWtGafRXrwyQzbvfECKi+FZef8s21IXg0ubXKGsIDDKV7+HAE+Z4ZhyB+XTsG8m8
3Z4BS1L55wmQHXbeMHbTNFmj+aMyZhK2f9y8WzEJA2K5N0Zran9+z3jJpRU45Azvlmm/qJPQCwi/
47FBJGD8/fJeJHFyLlVOa2fza/QCACeWAyovlhuTMbYhcOAMl5zRqPbj2zcO7lVb86NfjUvd3a5R
x41k3ONv+XzGCQiESSdax/K/U5F7t6vTm9rnVKCkSci7YmUirEGIK2bfbC4C+y+Kk7p4uKrO5MzE
x5elK7Obn+ubdfoEioMRUG3OQCn4scQoExBG6KqOVmS4jRn8nxd1QdAuZFbdYOBDsH1PwnuknDjc
Atj0GENTGhQZEsWuATh5czwCE3VLvHs837ucTcu+yDW825l8F3KiOx9pGFqMXYnDwMRwzsuqzGNF
tvy3qGRkz4s3sHkjYnxPVNlAtQOolry0ajBJbi2So/73iGoyOPcjib8EgSZPrg4tqj0SYLinlOze
gdcw9pijJZQkCDxh99dF3C6jFkhqX9tccAHKXqigB/uPntJn57YYcYQbg+PIs5GTTROCXQbtDYRZ
1MVv63LXS5wNSIRbGUFNoexmWTJXGggyjQTIdqEQUw6y76cJOLxZ2Vix5azAGnkr+R8Oo+ZeqgGe
Q5PXmsor7uVnViperDHHnvQpjvQ6OixizaGFG3Ed2s6JRqZ+7HOVN7K6AvHZ5m9FwEfccIo4UJv6
vY+W7txx7ZFqU6c7KUj6sDBj9mmt4qIHDUzxretYPBvovU4T5UinuEAL5bPR4r9y7D9Dq7V7gTgW
W+Hg5MtUnjLhQ2XB+tdwecy1c4Hi4NB/gXOpfRVrljP/inviV3j4Q6UTzB1XlVyAxhMXEjHK2Gmu
xRQ8cSy3iS7ocmKcAF3gQ7u8tK/IRy1ejhWhxkvsYS3iNseT5nGYZQtnWeVTjQQ+m58SLMCnsYfP
8DrU4OeWXcYC+6G7MFvNqwoy647syY7g/OXs0Xd3DakrYl4CKmzJKehlk2j31XirUUGBp1BzqaWc
5ON6bvpO04uFehw2x07MgD9ZxKbB5IfUMl6qbMAKeok4yN4tc+VjVDjIfjTuo+k9iyKswBov/gpg
tke2Aaj24msgApCQHqD4h/oDOSsQLzW3EP+B5Tri/Wc77IlD+w9/puefGNn3VHci1t0dKP7WUFq9
dqWRVuCzZQ/IqhJxfxlBigfZfFOflw1zz2m2smn5e4dmw2DIHGUhpIPCEI4Aw9jThSfniBPaFVr4
i1Gjbdvw9JmuAIc9FroM1dAIdo/bNqg6OQEddI6zvEz3GulvPgYw5MWUxqloAIR83nI+VcKuxKeb
w7DAODRBCEvWqRD/DfvH4mD2Smp3/TdMvH0Qk7NoKDoX6Sbvy522Yq7gHI3aGNFLMd7Rowr0lJLA
EDs6g2n8F1yWwR4m2HP2Sug3yoNsuZ1ASNuqisKJjf1izNz6Dd3nBRiV1lh/cqJBHqx15BJwDqwX
od6Xkuzv9LbfpuZI/CJnxcUYJ2oeeQM7ADJBQZIlDgFRI+E6iffmbIjSlN7Z9YaAwOmjKypC0Vre
OhDg/nrRjfJ0TDjvSbjvbFfIl+jecU0ruofsKs3ULE6JP7TybT0opTOv99bOr/5t0tPb6DG4qsqQ
tXcF/8KtY0/GlXdfD80Ucao/Yp5CHojzbeT2RMQZ62MMksits/lNtAyoV4yRHEP4DqhmPnbqetTB
wyRYY5nl0Tk2G4UybYvgxZ4CJnIgVukp0hp51x4g0jZk4W6yYdf6xaCJksbLcGgapZVMNucwYvhp
zCsVXACUe2CoS8sV4gcrb8LPQ7Ch5ioTq+HysDVRXAYD/eklNteXUpeEVy23rsF3VnQag4RiUUy7
O4kiMekokwuqdVtDnChV+EFISVIFHSLoosat+nt5a4eyXNYml4NRxtcCV73buCeD1o/cuc32Dvnv
GPktEo109sPXe8CGu1aSZc/RDL/qcbSti/jYZwRIL9e2PgPlRGcCrhchQ+LRQffy8iHYfy471eo7
HPjePW4B0ZfOpnRkiN71OkUe7EQzR0nAoxv4MyGRZvkNujfHy+Mj8bYBXO3rQLNfQ+4xv24pol3B
RT60hNMjFGLKqS+ZRB8dKxgabU6GdYg6omJeWA0ULRNvg6xG0yCS1PKZmFXYG9maDauZ4Ja1Lr8/
97ECZtGe9KcHD+XWofQv+Eh4TKHmraDV0vePkiZNJt2OrQCEKQonuF7knC96IKeYlT5TKYDARkQ9
aC3pLGzP6vR/+w9GYeph+vNPjaQ50diBbGoj4Rc9MqDjedDW8qn50ycg9qDKocIPmnJP7T7KOKMx
Q1dqZrcKE/7BDVReECfKcsXEDhwlolqQzO4WJw53/kErjMzBVMZB9aeHubTGHQE22hlaxVwY4UF3
HUa0MgA2IEnuHsKf3vGvOz0XPUJpcVxjzNrbF6Iys6xVJk887BbSxA8gN5Ta5jLsHYossWYZObwy
4HzRO8wuCEIasDtmiJRBa74Lo/85h3RjGe11tOttlUnQTltker2SJwCEP1R4t26OG+G+pmCb17QA
mWOMW0VsvRGwS9PlGrh+NS9aG4BqlToBY0MGard99gSliDqcPDalmqQXQRej7QHGP2Sfm6zvpp8B
5kbSTvH07Zi+pUOZfHY8IZ2UOG5q8Eo2F3spWIwrTZvc7xJ0ygu9y4dF3N5IimJ7ATyF0IEln6yi
+tvVUQgwwOnC8p/LwcBEJaYtJqMqoujMjcPCG51axCvfvsdjwdgFl6k8aUBSk/UfymfqYvAaOjPH
6J5PU0uOLlR1yld5LpCauirL/S7gDY7USOwz3byxEEw3o8fN6uKGFbmjueGOm7tUb/fwUoyuYfwU
zoTtztGYDXow3fFatSnHKe5LpRvuSJAg5rwC+ybZBazo2ZFOQk1NWO/bcFu0u0aNvVKAYzJiZ+Co
Lgc9hosCP739BtYrV16M8XBjHhmf7KLWkLjJnXPcAoQZbLLl6g/gpida/e5gzTqnKGAdF6TqTOI6
jXA5n8k6eJkx8nWSb7fr5N1IGCcpC4fRCiHDAprb2ikxudzcD2sdttCVmq2SZ5OiDQ3uhfWjvzrU
ohlaiIdQL5YkXm3+jG0cMOXCpE7XyzkkJbnfedklUIhxTYdUJmIvrSMofb3C6+JRurWABwJS/XQ3
a2ff+d/Ux2QwnbKvK2euPMD0fmBH1glpCJYxpaxDV9ib3HQQM0DbQBr4uE6i2ne/kISwb8VexW11
/yKMcoTWx3E3w5h4HbL5lVEGa6uGe21kc1DrOwB6pY75E3mvtfPuewTBR8j+Zt+H/RLb0SdCoFGv
r4DDM0ElnmlyC6s9rYZqgQPHrM94bl9BUgD2i8GJhC6MIY1Mb6CzpkfhkvNeUKNxoDpif5X79/HN
yq/KLvwHe3DYGfY+Ntnv8lH/VTY3Mm9pBDqLMeFVzJXkqc6snc2bSj57Dh28PujSQCnfQRU3OJ5g
ruSbd9MyLzEdGrGVnVF2wPuZ6x5LrT+3cadn29McpTQJ/aTdvYCNDjykClCP0E3RrsnmbhtcBGNl
EcQTPHkViAP7VF/C7U5ITOMODWvbmWuNfg6+lQumD6OpXUFG1OdURpfJiBbLbsqehyUCEfjelYvy
kLJNohOAFa/HDpWctO1aqI9IlOd1ke6UGxCrDvXoGNlHbB0Q7IJaH/Y0eyTu94aCiz9gWB29ADal
7U8ygH9iT9kSTb3kGP5YWO57O9mwKMGp87KgDspAyuoe0wRge+IGxBu6RzTBhJjBmOX0xPt7HEZ6
iUJbRm/956Dv7O8GrnQA5po/5uJ/8YmQrs2C6t7wk2B7hRHIBzPxvuWRz7/2XC7oukCnvemfjy36
fFVT4+cQ5iS6IFU659G4qX7A2MELSRtOltho3rQon2cBSBkF5T1yjuqENjqd82R9Qqa8jHSaCguE
Lli5r/+NVyzLoC2+YsAB22nx1gPm9CJFlW0usK6TYg4X6g0eEwmaM76SywBXlnx4kWqrqKzjBxPl
gFzvRVItaRpswCOkVAryIlY/3ed90fzZr11xTUgD9zs2/ovePDUO3VeysCGIKBh22fKOl9X26+bq
l03zgehtdZMySjdl/fnLQebRTcE5zll3ASliLedoZ+7Y7Kg6PXUZ3VPZN5hhG9qzE8JmbhisrH92
SUoS+8nS8Q1VE8d60oiMCW8qVtbz0AZ9hKnZ2KZ3zGzHCMrmlJdjrGOYX4wSLiHqnJ3B6z1b43xH
Z84BCuCYZM9105HG+nW4vb5drQzejwsGz0XSOOQw7JwhBY1LymFgDm2dhACcKuqDtEVKIDs0wtc2
LoQh3FKAtElqRLxsYs01doz57PyzvpJ0fN7dn3sG6EsDIKkkcA/RcnzWV2zBvotSrcmiVhy1iSJN
eYMLFY+mn60EKpW18xEbMW+3J/ds2RbmK1DLG1WhJFz2kFdaRirhfz0uk3ZJcdr+Bwkfxp4GgOrv
SisRHGqa5Ho800eGE+VigyhHBbn4Ix88wvFYG7BTgRYH8v//VHOtfLVQArmZC/Wgwie0WEDHUTrZ
XtVC6mCpOPsWRivJ2KB9UBNfStXwg8QoEUywapgpR8i9ZCjm9yNBWTKy1aSrY44ild+y8KNZjlbd
DAkflfg7BW5Ta+rax5FBKfetIZeLyHNUXs2FlZQpuzw+J0/S5fpRRuQMLhO8kQonhSM+/pdwJm2Z
rQfNqPNNtO4LKJHZk++tcN1wd8m7FnPigVJ/n3AZ7YoyBIUI/4e5+OrXTGr5GaXFVE+fbTbCOJIR
Wn+Mq5K77Ol5bYX71D8avOkJqloCnAEZSFw6R3evs3j6KxAd+McT+qpCUbMSsrykh/JmqAR9VLLZ
lxH5kuAfixD0QN2JErr/H0InSjAs8y/kzIRudxdi1SWkE8/gUF2NC5QzxAQ/1UnPVZogeSWPmtuh
dHuRBHhu+xXIpPdHs7Dl9h7J27B2cmFkjboL8/qSC17EwnP8BvproLOjZ8mBILHCPJCdZbupbIpd
vpo6jDDPVdl/a2DjRBS2X7O42u7hgYy5nnEGnz9iPqa3cTSsio1ebSXrKOtgEVEVn5LikAz6fDKN
LFQUUmh5z0inWp+PUZRkYfbsMAyLeUK2B7Q7xjKbpksGTfLBars21FWHKdTA4Gn+yZoeW82zycgE
0UhCeJrPOOULdCiEsjmcW0Nuxi/naJVRbqzk9QTIZwvTOGp9XFU+U3nkTaoBK18gvkft8ttfkHlp
Rq4hlDuYQt/Sj9nOxTWtY9ATc8uJ+I+G/FxgLgAjnnjgZV49h/DfztOWLOAO/cJ0oDxVY8vfzGP3
NU0MK/v8SZjhESdV/wY/6bzt38ePab0HQxPG5+BKOntJASDogIW0PGrbq2okoDzdrYN7VCxxDIxe
R9aOPUpuwq552GXyz3CiA/2FMafyR5VyJmpE64rVJtOd3BFGlKYYwa+CFZWGhgASx8H75NJeNq3w
pj+7T9N2J9V5YwmLD3SvbjSLGavBwozCQpr86pBHLiw0R7Rk5njcflcg1OYplymnC06jf8BB5zbe
qZP6744HC6K12r+BecLVXRMtVJcS1KJWPQYkN24Ajinhi3mY5OpknjkNactv3XRE4sbT36WqXe1w
vOAsNV2ibFBEibC8/YriR9BagEaWiQVgLsdN7wDEuhm9igAkmjF/cWoJqGtYk+46n4KWOHjhSq4K
0d4aVfN4wuTUuOubMikj3mGAXh/fx/drHnuE1Ebvqu5ypnW6gGa4+LFPoxU96fbm4xDOAg/uLiu2
2m+6MahZN7SqPEpjuB9sH2a2i83KArUX+qoRR5ajTkYl7CLQQRUhgL3ayb3HHAkTkL3IetG56x2Y
eVFzHn/P5ejQ6h0LaFV4wjxkrtl2OtefiV+lPouP5p7/JhBidFMz5GPpXkgYRemKrIPoyMuzC6Eb
iIELW9suz1uvlR4d2Cafi4QRdqggnPnpGk+REXmZrKHkrF4Apx4ypZDB8LmGMveG1WuU7t4m/O4R
RQ1fjY3mWGHTv3tGSaNBEd//Sx+c+5YuXvP660PzhzWawmnuO6VRhRgCcx+dCfeH2e8/qgBGW+TR
jmsEW5sp53M3RalSeJK1fTkVSmT8TtW2md8VwNn+XQD4reuucmDvS7PSkQ72sRn4kWp82D82fhYq
/nUW9HyuSQy2q4kmPYRvr3NtfwnXs8Jq+RjZ4ma8vBfOYVXqSlUHztZ3O1sLkpNgp+sWe+5Zl6pN
3VgR9pjdBgADof6R7NIsPX5xx+SmqJnqStN/4r1BCawe20K1PInVqt5vDTaNN64CQ3/qGHz9pX2d
vbqYab3g8rb0w51HPAiAzldoCseW40g+VGHV2/weR/WoDjFc4o3ENwU4/mTXU87mFcmcju9Bce0M
5lkSNXbQHRLUzveZN693q7LraHNx9g8O0YvuR2pvJVSfSFsfkduelWkZCjDIHPuMXZjqjx4meaVP
/P4VzIetlPbsZ2MO37070QffA7OnMZkFERcyMOJdgXNNBsL5dGuiDvVv8UprqcVNFXLJpiJ3sg2Z
kqUFjbjwkRb8xtHKCYSzvDOGwyhEvu1AN6LxLSCURju1R1rScCamkHQhaZFNguQaQsWCYQkLzxYx
udclBBrOIQ8vOrzvRDsHAZSmhksNJj9Mqf+UTPj0rLlwSD01NNqLqN5qxsNBsOAlyL67jsFhMAGt
YZiiPZ14+y+OZgbEsD8wtDvWVm/N7Yw06okBqmCrAgLiyCKs237fT7Sk/2dIwhq/Vz8hP1PJDo8g
XhW7Fet/SE2tLapksbHEg5SABQ1oF3rb1mVDxVImKaaR94gi98Yo+gaBilvoDTP5UnS/YxbJ86Cj
1ZvbXwnXmyAwtv8Cwfe7+s3w1Fr1eJR0mFvvef6uCsPEV7A8jrxukEEOW4csKJCTxZweKpk8Bp3L
VpQmdc5SK9w0xQvHgpGhyKURFbC7fYIgh08OaAY/sPwxM32xfZPUFiLfQ35ffMdg9Z0YC/AVDOkN
WWTSZfBt0GnOxV7/Rrlc1cyw+sOO8XdNc/0HdrW8lX9zKmrGu/G01HfUUMqSOWkjkY/aV6HPLFS4
+hn40SYLgoGO4p26+gBy5skeLdDbKyz7wLCmvAw3mrJpUj1FG8T/7ZLeaKnOCL1y52XOfpQtVDod
g7znQ0Db0XoYIyh9l+rj40U/WrxuU6t6lFJ4Fk0aryhP6L3Jx0DtlYC53yn0Sg8zbmkLC+bXOrpJ
TOeihaGiazRlmu8u2n//t3KyPfKP1bzhXLAtPLjg3+VCPTTsSVbwoZChju4gkQEy9HNjaRYaMRzy
4jTaUptJL6wPCErbRrhFBxNObuI1dfHErel2WF0V5ol0sDlrLQizLGdnpu9eghRldrXreThkEmBO
za88h0DIzqEXyXF1I7YRZniEG2j+mKNEKhX7zFVycvZah+hQEzXNKoGqOn8EtrlSCgvb4zbR8tAW
AchFI098PFYt1EieRns1t9LpoTTWlCXfy+1mVXCpy2m7BiEFs/mJMQzHiqGQ2Nxp2NaH9IafwPUL
rMlOXvnKQCU+Qc2YdSGi7fn/EBTUP6jI/8xH0eaw4NxZtgqAkYx9rMvb499krckQsA65DK+Kuix4
rXX1tea8M2OZhYD9RI9bfSZQwihoDnhtUsMhaUU4GEYVL3NTlorAW3jFMloPGA5HQ4SoaSvW4dYS
KICd+5kGjE4/JEHvNVF3IE9reUsA9HwxYjoVq0bD+n8pMMvF/Lzd+mWwNRboLniNGRwy166ZG5nv
BSEyAGKKAaWvktE4OGs/PZRGdz7pYlW9FcV/TYBZ0WyQdy3m8QkakS5gPV5HI3FayFf09tPLZYmb
i1voS+NQTH+iMiIj3xmO8rfBw9KY9rGmJEh6lkVj5a1g+ZW0lM5ov19mEGNBEoc6ghrBM8iuITv1
ox96hc0yLKb7CnjCUTvMiJiByEphs9b17YF695o/HgGUVboJG/ns0B7KB/1FJXPs8bvDU8C3yoi2
WLnOU10W4yVYncQalcG4LoeNkL/tTjTfkT4aZwEZuzeTjm8GhZ0XA8xq6q5qESY1hcI2ThainYrJ
v0Z3y5mwkDUy/jWwffNkdMyPUcA4a7y6HIO1flobw2N2rGOxJsV26LvsFB0rSAlnNePI3TeapFov
HR2PBceB2g2gddMtLagL7Hs7ZtWogpXN12Rfmbgl86l3JQLRI/vOHBawVvB6rA/YlVI/FH+8c2bX
RTHY2O3sudIa896Q8gAN5bJLdGJpFW9+enP3l7FQ3vTGA5EgQDMc9+KQVmkygHmtrVCrjk2b2YkR
E8nh66ajjyDzJqv/OVABQrCiS38yJ4HnenQ5QH6mr7pGP4eYTOSE+uFdYlyo6SsVgEQKXw+8DKiU
Usv1wyokG8ny56L4cWO76pW+bjxAbX501g5BP3uZ2nNjfvJ5xpQyKNNutrDMozvFyFnBv9njrkBv
EdTeZgDeAg6+TS9HtV6JKXRfWin4uNZSRIJf+oaD0yHUMurxlHHR99Uut0kWhHZbJtGGrmd3omL6
NIkn2PDxBo4UAJ3YEC6I9iPN/ongx05TcFJ/SUi1L+eiXjbSXfbcnUaT9vuKs37JNEDmqNmUy0Y5
saQPUVjeye0NlUO7Fjiv/lZEQnwwsSU6/1dzrvWMnWnmHPehqqaBjXCcNbXCDqWdHStcIaxbdnda
QoDkCn1m78xssPV7t9M8MugFlKQXwwXsf5O+kS4mhmAHIzx7BdOoM6IH/JsWpT5IKb4nKL40cSvs
KFfRBpSiIKfC9CBHl3uuWUowM4mUVULABP1CJT4VSt1D5VFw3ujs4IswnW8DwTCDkGkLxrA0jfeK
VUpD9fQk10m7lMt7R1yFVzaPo2PnXgVw3kG1NYLKekar8AiRqDuk9cw3EgkXmZBVy7V8+EduZKd7
ncKSg7st2l6SKjuETToAbuIAnPZPKYSE7Pg+IyjUjHJxuBub6S8dmkx5pOzni2ldFIpzeYwW9cF4
uM+xUgdpTdtzFgBDcZeKU/JSIOagGJLNbnDkjW/hXgcz8JFDtgu5zrWFSYl65HSF9PCj+ltwdKAl
UdjJzvs+9mM8JeMmR8GJo9dh+++U8/fyLc7b6xPgUvz0iDTM/8C/FkSiZwEQpe45+EAf1EAuDhrb
Z8XlWV9APmIb+EEEOQj9QBwUqyE2z0mP/C55uZM9B2ZRwAC1o0O5L86nWDNx8L24Nve13CW1MG4q
WqMep4OUMdUOR2PzEHBqCh83m/+3abJQUe8dBaD50ZF9Fbioxxm0RdUqhl64l1AW8CMqfA18ddTn
oaGr2RW/zvzyWYe9U1WGOR2aAeIvzWPwvtocJPKKInsISsZgQVJjjdfxvGiEFrPk9ajT1FoCeMdY
TYRcnmIXkayNt/de28IZw+gJjdTITEHYwh6A3h3rM2ta4l2jTuAqQjqjATdRXGvvTeox9GpsIAnU
vV0JyvmSCLZYh7dI3MqruZ/V7/PJvV4KZlbtkj+G/3zVZ1By9uy7YMzvLGDJz9sh4NL7VssYjUNc
kPX+L2f7szlMgdPq7FjUbAvp3Xvi3Ffi8L162bDh0w6mZwJ3Aow9OHGlfn9ga9iIvoBWvsocjepA
m/Vg4JyvmrrxhyGl5Lgn3SIBtj2tdkTlhq50PCDgAJtF9BRGqPuDyhqr+0vzFss1IkxNRmBdvxsj
zayUImi6R7slYaGU9RRQOOSBrQvDZEHYCC3lT2aFWidAmybWfrhdBaoRBv8qmTfKx6ANdpN8QOma
n7IZynNxV0rPdPO+8ETteulLF2wXnQ5KEwSNPgoHp+aR2XJXe7OtzYo+BprNCQTCmtRMt42hXhk6
TqU/9lSi0NM2TVAoxu9AOBt15S0njWzeZ3I8FoIlBqB82Tiul1HjcHkCkUPXA0GpTklPlu1cuspa
IO8gLYB+WyUHJeKpW7NbXGiVzY9YGhmGdVBTkYnkxMDbZo5gvgxr1aCpd6AV4SqTQeiztNs0q0iF
kdqvPNLr7j4FlntPBlOV+rMEadpWV98iBDqwocNmwm1duHEs2yqVjhchYV+6/WNMUdtfDGPS7EFY
xIsGcNMtD1UlTuOIcAMck9zRS/MCHQWMQa7vECKzKj/MoQR/KnS3Ok/aziG6yNF2nFMVALLty+n7
XU5T/RbMYBq2J0dsfp3t1arE6dnDxWMmAaZmc11JYddkJG9zvdqXIHong9/U6nXvzx9us9VDUSh8
2TQrQLTd9zW/8Gt1xIkGMvAr0JbAeGH6SoVHRXkNLO4VTvx6KLbd3Fi+F6jRsn00FCwiKiSxPMmd
gAfSGVMjBvj4p/17Pezg+Svp7NVxOIquxGa5Byfo+RSfeqMchwzWZZC/ueb2SS78IJDdKXdupzq+
zAWJ2H8kHuXMu6tfHwc/A/VUtE94JEfjGzFoJxfyIPR9VpraQnYCMo53+8xUPiLBL6pjcun9rzp7
GgM5awq4WanT/auGQUDCoKxfQh8QzKErk4qfIypEocAoxyPsyK13pWTrFbgH4AEDUAMwq4IBsndO
FbtNEN/sXuqjUEHtabWbWzGbnjDoGly9/ZI+HqawScDkgN35Pww0lUspSCZqFidRg2wSjb1R2H0I
KFCIAkiBqcGuLGupuFl9IolcwvD+er5m7QukjYxossk3I3vTw0IcDcmZ4nReC+F77JfW/qWUDPLE
qNYEtzxvUFbDgoxL0sFyYntDWRfKPy7Sf5cZJWBNsSapXzUCYLFD9oSLhODbUPPBYCNAIn6sOzQ4
Ax117GJqmGxnKu98jBxDOnwga6H1ORQZjdIQmu/3+jtZVdLcCgGzB2SwxoHADtzWdPvqqOYybou3
tPKDUb9llZ6x1XEZnOvRVFTLBS1ycfAtMP/o02wm34+st5dky9PBvgxrgZZl7EFMI0y/5OfMgAyE
AqlsDWpP7qswVSGzNniKV3egk6adFQsIHdNFDz4QOsM1Y99f9GXyubVg1ySoPaVWunb+ACGQgBSh
L4R/vCLKoZJKsLOiO+YBJbjlW+VsQclqlCdZuS6tu9rc5O/yHpUVRHlEqNYgJbCelNtsJetZCrrT
SYwZea1T/+2VjiUvObVsKWN7dV1h/PouD8OMtAZZVrRwuTicNQCMZWjbtpdefwNuOTiQvHOjl9aM
JjZIMV3ZkVO0z5o9Fc0t5h08xFPLlkTte+HEKjbW2oXcpzlQDuRAYR/LWzKkjkZw/Bd62b4WxeuE
NKrgaZ1DqBceRhloFy7d1HXVkJTXlCMazbLZODHTMGEUqgPFJCicEUd4orSJtbqa3+dnKGnst2oV
2nXRG95Vcf9fykUBlrRQnvrTWgxo/s4eA/YSwLmzJZx2mGW2ol872JpZFjWx9g5kjIxoFR9EYv6D
9LSl3Jw6y81tnXzmK/CWSviKRvbktr1CLWYJ15SHZehC7W+Pi1FkJ5VaNoyhntOXa3TxoFDDn7HG
ngDJawMApjq63dLQqx9wwDE5l2Fa6VYXDTrv40nWR7H3O7vxy0Tp2O9gfqCIulN3B3vRv5KQhkJ9
l7cfaNrirGcJs9uiYwKsiBU9bDwvLNg/WpnUlh4He/ZwmoKqrBv+tTNVCtEtdgk3OZJH80/+qJA2
55aQ13MCgOU45y+u28ogi+rc/hCDyUZhhKQaS2RkmVNe10pQ32ery4/RdL5hRH7XA2nZapbRuFoP
nqf83SuVLkuib+hK6dCpPI//SL87JLud32FMSTbLynK9JgF9jMU1JmsDBiR7CxBszop0hOFyZooD
gTSPGj1hYqo3hrnZDAsmZH9/W7AyLYdXHf+Yd55FAhLE2JikvAlc2+VXTwp8VFm68qIHGq9LA0tF
j9EkXXnH2izQTz0WuxQcL+n4bbJBiHFi8yUYQ5ixBduMW9QerAPqUqYKYae9mzF7VppaNEUL2JRa
87PhTPaY2D8zHSwMe6BF5lrGZpEA39QUPL/DShaIbZE4BOzJWxAEo1pxJmv/s0a7UIq0Hak5nuG1
biWr92CY2bb/CtUhAnPAYpt2cOXJn/Ee7gwFziQZdzaDByx2TWAvMoiVwvYhCVbAk7ZIm1OG1LjN
dh0F3hoIG8cGKsLr63ytRtI2YL24UAq7O+q+d5auSYpWdeLEVIjYgd2iF3iR8/0dDrBamYbK5QSg
kqAFlJ0BgVbJixr3QEMBHT/CtAu5xDnDXjPpovEOM7/QX7nR1Ct65KIfK3ROpW/Rg5vJdYl1/21r
ofRN1qFZ/Ge07MxJFrhe8NlZEgZ5C8nEu/mIGAh1QJ1KO7N06W1okFqSkm46gjzr5AFuU1qFZAJv
2c7QJBnx6KXKA8w8JTjN2hdDrM4JwT0M6crcRike8JkWkMAUE2qyHgdW2XAekiTe5oDSiAoQWNW5
7XMkf/mSVY7r9vzDtYDEK7bf+9w+Et+co2nflwh0fvQ1HCkzA3ZpGDJLrLk0in2MGqnYM1hqeZ/8
nr3Q0C/5SwflXFG/yqlNlkkDxZGDcQxbm0eR3URi/Sw/oKOcCmWwW9HegQ8EE7bQCWo3AlM4+DWv
R8xyEU6VZYt6xbFaMDKovNd4BN9++W06PALGA5MaftWQPLHLR5OK5oXR0oVMhwKEvTD6HOTTiPsw
Ljvz3Ts1QaAYahhcpynfk4J7ukDlAUTL459QFTcxOT+mHx4rrBfVyBWzCWwfukvHziaVn0NNsSWj
QEtl1DNlnsnACJmYhBi0/TUODhceyBxVqXm2CT3n5OV7yQJE7cO2h2HbBHmiuwVIXOU3MhPsfY53
USIsydWGKobP9rfhBA/1BstO1BVYd4gaHku3+n4HT9nOiMnAyVAH3cZ2TfaRrxGUIJ+IIxxJB5Cu
PtFWvW9V8j+gT5oGcIhkwyT6oqXm1T5QYLIJuPzRGvL8ajNh7pBUkBMv15nN4iknu5lhNepomU69
1e8rNKRuA/OLzLahDsWT10U5SgHpokxPXaCYcJyi6Nke6lgVyUQDmjXpoedM3L2+KMkeGtuFiHae
xSxXIhZ+ejphionC7/tHb1uKjecKyeVFR6PJaqJrw55gysZtb4eJjI4wpOJEFne34O2s23zurRCf
TnWXrsKypqo5Mid7CHkoits29OaJf5M02mWvmaezpJX2NgxWjkT4ecTHTq+10MoDbyyuHIfUDHBo
vTVRa6RLsnyGGZRUSefmE4h7/l1ypIqR4YxOZDND8m82xktCB1OWqeIhZDHQYsPIeJ5/u54wdSyl
UP4AysGkM2s1llnjJuzJ/DR32Np9tfrpJwfTT8U5hPdAp7uALvVX13P0h3U0IvxSaQys5Cz9SsVg
1buKjD4JvEe4dy4T7bb7hT5dfZjWZl0XNxe95wB/N/EYXmA5qvgLxfrtOLUbsKSBiKRKzmuoVP67
rvDJyA88qzg+P0Y5kEAQ8PaGU97hQncYxZ+MYg0xLXUBNJS+nzfELYI31MzZAUOYgx+DdeZWt2AO
6ODI4h4d8eOFFiqcCYpLhE/jeM/WDvLbmdmiftdAElxV0SUERYSPe/PpVEseKiLKPxiLIs/2qW/D
BL4ekzvu4jq3lsRFYtzO1xOa3sydLNpGNXZ+hlgfAn5mhpaJrjPunopUq8stD+6Z2xpF25yDaYPn
6oKyK60FofL4MJAjg970xrpKFvPX5vlHR5Tj4M3043lb7tfGMmD+HOerNPp9kf56xlvxFIq5N3z9
AURjZcCmqG52DgdiQR2c28j0hTm90jSPlh4hTQeiOBojIehuEiZbSMVLyRc8eGiFcT/uU2y0RGXU
tdH+4Tr211hhFy1KoyHspHLlwGTr0uygtj+0uJ8t/+Xl6x/BgdvB8XsXNPp+iQ5ucJVF11b72FSb
aRZ8oqCqaiEI6Ap79gHfDqCvSOJGtSPpko/AHkLl0c5YQPZu0r0Es/ffEMcI4NPzb633M3e9QxM0
qK49f+fnaeqA4Pw6Ikp44aW/esVbFZZR3ylVHTq0i9xKSaaiQxUgBUt1mxjyErBp4swWWV4MKJvK
MPCG4s8611WkBqEu/upNGEFmVdtZrCzx4/rWA4Xdp0vP0258YXnzp9DsYYuWihIm4tKw6k/cdACy
K6y7FI5OPA48ZT9pEiQSx6GmjP9CdhpTwjZCVa9QpbkkLDPYfCi8dHrxERjcbGu2HOuN1UJB/Lw6
pb3jVxMP8eK7vfCBh5wnWDtFORtN0dnZPtbcAGX9/zt4uhhMFTWY3TjFmetQ2iHIopqTtkCj5YNA
zdU6muhG/KdYI7ubxru2kYEKcGGj05JVzhe3wlVk4KxIFlVKglYCJ9tAM2ftKZp41Xk34BUllN6l
ZBc4h7N1KyYXeksRR4ey5TKWFplY3kFU4ovgs190ybX5iJB3/qDdNkGazIL0ZXiX2f5guaR0VzaL
fQhKFfCyYbrdvq8XLR9f+eQvglWtFxDOFbbMSCcKF5Uk4P1ZYK4jwDRu3iZpCeB/vy+QYBDXqeEQ
DVzISQK//PJ2BOlBPWGgT8iej7p1ugUnFRjkw1VwQH7EEDNCFRTpaE3FcMKNog9Yo37LeWI5QEhn
9c+G/e0Xkq51Kkp4VcWfPRohK9A8/0W+f6J3Da0MlD+GEHYiqaAvNwEzB75/S7w1yAQBUE3URR/c
nhXdZ3UllU4eYWtVMrajZBtTdKFDph7MrVTeM5IQVsYtmbacW1xyWbbbAuWlU0uNR1FjLvDdklp2
4sHt5etCzaUkD5V06fPgqPwSRYpkO6Uu/IhHY8T5tQgyQl0/igoeHR8Vpk9kT8sW83hCniOhrFxN
oxNzv0VG6exQ74LSPfXQ63YL3F1NllFeL6nB7B4gub4imkZ/pZzfS0hDaCVxYRrqE/BVhUvPACrp
V1BgNWofKHmCXxDRbn4sy3ptUKKxbXXETXByCQfTjUdiO2n5HQ6yGGMohC8v5t23cu/AZAgVWKMJ
lAMkOYkLIvveB57eaYt7USZySgj32uHlUD1aOjStJmqZjYI9tvbkw0lshB2Nn1kGtINAOvocbDxn
aNRrWUN5B72dXb8JSSpFq95mwbbinj9AhtSX7FDVbfkSwkFU3ayVIYtSmSCJDuJ3M+s2Ywyh90+z
B7F0KPco0VsvJAYY6Z3mQmF6cF/vjgdDSqR2d7Ck1NgN9OMbKPUR2I8YpKGW3qEZTF4ufUMVg03l
KgUuqNUvBSnJK/HL/3YHkfrNyMlz1xVsieZ5fVVtznb/VpWezJynIhGS/UFXXhNQqT+NBsImyvwP
l0JwIRwnP8MVayyq/HufH69DPHsmkdXo08JCssOGC+70ebU4pEbYIfzYeyk6Spggimf8ZmPPI14y
8srRLhxcDp0mf/aP/7Dxd91E5B2KicaiM/35mgiYR2dK2P7W6+BuJZ82k5hLOyPTUbiW8Mk4c8nZ
JG6rc9EGhsD5qWbbHGvtnoUfqWuIOAnOwznUKs/RNlXxYtSnM8Ku380R+0DfFGq++oLvwHhWaHM/
9JQIJGSRvvmypbmmGgBY+lpslk7rYwqpLFd9on7CgdluKSscxuzvdZjSN0WuehZsV6jx3aLOJ3A+
H9pkRRchBPlkoFesigb1CWO+qD7e3/7GoRXTrdsTMNDXKrTtMxK0MB0H0uF/996+iPdNGpz6lnDW
ErnP51/dar7JybKe/8dNDlq89ITA0rcJiRJ7O2iiBKN/uZdU7EdZd18Zg4DWROpwLQSvEIT1bRtO
YuQrA4kKtsVO5pREF3U2X7NvmG+i5OUoahbPYYaXx3+sVTdtac9+dJb9oT3dGR2k43mWaM2S0LWf
jMX1ap33I2BSaFZ9aHY50dbaE76eSbVd3dez1m/OECeapQoWlvrK/a7RBAT9cWtZcLRcuNLykZOr
PoJqt5Ti0G/Iz7+SrQm5dKgboSL2+B1SXsBVFVYtHRjLaDndgkHcPNt5msP/E/vFmJJGMjJaGLY8
9aup+NGCp8nCF/YhV9K8ldqZYt+38rAN1+/zqGidJk+KSd0RUtroXCqfUJyiExK+pNU7vpbtAuaM
3ALu7Dknhjyvmt1GNGUn038ikso/+C4sdPWTC9hAHTgUrzfqB8ZP8aV3NC0ek9gd7VKRp7y5pSLB
fEnV+rV+Y14D3S7t60QZgeUMd7kbSJ3dB1iSIyiuxKasVRGpbAbTUfigXB0uZdhBiUWh/Kxtku1t
O8dWSVTwHp/7azytnpJD1GXFVi4C0sRjBUOMmycuWGbfBLKm3yihjytxY5iXcHF/7orPXmZ8pC9H
wICM+Kppz4NCH5I+Yhoi98KcHXiBT3ixgoMk5Eoew/WwB0iNVqeFJ1ILhhi/cB2WyFer6PDQJsu/
liu9a5GDBQUKbtkIfP8qmuSm/bg8ufRhnPwOTE2GtJRftNmkvBz/icCzFGqOUnwr+uTMFODUOSzH
bPoGdfCZnklIavu4BRA+GJdaBrFoZdXVjswasw9P9snZUOD6TmmDQdyrCvhCGGMdIhDb2Y9qprRf
K+pxBqwKqwAswXhI6FMs/oWRziSvohpOKqZ9wmFlpDLPKqTv/D913qfjXRaZej3AF7ELIyJT3Du1
RumvCvHwi7eeh/jiOlvSH3YYabI11hgqaUBiCaoins1S12D6oVs4ZGumhzyhsgcNYhD1mO1UZEwg
zJ9vkArGUKch7UmjtCYox/EOGcLhKpqDhBaeJtYoFMJleTDM25E4wUPcNIxpApgvtYljeH3AFm9z
fuha1TZWSEPBVt+WfWuYu04N7cqmRSITb5v5PYReAAfn4ZJKuj5UxxNaD3LH2TB8dDn7/dmolFOB
y0mN7kJXjCxtP820wt9z2RtRIG79R/2ZoqOpE1Rw3POY/khVRN8I6eOlPa0H0q19DN/Oo2X9sN37
yVjdgjhiNFue3GLHxYXqP0ZWkTikcr6GRtjzhZD86opOc6unrsCIFXheMVasnVU6Fm+N6Rb//Zp2
JNNagzYOmrgMWLSJLtJjIa/6ttdqCVUepHiWsSYAYy+joIBpdFIWCYV7wYmT44Ow5MQlqbwxd4S0
NbkfNfzZsEDsBZ/NM/ZesEcVTrHejC6uIUti5Eh5LQslqQdWctBEkZ0oHzqGhwo1ATge+kDrn8bA
5lbhHoGaBxqXVfZwWofw2QGs+c0pHhaj8Vc3VHlaWc330UJan1tTDOWJO1P/EoyszMHQ6Rwr+7Qv
LausaGxHDcle+2gMUZZdfeKGkS3VXhAk7yzCfGA0uHCtEmcE2fp0TX80Q/x6pS34abU6ZIC7ZDmd
IAzf6u63ESM7rl9P9muN7UX5Q9tBF5EAQEGelhStkwantiqPslKhmBZnNILkWe5oVJdAhTCVQLoG
tnd0nDv+vo5g3nQEGFe9aAiOS7/C1ufh2qBL0+Pz11p6Fe0CYk+bGQ9LaPmBiFspqbHYNS9rWn07
VcVNdkW30i3WZSQjoMt4H8Wq711kAi848qfWFfF+LFQifTt4HJQC+NCcugyrP3fi0SwT61h8cL7R
wSEugYDyoQN8TFgXLbozcbmlYDvWzSipOza1O9nixiojUJplwP86GdK4lqMVdzUKxcqI/xfsZ/aH
xlkjEp7bp5AtaB1vWrikD72GpOhAdHDm0uiP26GmHN+R8WzDnlQNvgbpi+c2Qa8gNpzfN91udO2H
1AUF3Ps9d0Hwq44NpRD3wqdRFTMkmc0tuqaKnCaJXtFDqX956QcHeLcl3yNRgBcX+SCld7YLrrem
2V8U6L7P5wVsZzgFMTFM0tPl1HCbZg5pvGVJJqAWaT6WrHG23NsBUTXn38qG63897Moi4J5D0bQ9
GBl2jQEFPB2nOPjj0CYkEKh2OXVdzlKBVuJ5DWzFGGCMLDeBxlutribsLRsJ7aW/ps638szTCWjw
xHSJ34SULFZfgQNBo7eYxS1BnOo3GwWVeOvTB/xKq4ojoNBuXK/B7gtM8sKcWoyiSoo7ye4pe3Ch
dxW/wWrh+6yp5dZNUG2sUOGBKx5QFqKBFNIJytUFxG7LcrzbmxlNHQ+3HQpK4ReDYQZ0fTv7R1Cf
39ex4W2eB9IDb4mqLN3CcUgXUcadMJMM7wemp9ef4lieJyKOk6VYIvlA7SYkZON5tHLw2WI+/Xtu
eoqzm/lswt4rE4mhW44xMw9nKMCU6fqTGORkFPG0Ae0VYgg+UVkJyw4ydm5Ys7SwyJ0/g5PelE/w
e22fYNriX+oGrMuito91iJ6s0AMfkMk6Jf3awOi+2pJoxeSxjSzWmOzToChYdYQ9r03K0HggZqJV
yo0RHHAvXsEQnzaidExSu5NyZkpILaSL+OXwOi+uCrqVE36WIO9pDvpMaD8VY2LqP6y7by2ZQH3j
0yVhvp/m8KVPDeeSZbL2nivhopcxC7RCQ3j/lgQ5YIWSx4b54bh7cwnWOjBXEGtV6y9yvqi5nkXT
ifAidH+LJF7jeSdocCER88eI+zYb3RIKHBFsZxeNiRmISeOqH1HwD0rioPjlO5likfC+FRaMISO9
BUXTUT6TN6IEigwd0Od2fP93x3kBCI+Q/4FLIidp52QaMKTm+EAYqBHkinehzRXPJwQk19Vej6hZ
yiprvGgG1jRQn6wE5wn1hwLSQaywyjdwB91tM84XmkGuunIPxOlGHAyHCW1U+DDi6WLPANaJ4usw
lkQRoDU8lH86u0fhJYJK4NQ7rgg7CJK/bdCXZduHJqbmKG76Irki4QlMim5YHTwMVqN1CWqEpSwa
6jt/kKpTa9okU+Y5416U+H8G4Aigls6nfq6VgJRoc/NGTe2Hl2c6NUbGnZQakvAYCMIs8vSLpRyG
7aLfDzCAgrDka6df17bTOnUPtoHglEOr9uDt2WFhKpG1x28hBqj1T/5EwsRXmFhvCU/jiFCsqRjm
9FM/Po2U+/GsC9MoH9sJ9pe4HKZtt3JB0UuQJueX1RnTp5vKAbFf8Zdv9OkPre9J0HPnKUaCjviI
yHAvpbakTCgTDSz1wRNPTF/C4VLiuM5Tjlj5gsPhr8p9NYywmlsIM8VEaBgx+f+gqVhWGt/bozQX
91ykFqQY2hNnFoc9VcrQCWrp+SmqvAvi/b6pfwl6NHvcYNXj56GfHvEGSQVNiRMhW2OcwHeISoUm
BBPqg2UVk9+eQSYeul8AvLkmqT/5lb2msrZRBCvBm5J9lk9MxXw0PP31Yodgcz1IRyXYvdjzXxZZ
oUMk0sI1fivbIZJQO5fjtVLqp3YrV/YcRMbD8R+VH965pX1zKo8bkiU1sQMkNnpAL95tIRq5w0ig
pzK2oKFOY7ijI7fw24NImpRSEB85ome4ZdBcPrhx5jjyGUlXdpFcMYWmBehm9L0rXU90wDiHZd/V
90SAPS70mBp4dWA+iQMiZAIleGgor1cbnflpkEcIoJK83Vo7aMOfZn2KRuh7Rt4YR+n8A0nobmfn
9h9KIdsYPjNLjTR9zfMvsc3QepZFPUJEEYkXfDJlnzR3tjrhW8ZbRvHqUGulmv6CnWczIUUqnYEC
FZyfetlUtVgBBYlA7vOQ2UEhHLb/LnRLv7Tzm7uERSe5nXNJpErGvPkil4RGwufM0ge80rdNE5op
GfYCiq1tDJlvALr9CBRJ8rJWGBzCevn8SSb7tZmdk8s/ZPAeqVz+Cnw15RJHe8QpRzbmHC0ujwsK
ZNkk1o8mU9NbY19ii4nVhTknHeZGr9LRLrRxNgceekH2gP1YBGAOWPMsqF5eclLlDWY4F4lrMKoc
vHttlHIlFoBfMy3XUHkaXqcdDd5uZlg9E0KFJ0Ia9Eg9oKfjE0EHnDVZ9iP4A7UejVkdfxkqDnLq
/vIUtw2bZLW7OYVV14GeXbH/aigtiTzpnDpPQ1fWNaHYOtK33rI1L1/glbPnsVSL0ykiP/xZ+JWl
I7n1pMdo2qssBUW9UPjexmv7AA3P8Nx2vdMneUNj8TNUHIN2onHjl9NV390aS5zIngtbgDvdNpeK
K/cqEXrz0DJnqsz5VBrefDLnhG2Bk3IgtCA87j4Ghr57GBWC6KhST8HX7ri2S3PA57yvaLCAUC6O
4VjsrW1FBz7GYOvZ4e7S309FxDc7sGEEtZcwpH/ntS68cEginP8Px4v3Peo2jLg1IgoN3lZkOa4A
pofWaXiKYYr1TsklwSnI9BvfvfGPsVKMQcEFL9LXTPeHAlPdicN4c6gu1hSK8I6qO3kO0CbAjn/H
dwniRWnD37okjhaCTqsHgjnJ3xYhXK5s/JldDum6GP7MEsTYKmUKBfBc7blOWSzJzZw+Nv1TzGSM
f71x8F4JwH18EwuIKgtNAD+mdtjZyfTNCqdXRFRn/O6W88qu3IE7Gxn2sZwnxA966YH1j+MDG48U
WUavmd/Gua3VphektH77cghdQE4uTwC4npZMaR6SSJ/yKL1+BkzVDPHViTQVLEsJI+U88/sg2aPr
BgpcpXYXuaijpdfuTih/0h1kcMNDWPr7FaaUvMymebSxfIZzwcKU95bWpekrB+C2PLhcpxt0ucsW
WrcmeJuOWlatewbmMiXtLlXkdcSDp2xNw0ZS5ACApwKuowZpaVjNsTC+Pezf2WuXgRwr4E2lh+SF
K9eTC5NXDL1Qzqbs8fD74SvNZS53/AjpH0khdLrEeib0Zy8sjYGCzse1wC2dBF/GDB0hIqT/mJ9K
yUztN4c2aQNLFZaRIHw8y+ZyYeP0vTH4X87AV77d3hgjJ9KfV/AP+SBVh2+b+gRwwDijnORFflXR
tTvm5lis1fnHenxmWRRuVZ+Q8dDcbiHPvLh+QhD36keZTeqv9GFx0NLuYPMrQQBm2uVdd7TlUV2s
kArkbvqds0xT7f3s5cM45g9U7pWvbYaJI7urqQDu/ZZd77OPCbZbLAzgNtspxgWuLa35O3npGtP1
Rc0/4qHPJEbzB52NANKE491WzJ1aCx0H1aB2T8yxHV1XR0RyKPFfkk4znRUSD//S8IqbGvXk3YbZ
uHxzRx3RnsQVFT3I+Tct/m5BnWlDUS9yP9kfNr0olxezKTuk/iEn5S1iPDCMKooWYwxKd+kouUvn
odlj49BT3KPP9kaiM83ykuBjh6aSHwfcnCp9CvJ73fTklbBC2G4D4YDN2DvQRj77ikBePVaxwvxt
ul5GhtKSB48w+rg0RsIy4IUdh4Sn6+jPSCZ2ERblF5fBDlPKDMptw2GCEFRR6Qath4kLSvUkkHDF
0rehSkREv5poHiNtA9sU/S5Rgmt7UdOJNTd105ZPFI3xw/83NZ9uEhw0IGAa0tUUwbZntPgfsewu
HhobeW0gGCK0OFne2+tcaSihwWdtpgGcACUtYn9ddFxXDwIa/L8QLxkqvJ1uB8HYpW9f7HNff1SB
0kncykIXx8zKVre173Xa+g2hj5n/Zt31aJJSIT2rdKbzsU4DzgfPwAGpj7MhSs+K5DFb54JLkkwk
Ac+7+ofxKOryryn8CQCRV7CMSDa9XBBtFr1vwje9PIGcHmu2Jpfvgbt5+lOvPgDIPMXACmDr6+8S
4NRo0KMuUj5R2dHBnX64ZKU9oo0pokVaFXQVfbxMDh4KzeS62z0SSk4BjxI7WoJztp9y6j5MtljN
5RhkZRTNIdudf6qwRIqRrL8vLqwwLrv4gz9r+uTJB4ZCzmLuXrJxjfE2M4x69Bdbk+vumcIFYTpn
0cWPwSjRuT4qwAupoJ/jKSpP2q1bBUN6+KjVa9xUPIxPUbMeAICZ80EEwHZyyOAYUwxh+yL893Sn
N54llroY31Oxpi7VeDo6+isrlK3IUTvOr+UqoWWmGgTTFVCqJW1cICvGMRqwBY8elWUwDYr3Mbl4
q2q+ga4QcyOAHZuWerlhfzFRuwjDpOF/ln+G4yhNAxA8lcvADOlR0QNHmzqIg6EkWvL/6+USXY/E
ozKQ6ykQ9lwfAgJ39Gb605QGUOW4EFUCwAr5M39vmn06QyIE8BDiKiG88KO85B+6gaWsDA3yhCYi
HYy48XydYRDkR21VL5+MtEiQ4PFbe/NKo06CWPtrdLoM7sHxprjkZzhNNhcKXtip3LIsC6P59Drz
MXMIX85ApaCM7ipzOm2+hirk++0IyLeEkzQ8iVZSwvPM1SadX6FufI4osV2CLOIqMfhsezFw1pWM
l+BXd0BfSuE9kY8KTiet4kAp1COC3nXatC+rDrAqsqlQVJNFL9x8wid5XWAReeY2rAvDWh+mlpox
xTnAbzINAQlKrt44J2LY5dgPec6uGhEePIxL9YFyT2nwxE/LBMnZMTXEAA9mbi0Cn/WtzTi2grrZ
XMCqcSKtEQFyliJ/kN+o29dd/8+A5JvjwWqR4RdpEJZPfisuo3C5ET4bqhjoAXWT1//5S+zO3MZf
IqV3Dcf5Nlx8rS7SiiGTMPepcB4kKYaD5ReCu6PDKfM+gLQ0uO3udAiCAMrm8GcmRRZxM9EoRDX2
D9sOI/GfGl5QVwOiCiLYxmpdbWebTLibMfa6liuicSqQIt62lZIHS/ZHwb6gFYY9LcQd2zKcjO+1
E8qm1CZIzcvQ7+d50HaxWMstu0P1+RbsE9lzuU48FcWl4UWEnU4UUGjZbS4/39P7SvWg8n1sdmFJ
4qGLQ3JN97Aj+ZuJiPzpw76BAc0HtiMeUFBcnoDLUS1jv5JfADEBG/vVbrjRPpNaQzBq6xz2PsSK
0j5hV2hmQPwtyEGy/wuHqw12W/vQuntypWOvfizYlPmGow7/gDzvJY32kA5OmB7U8X2PC9lZN97F
Awad/vHjkZtvpYkLhSTTqclfJilcZsfGbvi20GPbgy+OBBZ616CdljnUFrMblZrUXJ7GPP/lITGi
qTb667+tKUZHrGEiOxA9vPD59ghP4VCzf1OKU8kfGctrB45Vysyjdf9YbwPoO5T9p7pzPbYOBrtH
MO85jbDOg+KLvRVACh8POi7uwudsFEGH8D597AWhSprNDl+aZscZO5yqN/jL29cGQs1TezHkGilM
hRVg/LJlTdz5s+rrUrAiOXTxxhJRH7SzIX+Ox1wAjspVoJdxkIzh3n3JZWykJlYxSDltWgrEuhra
MMQUSIbXNJWT/cRLE1xT6eZ0QFutu+T7DgJUSvVpk763bZUT1by9T25qKPyhNL3eOlpZ+yFk0m3K
158zFUYJx82nZ+gDqSymWOSGN3BAyMTIMeNv25pQtqUM+5ZPaVJU64bSIRskC/IzNwKJcqcwT0xj
+8H05dzfkUObyNDRt/yoI/o0ObCrv/W6/ddwhxki3oDgj20XhNsGKLqOYgOxjP+UNUx4xnAgErrr
r5u17l9knIgRjHgwHcvnM+ZijM/BsPAIcCZFtv8+wg6ybNkQ441NsPTOpScPYYcjSLGPZZsrjDMs
yX0ekPrpiiNdISLTDc2nPZYGVQ6/68//7s849RZJ9hE3qIQX2M5QLJWqgCdkryabSAaFDc2xw1Eu
61AL3DAXXVhmSln6gWWqMYNJ2lQec7pW2YYfooZARTeYdQ+//dyvL7pCDArnwvXpPCSn3SO+GHB6
hvUCEhdZ2MPRAwR70hjpgzUxV61H7oGnSQPa+tpmMNcDK4fjHmtRFuXJ5X04MFDbP9VViKU9x6Qd
YrJVZn1icyNTho6MRWYDZaCyBrEMk8OcLqWJx/4Itm72fqSpSbSkl7YZQi8rt5nj3mt0SaHH1qhL
Y+kzB4mqMx8CHkEIvPSOOWw3pFXd/iFrnIddJiIIG1WmSchjgLMHAzycuIc59KhqpxuqJdMscDXx
P1kXUviSdcCq1wKka4xMPpCN/sGMxbdxrkgi3xaJjGRAJIsIhQJ/VP5zbKGvpz+0x5/66QqKnKp5
8+jMEz3GOp5GayyIBNs3GdXVevJWPp+P1umZNwB2w4DbghkrsZgDkzP3/HEKy/gAySxeXVEQFQo6
JSmzU5XLgVhm4sNnaRVaBv0FXp21VuiMK6SDcBEcdOdRJzQdg87INBTEMV4UjMabIW0tcj6e1bUi
eiNACPIV/RIiLlP4WBCx77sLtRhCz1V9jLUppCwA3Xfb04XHBh8G1BUyrB+tf+Nt6rgwwXjwaHTU
8H1jPcXIcI3tFYyP/yuy5XfnW9SbVS7ExjnbjJ+rk/Q6i2tD2nbPR+LFlVcg5cNdREhdaHhxqn/2
5FBa6xoI06rpdDjYHZCxcwUQ0Az+qWdstlGfn+e+7VbSmaAMrQbam5//jFduxK1GwClZ8ze57DAP
KJo5u6tnpxz5Pb5o2Fv0+nr47/ouYm18T+4kwXT1jyXGz279WnTifnTle7WSlL4lfbJLJ5G82Kja
W2uwi6c4X9qj2qiZsO5VkZ2y9jiYKVkmfYWnXJiEwk28inc7lKOOfPJ8/OFy8TfbWVha4qWgPvbV
6DCRgZwP2bYeoq61TyG7gdj+CmjtTEHoT+f13w1tb9D/PyePHNNtm//8aDL7Q/t6WOAnbbVcfieX
FnhrBIRoW8rjSaeuR4jsQe9ZGb2c4ZCqMT87uc7eQnI4Rm9VRxBWesqXzdktmLLw+ZtLG7/2nFq5
dPKCjbxi+KLKl1xt8XO2ee5pjLqYYr7I9xbBWyZJ7VYqRSOJ+cayhvbj77FkkTZ8ewjKcsN86vnZ
g1ODA1lpn4PG0xGJyi7t5izA9ROlgnfW9tOcZ4xTmuAJBdb86Rh4n//YcVTwwZ/G2ymVy6rOZcVi
prAVDfhk5FLrHgpG7EvncYhgj4ztW1GzKbQTdieG4XMF4DXi7bNZUs8XnHGS/9jq3EYHZksdV1lt
ht3VyjdMHy7/48r/quVDQ1w3fkashh/M7a3559r4t9Ix4/SVIjyK0znIy+s6uZCRkR16+t1/uaBn
ZH8JH6/Eq7Bv71cjyVWk2aLtQnoS0hMgC1tPz0opvQp79cMY+M2YIHuHj1Gh3cCYYIDlY/jUkbu2
gAqIpKJL8Xtgn68QJGEt0ceHD8n3uogB3O0NBTz0UPnmutYhrLBR7fduD2YLsouCBWmuUMjd6b3h
cd/W+v3l9j9zgGqWQAfXivpfhfujbdWuCc/ezDYbLGzq/iqlbccVFZdKAdAOXgX1c6IiDjWJM4+3
mMRfP1QNLFGfHQUVxl9Mjj0OZknHVgOHolhXPqvwaUt7YKgFIDNbsBiaGMAr5wZGMJcTJ5tp1Lmq
U+AGXt60I3HsHj/v02pzkQkkNYJlCxgPeSgu2EodIkxEniMpfTuEcYWE1RRy5Lpsa+qlEv3uKCS0
XQCbL0WKNJEG+Kvu/6/EDISDcu3ERWo7So0x5YbEpKhFHMyky5FYFmUMDUyS3aSXCo7UfGL/0W3W
Bs1hxeINsNDtsTJmqzEYDTypPYG8RLaTLfcyf91cVjR56WbUOW194IRaC08ELnkZtX55IngJIJQE
9hcoJi9ZKt7JEnAL8WUQMHCqCHjHF4dFuJWLi/jWiUCzHb8NU7JfiHP6Dt5EzFTSjE4g1dsPWnWE
EoxZFufwQrYb4di0q7GVrKgoYFSNtC+R7Y9DnRBR3zBTTZXXUqZs0lf5UigXALbYSiByfakY4hOp
0kkUXu3bT++qXuZhq8J4IXT5dZ25Ib8LxE/KzZ7AfFcOg8nbHX6rhTdEpb8Q4qRlchJIMkqS9tDk
E44UO2C3qmcxCCQX3TNDLNusYhzfK4mDldnygva0dCERVup7AG3ew5eED+RbwcQz5CQLAmAP9NxH
duZsUYoBfnrS3UT07KhvWULBjTWnfvTom1dmehejuiQmynagc0cz/4XSA1gCNB3vA7Zy0nwsUzuK
3wx9bxujXp/km720ftHLwZe6ZpSxfKT8Pt1UQheCdP1LaVBNZEBZ9KEIeGjlq9KT8lq2GmXgN52i
OAVS++D9A9IJWwejEQRPXS3y65NXRLL1b2NsJhuTS0DRgqRE1oFnCej8IoO9BwHe2j48KUbqj8Hk
MGx1XSw4Dy+KvhnLe4+gzYnSNqP6QNQZKproMAXzASumSixn+kX31pI4w1k8EkvGZ0DaJ6ZLSg0p
o1BaeVWMWu8reZ5D0Yt8t2mK/kEk1WrKHoERMdgr1HC1TlTbTOIWLIifGF98zmudedmAK2Um1Ls3
aoH744Te7lE8CxG3RyBcFoZOpZPlpyTPkvgYEfxA9iK7WTEhME66h2pf3LW9iBdAv8NmZJoLxThy
vSd6wIThL0ccoxiS8fkugXHXB9tDeSdFU8syptuQ8FnsNni5tKvP+nRaqDVBlM9G8NcL7zhvX8D2
mz03oT7kT7q3pM6Echih8LzXQ07XT9rKU6h6LKMd4ngCRb5I9JLNw9NuFg+CMGxMC597alLgXl2O
CnTC4AwtFRHIIasM2SFx4PhkerD2hNJL2XSZlRJ2rLLJ7biiz/9m1w+yotn5gK1jyHMbpgh2xuk2
cUUNNkDdbejFUzn4HJ5LI51gTyiECKiqIUcwhEU7vx7dn5MrTX/0gYtgSU5gL1GkPDnHhxmWD5WQ
48cGKrgGZh9fvLhKOVAu3jxRE/eFZOc8TwW0/WQd26G/lw9HOvu5DEnpnl5+br295ao1ATqXX4C9
sWw58O/n8DJp2h5+TtDVtxjY8Jx5xQQrFpR8CXM+eXtFkutEbgdya6sszLSlBj08HyXYp1dAV88q
BruST8P7XbIMnQr5P8JJM+QzdaS/EWpR7wtcZUpsGiGT19Sy76C0W+0H/DDAsPKpY6zXaGcAGr8H
EW20qZ+eIf+bVULSpx5jc7yHKfHF1fi720djMrla0XBVn8PEes3F1S2V53GneXNZQGCoSA2oZPMi
7vqVNOeGIzBGVxeCevMAgQshm7eioQHzC0VaM77ltnWHuQ0AuvqAakpGpu6o5fIBHTTEpiRU3QJc
ud/qCuDoW7WKs5ZCR/Rcv/LA2JsRiBqdqm2ks2X93Z254sIyK4pfAwKZCLAQuYmsRIFn2Ezfk1fb
jdX2xz7KAdhfa7lR/zBxL+h1K/cscT26uGupIS9YebN/qZbHkcI5LewVVlQrKcTtTRdAB+XtRrKn
5efZ8LX68Cc5hTnxpY0+pUA2IlQjgNWgYglt3f3tlpy0U2GsaioIsTFJ13tinl8Ex6ZkV575Zykl
73VsTbfV4f7MNnCPyWxlOa1qKHOUdpGzDfg+GN/THgZgdLDoO86daVy7gtGI4f2HcK7E3b+40qxf
Sg3Keez2/RbjrYAlNzwhBloV/3HZMwujavT7agtMV5tITGxbiIHyghSh8tUQTeM4YT+pDxa5XOkk
D6/AlyPkbqiClgeCqruvIsodqnRRt10uIB/PNAzvlPal4yKVlFzzSxeel8+jGv+2MNqkj4SqhXiz
HuyRL9c+3gvSv2Qzobhr1M1zs9TKxFCuBwjma4EGDX4OIbP4LQRNRKqrRaI2+JPcka7eKMy9Il/J
3UU2+vROheLLSp/JmWj3tri2zFkZHtGfHUFbbTvfqcM3ZYiqmBcds6eFav9bTA564s+PVC+GTq1o
XF3h7hg348J6FZ1JAJ76gIymppGZpP5VrO3I6iLaEBVxKJgD0ujmNh+JK4X9f899oQFWKf7+Dn2f
fGicxX24nDoYhYOo5McVH652Fu6HcBHP5O5OgdQKnAfWM2wUXgDgrGxaZhyHM1wSg4SC9U1zOEXt
zDd2rJ7qXYtTj50BWBdB4PvpwWZzRLNZ69/aWHcrAJlCdlmerkrFRQ3HWWAA9zkgo5yTJVgebX8d
XMhnJMBdRGMJrCLEhifXSSPkOHLthfsDhF/FCkaW1/JFkzs7FkF7Rxi4WsXPznVKyuxZt4pUMCLh
tgvORa0iVw1lzGxADmDWjuZfa5ul6q/k35CHCqfu6K7lGmiD7+Rpl7FZwzM60PXmtjMv7QLKuQbl
qgQS/on9REol84bOXMEPwb9o800f6i+93jWgHqX6ytXUzlKv/hxpv4WFTMBCdg4+jxgDx4T0cgnA
VyEu/dUL/8xgH4bhqYOgLRUBGnfqr54ctgvukpRgHbkyH/F4M2huzrZ8X71IiXp8oUM6Blabm2+D
9ci4zJ0W6TDWX6QDeFBfCn3fA0l/J+3ZiOJLDEb2wBklZ223vI1bGKcF1ehl8CTL0LCsGllyS2U7
iwCGQNcT36qfE9BuiddwZedMNnLOkWhnQ2+yR+61n/uLFE6pCsVznJZBTOZHnuFQZv7cTOZNQtBE
RlioSB85rCmuCSiiHU10iIaPhCxmdu8Eu/QAy7hpfk/jAcEVXwp+q5mtzqjWiYb39A+G3wKQ71F1
aylK1tLxn/Ya8EwDgTmECAFpPOVEXfvVbNaU9Hog2O+nbjQK7WsFafa3nOSlkXZG2np+5xBwE3aB
NV5Sr3N633FHvUz6jlBnhdlRyXht5CinZc2tDOJ4eQ3SUil+NOStyiDUPueo6W4XScQtUTAhhnBl
+rz/f7vu2Wn69cNXGv3P5GYTk9TzJIQn95MBfvwOwdDCVF7U5LSO8o5TjHbiCpxE2gUoZ7OGOrqE
hkAoYWKlp1g7QqOrN/KxiVW9/iiOuEwrUtaCkrQiZ5Rti3yY0dT2ggXsQUJApM00qmYiLJh3XevO
z+15RchG2fg8ChooenS0uKtUR925/+u+PfPMB4/KYCnBdKlIe+fztmeA9kxx+pOXgajQ55b7na24
CXid53F8Rbib1TEXpu0EvYZ1WAooFn+IHQzs2/yI+y13H1UxIEkASmSgCbQS1GrIAtUcZNhkLz8x
/pe6sxftzuPadejX4xinJubMKZ5q/C6xZIK5ASxW5qt1y0AarHDNwuFkRpa22TLbVzuldIjyGg5E
oNBLCC/Ye0RAxTHytkiUcg7XX/RtaPC4SEWx640h+r+LaWfKdgACTn63ocY32kTtnEh8DdJKbcWs
pRFm+oBAmApqY2GDQRY4VIKWrJBLShqZ5UThhBWCBEdeXr3D3hJwDQN+9JmYVGQu+71gwHdDg0xq
K/1G7Jo+o6cpc9zVvYvbyb1uFnr8b8KHz/oL9AvlKJFjpor6Sgsqmzymmz8xjtmUXoq27B55+Ue8
hnbRjghAk0cw9uiz3LJHiIyRDG72NNqU9QNoOzftpDxdOyRlyYTL1oxHeYFu6OICyLKXc1qRZHMu
j0e2PFZRA4Q0VZl3R+nwR+pF8sXV79qW+xr1KK/OpvH+n7Hwd3s/JPKJtkXmOyAcnClQ/PgGabjP
wmC93kSjcqYOzBTdEfcOygWDeUMhaRnRzkaXRAsFkbcgxzd9jC53T5tappUWdapGSgRdFWq03rg5
7cMBS9i90uVZ6UjJk6Nfa9AkDFhK1ZM0lAZ4A42owzkBEfqCpdk7g/xsrnatGvNcDXsmR4RhVPcT
AncziZoVqsaU3Rbr9i0+6wzxYyXqqhBXuNm0RhUuDhswCYtg70joozxerXRhyVWG4Yk0bOZ9SQK0
e/sEN38/LvtXtfaVooU3A+y3i5xSPZorc9ez/eoeQD3ra0czZHUzOBZis2l2o9ZNgpQqNM5b5Ftr
mCB5aSuHvVz9gq1qzT8RPJYz7GFD60jTXSVW9NuI9LXrD5CcMiIF6FG7XkAlnAM1jzSFZjBYU6Qz
cBJk9czGZF8bMqZk5E6qinnY3W8nbSt77pwM9nCU3hIfQWULBsiSGPm779PV6TEwk0ak3jTdXtog
1PKBPo5mNBqgXohXMf5PlU/gGsgqCDnAJICl52yJ+/bCCjOCV0k0PGilHH0mb/Om5w1tlHqCys3E
uLmIaLFvLZdqbTk9Ds0/pReSY2HWJkjUjxOv6fiKQ4iUrWMmk46iFn1iHmn8//cRc8CSVFsK6gHW
iJnrt5aB190SfuR0ZpuHFBosei4S5Yla43NOL7s+HwLErWSmWTodC73tC8OCPuiP8Oa6hQjMixMx
gW+seI6D6p1AeHsHutOn0LrYH0sh/FWYmiiV6nisA27P1052BbsWBIWGR6J1anOfiwRa7DVDiG8+
kOb8voaOZEQJxLzHStvD6kOvtzAT3USC/mmq9fwQEoM1XOB+bHQJFxYcbSKB2tfQjoiMJ7iu5opF
i8mzoyB/mTWDgtQz69sziTmcPdoPA3ZGKPxmP0aitOKb1y/1Nrz1tI0laz+ctSnorIbtTtoOJlKS
HihGoX0RPXe6dWf/5iSIjtocHUQeWEGiTtmEKVthfFQXj7HCBTU9PBcM7DWDUAER1HD/kBxnSxHF
tbXO0fHjCksl/pjMtKMM5qfbgHzLFPmDJ0WPnQEBExNe4xrU0gdZsxx89t2CMpvKyV9JV3YkDDIm
BLiG52e1eCnMijmfDbo2H19DLbz4+Y4XnMUNaGQhG2MOvR/9tiY2SjPgl3h1a0PD5vXSriFLseEp
7HTl8WPWkV3TW2bzqC9eQGei8HKOccyL9FHbBk9V+vhd4YLzfufQEJmSBtVNXA14zE41n2LZgJHa
XkhVoaVD2eA5oCYbGMIeu3/Q7z+sRJvv/TPAJQS8Bvgd7pUTmEqEsOeMMkYjeLz7zFFXInD0WTbO
i7feJRYDfTmZchMpWtz+QTMvjtDcUy+C3fxtDXmly9uLWGYfG0lRJdLk4jpZTNSNjxurDP7i4DpF
bAN6J/pGIKNl3ab2qQCgKkzRMlVPPaQK3+qe2dcB1NTLADZ4LJ/fiohM0hdg/YYI8mzs4o8E/Phy
5H4ufakDUyuDZFFmr8oQHwp/zJz657/7/bsO9F47zgjBKRqGNGXwfHrPuQYVnoXlZqtDgnwhbTgo
DayEIytHLfawe9tqOf6deyAvpgftbm1QMgna6kGZRej1NiC4CROxZTXBG/XrD4ItOjyktkWBTfGF
kMkSdlGknslofszVzAUrmQ91KkzhyeEMR3gSaJy9z96WYIKD7mn05KVeyY1z3bbH1WBwbLCRfZXm
UVfjOG+XjK6mjNCKsJM150QZFZnNCoN5pf0tPuEx/xBdHcGd63ilWDY7fLt0xm8ObR6pjxhDLpdp
R6HwRGRN0H5U1dQStaBhLfDAdZ30ezxh0/uJb1m/sDSGe88mSDPIsI5MpiCASTgCc5gC0R66ypjM
WC/Mj8PZXN8a5GBftPGFNu0HI2segvnw0D9WcDblwmhqL0JIrqY7ZBXb2BjNSrhrQ8Tvh0OCuzg/
G9UXjkIm35Z1LOnJzbicWayxKlRf1JBLDAyQXi7PBSMr2PF7aueYdIMPt9USThNi3ljPcM5YQJvP
pjBn3jhSBINyrZmK6HqSIgg+YWqY/WxdoPY49WaALiJRxjTfOGCRvk8J8gdbOqR0FX9WMiera0vR
pQYEb/R3RjJpxP8H3sJQanKgkAGLiXfyc/yE+n5m8bXpNhrBhvkWnXrId+qzkh/LfeIP+jJjN7Y+
6ln2Z6XmceGPBqYkvBP9c4vwyKM10y7SU5IBZqQgFE1aUlhWQpZzuH5VH+Fi7h1Qq63Vjuan3C3T
wc+D7catYP92aLh2yq8ndIuSg6F8rSo8wdzOFXKE7izjcUKTkr9qVkPdnzVod40aX1p10UUolx2B
/fp/w8xLC3NZdHdUiL7yieHOvAnkxPHSTZdR645w0ehSfZ82BooqkiWVfgYlY45ScfgDISgkYWo7
uj1HQG5uAZOd6cubmvIO1JRaNNP412SJOGZgx6UGZUc+RQMMISPYAc5khhpRP/Bf5Bn9ZqrePh4f
e3En0+PWlakUR6lbnLrlVgiBNAeZbfoFBNfNJcpRNOFOwvoTDxvjzoB3S3Y6F2TkEflkffzBvcdY
OreEIpIkxOaDnOIKOZ9ZjdnaGsZuVC6j17MYOv91Axl8OVIJ9PJItTCmpZ1gOd7K/qo3aUqRaRwb
kPpqGP+rp0C679CArgXwJy5C5V20oakPv/oSow0ofj/189djWNupf3r5Whw3YnS1TvGYIiY5+7rZ
/aD3EFoCz7XiB9U/HfqB0UOjVVQXVSNlGNM6VfibLxefxRyl2IuZnOFf5ytAAuaAPJ8nbxuNSscE
7ddVMjlVXg9jgbjXyjkdCKFV+GmMgVy3ilXF+yOVIw/ZNksFBaM6jdF5SPE0rjxO4kpxX5HEve2e
Ej5RKD8zIPN4IvaVfXB7bmPlP9thwQWGiULeA+wrhtDzez4A43kt3w1bGf3UEQXikSw+9M2u/bYW
l5TV2V4D4Nb8AwkSoq1/yj8zbrIc05nZ5iYkbveMxmT2SqTXmFbkPUOIsE/IVF2Ju6AHqt+AsVw7
QgfpLb4uMmJa2rYCKnvggV189VZmXCyhGzh5wMEjyDEdcoNfsTucOeaXem/MveRBVleAAzfvSFDE
xdshKY7CtFJEExxUteeMJboXb3UH+o4bMfQV8+OGd/1v1p+cgc3eEwHGBgCec+iC32HyaNExS25m
Ig68THvvOJCoJPaocT3gEdpw0Y0bCKIYcJND7iiOKGMtAklh4V/2B4nX4bozujN5Rcq9vUGRfLcV
8wZP0ISeZF1nzFaZ6jHMOI4XOCnI6TaTAXTSyHhxCjMdtEwtbQoFsVO3vHhb7X1A9z2aqyAVDhlu
rlDJlcqDAL2PYJsw9Ss6kCrpRZ3iAKJXPZxdHagdqfjr9rydNSdqybh8UCMDkn6Feh3lG7DPjuvK
7V/LxhfwQoP+gVBuvcpK1RWMVGwcpbsb7uvXe+UzhNLgl4WR8wy06GFKebXbK8ovqSCDIs8TJNyC
htj9v1X+HV5jEaJ6CBU2VpsOtl2D+RXPeux3+TKsf0q5HONdENSYO0mOJeQXSFsctJ5L67eUeb9g
mjpnhuZYAGgvH6BNTVMP+Q7Zu+Us8lzI1uerpFhHmTo8KeYd8KWFfrOnMYJIpIdXY7hUQeqF9I9f
v2eqScQqEPsCnhs49Cx8t92k+R93gJet826C3+owkRwfV9WNCjnT5wdOmPJbTSrUtRMz0DVS9Xoz
lfjoE4jLoAfvCBMVSttVBp9kHHOz9hNGerk9o0cnqLWh1U13UHaOKB4xSrdm/9ejJDxh0qUlX+zL
xtkiavxDv2jhbg5aDh4SMP4fH6pB3Hej/e3SFJMR6ecEU0l8VSZ1SPhSVAtDyfbCovMn/5UExuZ/
d11fC9iQINzHoL9x9jjbGPVjlBQOxknvZKGyLJLk7zIMwUJGBQTK0oSprE+o4bnP4tJVoWKlaiou
aiBaTKwpzq7RD494hoZD84Kww+F84WFPSxrLrYphxgXoEP8YIvY+yhMSqaQhiy64yK+EQ+m3DnH6
H1oneghGAnsK2M9ML/00K0DJyo+bi524i4JBTiq6dg3JkvoRHFAYboOkIAA8YvVO7SJteZbgUCXu
YSIKw1ZomHxxonHvkFIhfN310BOPASnxPJWccF/2B5Jo3iQW+HIOkm+XU4+Pwg+MDu/3nE6fkvq7
F2fFWUehGHSbKzpc7Zm7gBSi9ORg3ynysZfr8NecKyBlUBASzqNfid+cdg+3Bh1nStI7aqJ5Jyck
1YyCkpiqhiSfAjClt+8mguYRyccX1w8AY/CtXDt+HkAO+688d2P6sksEUuS32hJewcfQzhyaP9fS
tdtqFKeBATdvIKa+P+m1kjAD2GpI4vFUnXS1OYDHEyVHFInsElOvPMBZW7Frw4SssdAVhaFLg3OZ
/F6Dp3tF9i2iu7/8x2l2XCdyhLN29eH8kuY/SDVWGOsiU3oNG89+yVSeSGQUvjtFwrlT7ew3HVq9
bcm0b04DOui7HQvIdz/odF7xtSY5Ye5l7A6UYJO2N0kV48VDPaduP2VjM7VYsWkDSnHiPMPXJkFG
p2VGqCwww7OFPY9RxVrC16J4j1kqHnzBcD348XdjQv9fs6QL1LpeVBvwb45T2X7qYDfVjVB1Q+0P
5hLzrr7aTCEZS8LUNLwahxWXEyA3nd0IhVfU//OevnkijzOo6qjbi6WqhVNdBxywn8BNLqJA0rTX
szJJ62Tjco2bO36CeguHNlXMa99N/SO2irsZO93iMSAk0ZwUDHIRyPMPkloisukPkNnJUCPVUN3S
b91WkSemM/To37HIVQU2+g5gQMP8hMjJTTfpwYFL6mprATFRIP72Ae43U98aLm74EX+GTrMJGfu5
pHJ2Z/DAoTKwf4J5BQl93ZiJptd4DtO9iTocTbb1xpfvmWvrnW8pGZW9xfko8iBN2mxDNgqk03jd
I42D+8E5dW5WMyhMKH+G2mm8i/VhISaXZdMO5ucdAZjhLbf3Hva9hIfoiOxj4iS4luU6v9ztSbkd
YJj9bkrwpFAWVUoWYJxEI5WOUFmAzlqlYh3vgaD/vcgjUGaIaechNU8x5EwDDgYE7whC+RG/oz5e
Ut+1y3jS+I1rjeFKRUKh75XQW8UUcgv4gmzITH/l8r/EeKbbp+8OS3HLcEGkC7GSeXrXsJxfy8Cr
ARs1Xo4kChqYqgjiQ+R3DNXtpORf5sXHXUgblefuExkRYGTUs3UG6bc1p/NcxtDZrvjG/kcpf0rS
yESVy0bT60oqMw2keH+c7zqbCE/xKNEEyanbeES8xcOhixO2HXtB4SdrTKptjwlolGTisMD/0vN/
m7fnxtJXABeYF9s9BCdDxEFnooLiiKaErPb4uQOS8ThixmaRab9gIlR2NVj3AZEkch5Jnceq5VnV
Rff8ZZZqhGkcTdXxbpamIJuAkh/FnyCwMn/GVbndOt0tTyH3365z2g93fB9f13TxHCND51xrYhdc
uzUD9tYpO974/oEFBndHCkeUJQIO1oW0zEeWLx3YsX//VgyTWTo+fnCOYnxd87BXDCSHMGXcUv56
VhT2YhyU3OM0ngfPUSpO2XJCwbmt8NQq1Mp+Dh34LlwpP0g5QyAPq4qALVu4Heo52QjcKKWttOdT
HCBLfddVq0hZPQSd7UnZycgh6S/7pGSPmc0HOFLPaCTlA67VnM/jn8QB+xlNHkgbiqm2fBLpH4tD
gL10r/uUUPDIbfNddkQNGbnmI24pE5AkwDaBTGsltB38rb/8m2QBfc4rzjE5XTgge+eyJHZY2U7F
+ztZiAdLjQKObUSN9C+iEMELCxWqR0bT0WJL6w7Fg3aqBVjcpmbHgP2iLwOL6qw9MDpbTR81+DRo
XOlMpZslBBxGFBVStvNxvcFCtWtbAuz8Py5kqJKDebxaRmpoRGtNFfTkLBoCX8wE4rMA9JMCGLET
CUM6EuMz02oP/hs2q8P3XpvfchS3Hb4mywjKfYpfKE9hvqqTb/WJAvIECBXdNoCIfDeT3xBt+2Nd
yLMmhjutl8EkFPo6LSnm4W2T2kHfpMfmRmhyx4fMxEOdXbU6u9F8hnIG5UPDi/FaHiHUFA7RnYWJ
wDUaj/3GFM8vsn+wEWpcePixJvd0gwIM24KfKYg0Bl/r5LTXiseFaOppLMZV2NuVc7vlrRHBmyXo
gStBfhuFNH3iZoDaC1iuS4bXr9PHjmT4MM8zNV8PzXtkAEEeYGBXDbomSuT+0yvB04iqrFfwdPmB
JjXmrjQmiVPFrHn6EX3lYoHPa12/0W75d9BZ8S6rptTKR4Er/EtYBYerBZVM0OS3sT/ZgJ4TWZmq
uJVHberjf8HYJV8iFVwcMDZlJBAyDjNWoUYgQ/mhrnMgy0y1fHcdO8jD6kFHPWHgWNQaZLcTIaL5
QieJXHJM3uv9iNgwzejv4XZoaBYQA1+ZNjNKapIa4aRbrGb2iJ2ugcALaGvGKMgXKdqTzp2jwBSI
lsYz9ImmLFivqNT0hdHrPPn5jKu/2ILrLRk2oWfKkrqcPpBvg9pW8XRKzjTdARH5WnKXVz4vJSi7
jDemCyPP3fEMKwMjSzACzfINVLuEiXv+v5R4XgdyohmvzvkfgbcLHvhkm2S0GSirLMBPPlLXkf01
iLRNfg4i2u0N4hEO1E12w2aNLHuMGqP1990LK2v1irnNoO5S1uaoavM2skGdHJtKECQpLepz1NFt
DV0YtA02tEjhxxI37zxT3PVs2CWZbQO57mBbYmEiwzlLU//lJUbCO1YuUEcmTsxVFWmDPHjMYTOl
Qk3BswfBhM8cbslBLP7bf59xdHlF3IhopckuPZYsMw1z0G+ZN4t97EgB6dKV3Vndot6EXerSFCS2
EaAIexKkBxxu3qeIBWiFTk1u9h5q5IWBiB/typnqXwJ9/77YJx1uH+cbeSS+hnnrxD7Hd0m/wIIr
iIZ2BRnYmyRfUejE3aNNpZwTKHu+dLDlbUfFuGF0dw2s6p/6SBb7iCkPHL2bE8BhmFP3RgencBjA
UYHtFI3+ULQ7Sk/m0lq5q2rMFo0LmgekkjV/LwsAPbrUcLlXCuDWQSP2cQhgvyeyaI93Eo3UeAhg
xlxTxZsWhcu+ttese4Jp0JZjtyAb0x2RMSH2K0MMF75lTpBjHiiemCh4LoHpFjqfncUbDo02jKlz
C6B+4TzgvnVquY+AUfNMkT3Y77FN4rdmhrvnYq8kkvorbwCmA7G85qmIQ2WPAYVnVdSzdbzT3Kk3
0IS9YXHSxTDwUIIg70E+mQPtX57GUEWshUwYoEeWQ4BMzV8FwOJuuO2YA/k/Ia7QXAKWGaodxEZB
UPxOjleP/X9bQe2sZdE0YzZm8te6e5BRivV24bQ6fFpXiqUko4RwteOcFcwOtue2NTE6HZfR2atq
JkHBF2+jXIk8K+hYuor8PNOP2EC7dHHAhkf6fzD9voBKdpQLNUpWPONJwGvAQRUEXBBIlWAeHnLd
I2hOf23xCkXd7wOrpBrqo68SyvA1+pVFOg3zLYSHqkhElYT/44fqTfJ2VSSH0M/5LtNHTvqfyDcu
0Fa//Esg5XSpvgjVRrKAKRoTk7MmkMqEYOGABGc9AFjNcpPQsXzMukvxj6fFf9S+lkl5kNZPZWvV
gze7NCbgz3iNClXn4g9dfA2qxPTYICrBoyjSkV3HJdQz5lwGHko1XrcR0KBdorFVQzRsuoxntUhz
/Kq5ObWTgQ5qK5hgWAOg4PhGpu0TEzddia9+w1HqkFq6Gyyd36tIiWlzEOcsjGLH17Yf2isIH9fy
R+kYKiN/mk8dQUqiBpaAEK+V3zizQznRRjKSssDqMXI/BDk8ZZ8GB5ifCrOoSQ0q85rpCCXbDby1
6pSUMo/eV3U7BPcM86UwZk50ZAQvMEfcplRw4qws9e9pJAmujPVNNwBIPxeA+BMXuP+EwVMM5GVk
hQxFflF8rKZDCCz/kAyYFHQb3s3CoUElxaRGEJGZM2VFIGbD3rh1mt4S0AcWe4TpYOEm+QYy+X2w
yYBEedHvV+c82vqAkqyhakw42DV3AuKeuVvrXl9RR4CUJ32r9BgNxABw1i1Oefu6HsEESxS17YwP
6Q94i5guk4fqee1diPrJQUywWp1wOTv1IgcOUEaC+uEDPJz2r0ijy9ZDZfTHrOAmYc2us+cPEKH5
8tgkEv9RcmAD54K9+OqyNRm67SkxYQLjnfaKQ+R+vDoZkgaPpUiAB9W69B4LM8w5mYl42EjN2iNV
bqtNhkabhal1JTspgxnzrXvmiPLAuXEVkcmWGW+kjjRfCdYdOkzowfkji3vgpuCYfNlAUE5wYoCC
uooBi+657ZMv9NT1UYRMaRVHMQK4OCDTnQKlAyHuBiKNRBn4mUFgGJZ+X+CfnqzpKznLmnmSEwbD
E4cWqFodOXEE+Z1j8mkVVaY+K10tuSE5CDTUEGcLn1v7kbDGdX8GuURZsX+4/hocPnNxyqkTH+1Q
J3sZ3jdUBzeqUc0l/o8wjCSLNxjK1Ht7fyb5mM6rhpRNJXaKRqVcFkwVItH5lbjmCWJERSC4pwwl
XecUfP/4W1tCUoHm8Mvs2nrAcuqse9sQ8Zuh1sb1xgd1M1RqwpTEkD5enoBBv03JmSX+4BswVNQG
rUfG8slVwBGYvDXxkYZsGyt+ENhDvRpVlQcjyJZxmn7zguc54bkHpgU5WvYEGgRL0M85IwOrvzhS
/s36Lb0z1P2SEOdKWJFnPutuo42xZmOukNFNFewPNu2xcLjg9DDQDryLXsg0TmhnLShUB7Da3aB8
tNGqfrBLbQlPVclAPKh6dauA4xQ5BTctQH1ywi+6OCs7vyeEAor0qNsrtYvtbi5SRGOIG1OqL0eC
ngXP+0Z+FtAW8RJ3bj58fapk/etwY6nPF7D/3lX71egRPYJa2cq4eTlm6gC7wrMp5FvmIU0Xv+ce
BtKwsB5thMm4BB6OVIhS+72amkue4xaxyDqvrd1i5qvDtv5GM0Ot5/Cv75yNXwYp7e2xF8Jl4BmO
lzCbFaEPM19nZk7CaT7GxeqZCWjwjSErN54lIo7TR8+oc4oyLjG6dxojjCtJoglvyygoyYJ09CeX
BeKmA9asH3hECP7XEPeSEMRmn7RZt4l7PqtU/UT1jdiTLod7STOarfNRf4vKuu8zWSSxBEB0u7F0
17VsMmKSVn9Dn1aRJ2ZQjfOsdLcUcpRvLv8RaB5QAVhEh/E7BSfKvFDK25pTLd4mdJcd0awLT2cV
Nz77OwAkcdH5bjgKPJKXTF4kuxsrzE6HNxlVdobwccxYdJ4reXEEANtY5ig2PasMfabdND2CZuhU
321swoLwT+ZvZGj/KuMC4vIw5j3FWyADeoEOfdB6xPz2I5O2lpnfi4J3IEThJMU8RV2s8ABH5dP6
7H5uCL0ny5JPLb2973kAsHLJxWasiw4fDBOqS7yQa6p/eiH2+vbVPTvAg6MPsTX3VXEHHbhJoXHf
rsCak01YJtxhKjaqT/1wyFZgsoOE3an9qZwBfqo8NgsG2DPyGvg4nx31MocXlHyyA/yVB9BIK19R
FES8xqCnd0BcDIBplfptcxVAzuFHzylPKwbtow/t9l5Bftw8H/M7atUV4VokmeoFpKaW42eiKGf1
xDxlIVklXjFBIjB+mONHEbVdNcdJrIwsH0XT9zVU4Ip12/tb2BB5/d3wVPtqr6niaceSkyplq1Kp
N/Ob/S/mJ/bN5pKrtwSPWjlaXvUT/4yXZP790xGAMCB1YJRGunGYKemaBudY6PzBSXF07nkOMHoT
saZVR8cuFfjPdnNI85646v1X8PTejurEkuvpC7CSTs7K/ShRRA2Ia23YLI+iDLz4ODxzWEaoURuj
EwNog88uWY+sIKi2kqEeFfP1UJhJ2CtBzrX/IUY2GJRUH7DdJs7vzd0TCDiJ8VABXJChcYi79ADC
2eX1Jw0Z3hijWTPHgnGJx8Po8UFa0T9jfDMOQcHUMrVI4242lEZz2r6L2EXOf0JexeyWtfFf8dMf
6+/8WZBGmua8Sp2WjqniBAYVqKmLoUyVkPZz4RTw5hM1D4UqJE1ZAWpdV8whti9X7Jmjs5TnnfbW
2VeAB7pyMvWoFZobJz2e4ORTfz/plty4PSQwrhv0YSrQstrc1sReVLqdhaVKTRcKAx8w5MLTD3/W
9BoIbjko6v1akUsLE/ipfX56XlMi4Ps6wGqUaQlqyKi6vkC6WCzfU4xKkKG8DdhfjRd/aMf7OqCz
mL+n43cRi5AyDTjPO+Hk0/iqZUSMTft4Nfvq5hFwDYh8N+pwGeQvsm+lJfNwQMLQIr5Hb/4joFQa
emb3pJHMo/KlGE5dniQAtj0wRyf6vxizi2UyNaWrgQn+j/cM8AiI/nyxAWMPIjF/RB9PgNtD4jx/
rz8RT4Il44XKilDHOtuI5nR939ocfmSuiRHve0orJGFH2UBvtQkIBOaBdjuxTIEICPt53sXllwfS
MBao2btSYbFzGh6ZZt9OiEcyldkD2C912wlq/zi9Kf8VPYNDBVRUbj1aUdnFLqDHqAvwBT3c+uqu
KdMX3JxsbuDOFdxp4p8nI2wtnWXtiXN66XQzdGBM1Wq7wfX3GN4aYk5UWfFt6YKA8jYnC77ifkzk
ldnscxHJiNILNSNaLQK9+3FEUYiXMBFnJYEbZrsuJSW6Co7fpYLHRhSt8YQnaA38Xrw2+CAz8u5a
NGIlWy/13eKy22ao4DLk0UqG+5O8c8lJLnnn0Vbdqdvr7qaGCMwYC41W7LLLyq+Bll8GVB6nutX9
oiDzHg66TJsh/c5mxnU42jLPqyzGrf0rM4MMlqYaI5zgyB5NTlSXyoPY6xt0MtKHuy0j4lkNBZIq
WRvzNhNRbWtwVe/8yD89xdC7+UBKAnZY8jctgUMRYpt1bzgelhP/3V230fxAAvfRxErH7pCvkMN4
qmNcEuPLSpnZVwl/lZtj8t2CVszalG0lznCUih4pRXeVHso9csckpRz9A3CRyOmNHQ9Pnk6yUyUP
hcU2aAf9FXDvOXPsIrsF4kVa+7yHDndoLFnCE30wA3y+J/OFnldwF/LcS/FTApZF7PMXq77eMj1c
DjzbRYIsM7kRK8tre5waNl/SeyylnCV6SnmXAbWlGoSKcMpl2Xh31RG94ksbxdaBj6EOmQ4R/DFV
JzvVEB0nfrx1/0C8c5O4mUynvVyuok8Q71LwjANPmuswp8oD47PHIu/ZCJ/yofEu6mMwWnXWz8Nk
lQlGq7fADheHDghM1LYgY92Oo6GWIIHL/yaCX9YGEvrNNe4gqx8e5xikTB4dxJvHFgB33ckcCTAZ
pS7NHyvanj2Fb2pUdlzf8c9fCMw9Uw0YJLpr0TBSARRNF9+dFgg+PXFacm77xbk8GeQ2s2p/VN2J
Tr8GF466yyzJJMWSuWexsIJCM/4qvAAv7muKWqNkQSahpO+NdW1Q1Su5mV+ZjWU/6rU+zEOBTbwF
Pj9cJ3aT4ap7V6kuMDDWgaUzJf7WAVQR3PoNRAPUFmAJhgsaOO7uopak6m42b46s+jRMeR/v1N48
uDbI07oP/HKS4oVdPt5DCj0dbcxX1mh13qPrV4jVHNKYdpHbAZaA1390PH/NRe5rMmY5Cb1x6h0v
1snNUMeedI/2Ulw0O/NB3mvwVqmsxbRrbza2EDpwhDJTfCXRiOSa/zsCAvjm+OXfSYMPNXjFKR7M
ODtLVyMuSLcHB+ISfsILCBLuVRaIyiILFjkhEQn1eiLR23c49fSI3PID+daRPOApReYRmxtK68c/
Zka5c01t6EzP7bfidcrpvcS2EQKcJ7bt80LfogO+0tWsrbndQAeffCNs49gCyZzzfGW+JENdJrVB
xsdh6D5xo1BUZUob1SpO+0OgYA6R17pmlJRLO+mltx5kne4js5gp+iq7kRXLWxge4Dgrl0kBKAzA
oDLXd0cZgOqNztJ53+Gm2gnig3+4boyWxpZN6Gi6sURDWnyTDUbmA2DDvMuUsi6nE57a2RjtV37r
8qvV25GF+5nRM8KZaiVTKn14uLQi7xuLOv+MCZMpbIyxE8Qb5a36OheCpLl21sCf8e0HkEtlq4nN
hv3uZh4i2WuoQ+vAYjZgcXtAoORiLk8dvrg+uInIX+7rItkp8JK17wRDuXSVM5WeVYkaO1OhA8Mc
WtNK3xO2BUJbL9OaSAnV+Oam3BsV7TivbgMk0bcpRKsMNGcj4Bxkr2CvSnCLF+dzcKFukF2bHHx9
QMhQT6p4oC4PLM3oBfvECIt0ZVoJ3TETFHhkv0i68jo5Nkkrhrg5JmtUtlSHRLH/4jM0BvhwGxxn
rp/twmN5A6MNQOgqMQRJN/BuBUXM1l2WqNj+VWofjipNfRiNlUUTntfpO3nng21k0oO6XzNiO+UT
pWVRAot11Z9HBaVQzRgPPWtzqlK/MfFb38Eg+VrLt1vuOMxcHN6Mnvc8rxqkgucfBx8p0UIQF4Ji
Rs0V2HgitNg4Iam2Y69MScuruq9jvvm7c8LwfIzWVg0Kc9w1FHnbU+2if16UlHKQlsvwjrV/H86a
nXfXPpDPhn4IrdI59omhUDG5F5CSEPqv6Rn3zFON92032B1XjSMSPKLuJwb9U2GVuFM0lZPYUGvO
QwnfOniXJWsZVjU+APNaNGpDTMrk70Cyx0HWosil1AlJQbQkLyHmbDAKyqVU4qzhBZ9EgLgXU4Mj
Y/v88XVukzLjCPblKT/3LoiE9Ic4Gwj5Le5EBKM1tPrBe6ImtzAYrNaNwOCMk8h+D4MRoNtYSKR9
AlFvn2ZR3A2gNRStWFi/LkSl0cewisQUaXBVhFhZq0A+qY+IeBt/1RanIbYLmd+Rz+satowFK5/6
7Pugwvx30PXLKUEydQV+RK9xya6y+6i4p4eM88Sfrvr6w0yCksUWt1S9a8Wn7WYgFHWO89Hi8rIg
ORv4Is0tULTPDv4cxpBDF5J1+3fdKZ2mC/3xmEmYohAHMED16xRyKoIt+juxNmMNbC6PAxHEQ2R/
reY+dbenuQym2Y21dwT3hNw3TSHMGqimzGi+cKWZ/s4/60pOTamHAvOkFVNOQpIx3NgQvTUl0QY2
+2ev7AFfZieQZsptlUhcRzpps2xNgGXB41B6haYSOxMBQQcbBYMQKpjpUj6RGv10dBUH2RUvD/pO
ScPpBbBPkxoInvqs47MViiVzrXcOaIbkkUel7zfJFKip/w4W5QYu06qinQoLEda718tPfrWtTrgz
H9V+wsit/CjsdrA/F7Foyw/WE3QVtEQcvauy1rGW7Mtr+txcVrafY9qwH7nfAG8fGAquT9sealBw
6j1Ga6bp35NIegeQjmwexTRoaCcAXOjH62IYVSKVnU/3kIQUyTsxOT63lMRkNopReV39iGw2B+UA
aP4axBVk3buwymOKF+1QNDfnb+A0veWj/OyTJl6uxrVdtAWSIpC1b4KiLNsRqUF0m0E/IyfG486d
OD9I6geS5fmNTkhz4tccJVUCJr8Ojbeo7Tf6Olj/Cr57cFydf1kWP81m3KQBccyidLrhz3IC3fPU
6Q0+V5XQpwbSYHkNLQONSuXsLqybZXRDdBU6yNJAJwb6ef7p/BiD1snCYBaobfEkHYh+JoN4/oN0
gFBtXraukqFH7g9aACWMSNGYVk+7WQoM47kNnM2EYvEx3smJ2Ib+kFQ7w0sNnUsjKKmuZUPfnaiB
FeKzrO0C30rRvJQA43+PVJ34kl+gzxxt45lCuyYBCGv3eFIixW2cyOsGHXJdLZyuQBpU+MJlEBh+
nsCTnxrTa4HPZsOQX0UJxfuMsvtUbBVqoCJmnZC11GlpV29D3MQP3BpdLq6HlkkUlXPC3I/w9uDF
mARzxUJk4zykqWHj4UjSJ57P0p3y23aUpj0KsaaJeDsMPbEwAOjdkBqdz3NsYV94hVJYtq8ifTgW
t2rMq/gTrnFZ7rEGgCW0XOWnaNqB1ikiZwIM3p8RBqJB9+wsVfiHuwzbUFGBkiTU2YaVtmWcznwV
aal3pOTYbOXPuc5nFAyaY26wo23kmyhsYTcjtHDnQG4hcvs+VYB26S6O6JgWfLUWilKurVbXGLzi
vNsOhA5JZFfDD2x79tn9EQceWX5EqAvpyVuhiIyjnWz2QCqAialrNzWG5PBJ2mXt/35cgZL2thWy
kLuNaFmfKKH/M3QsRzX8QK9s3ootTGozg/pT3L6nLKAqYauUZLS6Iq0g1qJBpGnKUNIVyfQ1TizY
jXXE5Mw6m6rHWd6MTS9o8yC/HGapXz9RLxwQcBBXlut2AzYJpa2dWJhLrhO+0w1/RNxWapSO5b53
NBqs/S5NA9AGiyoMvR4DFY9XGRIOlfuXuccgdO8GKHiXX6O8J99W0UggjuNGnwMOfLj6bJ6ugG6T
bEMgSUkSg3q8lqI97Vg30V8nYujZS0KrZIMjiYTYrgtMajYf6FiIAJm1EotdSSjLHVCejKg/x7O6
xk3heCsFvuw+9y5Z4gmXQbwcsb71FzFc4KAuSQMi4iGCi0sz+pfkdEzYx61JhHU96QUVEwgbiAZH
18BdTQK97SCBJpizPx63QD+CiI+It46owHyih1evf+CLNsvUJAif1hYuI1HrYi1kc3z2IWNQVya9
38nxlcqolIcf9y0t+cFhCgdPXqE6XE9gKYEnF+tACTLmZ6CosCds3fRRUiDXT629emvWFtxfTbOD
FWm1zzz9W4Lw/jYEU5Gg4/0BhgxZmOtZU9rBgNMIOuqJwCnODJTZ8f4s6cm0QPGHhXDH7e/Lo/fk
oWuAtJs6HE88w8H/KTdy5zzmKLwp3kXJs/IZxZoelApD0B+8EbVL2HqFnYSBQi0FJ8euwQQzG4DG
/2tqpeJGOtgj2Kk9X2BO7RjKMC81m37/GWkt/glPQPSoWY2RL3Vju2SeWLJM/Pn6sGNiRcol7ELU
5yqNsjXXkXtI1335tNrxpUFVtBNUCrmATn7NzvobVWOzJ11O9JxS4sbwbq28jdeYjsddNwetWx/8
7xRvoey/FE4Z/YRIOZV7h4UVBzktHdNpBJPCEHtoLBJn0x+yUofDeWmcHtdrIdzsugRm6Z6c/iWU
IEMJ0DMrEUGG0vY5aVGucz/tXNWTPWsa//DyifFoWtW0Zyqt8a49gLeGZ5oSfetmNpsyEQ5K2WHk
oHcG0KkODX4Zw7lD4TcRA6RsBuvoJxZYuGe0+sM3JuvytPqd0MOw3Lhf/KjtvUvRhzUHXE1LVHLU
UuwNXmlwhWh4N4AAXQgsj1S+dORvCtapu6OS6Rd66yQuiwScnGyWwMtBc/QMXJ8SrV3i92zFfAJE
2+GwCFMS09E9pcVESDv/bNd5YovOORjb3+9HeZrab2nNmJPo7Ku2k+FQle3vWuudaHv5rRPudIAP
fo8wOLA2KnMhFf9yYhsvg/JhYtvRpbmTWktVt8anyTWShHthyblJfdZ65BSLP509rRPD9r1O9wlS
pKhcNOoO7FOqd3HbB24KE7Kk92kNzAvCWNMRF7+xlb8BXkXEfgf9fAjkXtDoNlP7G0SGzJoU3Mn3
b00PG5xOMEyEwRN0JN1KVlBqqeHtYalugC9Eu6Uw79P89guZBKnltKkkLAIAlDgWLmociYR5Tn6S
BGvCWpqMM2hS93RA+zqKvxWwWOGGsIMCpYdvQL1aPUvgxD6lWurANcaBb+SwwBNEpVKYahuWeXx1
39ISi8ASlNe2Sy6Zh0O6+DEUn6FsLCBbz/dZ95+O3b+oLrg1EoB96JFXsj+Fg8HDIrztJXTmSnS7
Dw8o2Rhohs6bcYCQVY4MVpGqN8Y1RhwUBxdXrnzaEwLicMk79SjNi///Xd1Q3FDVFz8jMrImsxpq
XYLVrgfDuiNhW7yinKM1rRFuReqVu75pXqy2gELByyiy41lPlEF64P3ZEForf5hD6e5bEHNOPGDj
4pvtb1eliGt1P695HeDbNwqAO9sZ4/kEJoyQ8KVzz+Iv+Cnyq5TZoQrseS1nqJ1+9jL0vq2q476a
3ZfLQzsLFg2FdyGpjfEAHmbkMRG85pAxUj+mx/1u4OweSmEW7kjRQvBfUhF3mz5tIeiEHpnTw8S7
Dr/gsw73ExEoR3alzFLfM7xi8gjRMR3l0Pm3H//ey4dhEHHz8UQdHD2vDvbfIv6xsSATl88cyUvv
inF0R4InmEAJeWNrktwTTW6TjwGqm7JNMw0pkb1L/gLkxOzu/+uhdElAMzs2y9jiH3EjE0j39W4N
L4XuOA4cpe+lleKEqekjejL5KiTB0PGu25253YJ2EkVwVEyccxcSJL91FmD+A5PBY5An2kt4HiyK
TbiFpaPfdl+2JoGz5cbIAxGalEAyvE8ocejk7xDmClLZXgqUoCllQHLexzD1S6TKmPMucIgJUg8x
fBTD75VV+YDDwFIFyNQgwx9noh9caJ3eYfnyTnKVXy4G9UFXr7D5coyOjFn9V9f9MfwgP+8ZvNZF
/iTpF/MqzAXS6JI4WF3Boo0txRnh+1kCZBGw20KH4rahn2AfUcYewcORGSea1yj9GAvKRLd+1iz+
ECBkEIqvM6CQo8HeAAZj+trPLi5RVY5w98yfsWKsfqJOEV3djV7K0ak0CQIlMGxYB5QZ63DVAp5W
IgtE0P854dSktx70192wvHaNZsD3L8HRmg7lc8A4EOjF+wddMD4xvwkbfWC2b1wn+7gaI2wTMVEU
gItPviqQBTuf48reLdiGvSdWEDDFuMWJ8gk63VWF4JT7y586Z+tUb/LHTjOimrbey9XiUdJ2z478
qha2wkA0pL4gPwRutcBOR5BbNt+iFw7J8f0XTDYsIfSZFcjZy+agwWxY4ns77mYGV8VPcorfh5R8
U55mrH7p1zgZjjrzoNOQ0DJPN1gtP062u7Bq0bAlkgsTKTdATBStkXyfAsrX/lVRGoLZB0alS8iW
aDCcZ8+M24WYuHVL2zd7ScM/vNu0ZuJAysqbncNaqefgWQqaPXHBLIfyXuYMECEJ13GRlBD862b0
GKgsaZkqwyk99A827aFyaUO6sF1YYCqPeeXV1YNj4dw4UKmZmwRwwn4VHdvIgaKeVFndTRCmFKGk
rx8y/T1xu3u8afghQlhmRXecAJb7y8zSkXp8AU31Hy8Zhhm0mb9asf18k+nnri2oDKZ4m+lIq1AT
gwO5GWLFudK2s6rOWXxXs/C3Nf/fSIWFMpCQ4Nyjxw+YKAF/9b+Rc+SbZ8tUHtPBnGtLissoFLF7
MOzKhEQfScd3f180ZrD7UEtv1CqT2/YHY9mn5PMALAGZIq1k7/L9lRXPuPxOWiFrDi/PtyAm1SoU
9TLVAuJw6H08/Ikj/2Zdl9XxOUrehxQrfk5f8BxJJeULveLahwgAlV49g2vtNnuXKy49GgAG3veN
/QOM66lmSnFqkYM/g8R7gknpExSKZMaITqPHytGKDFc2hIwFrj70IXFVvCejZo3gtR57KIqMIIjh
RqyHG8WucUhD7Ouj8am8oxMEtVom9k1Z+JQzhzoyHrJuoDdlYR8swPl1z3A4Sdg8YD22BYgJ6XsC
sz3ef95roJz2NNlgsO0/oP0KopcWaom+2LCiTlGITjYi+1GVV/7d5Eq8OH1lNPwmZqXbalg/cbaf
M45KrcPzdHm8zGajhQEIl+RZDyozJ8jgpIMpeYgbMlBIumkXCMF54VfudRFrc/1hwY/lfM1W2Mts
hOzFscze7LzSD5HQor/SOMlcEWk6kv7kb2wpZVO1U9EClq3gmy940eIgE8JaDkEx92kEvKdymaUe
b9wWp3BqTwNnu1EJRnIJPVtbyJsFjA62acM8KODRzPA07RdRM3bPiK3Uz9PTFdMd99aml92viNXA
s/K392IUug7vbzNpNwolSUoqmfk6WayLx7egnpePxmlpQi3Jplry4LYkTIzH53og1eRwNpDTkAga
Eg9Nog5rFxybtOZT6uIwKVUQj023XJ1W/wD+mRY+WwesI1EpJAdI0s22kxhTjMkdOmiGsBOXp47s
+4t6wthxP2GaEWyM2bohip8mCVsfgnB4PVIMtPZgDp0K98vxszFTaTbUlc2gGZENdIVtGCM9eOZ8
7rHpTs9MDQB+Uf6nP7vbRcKV2rtr3b20cSW7HoLiRWZSFX66SKeSE2VggUBr6xTmBGma3C9lScay
zfT+7s6K9K9Arxsf4X9D9D6oJBfBq+YaBGjeOixHm3MUhhLHeo4pr+7pC53LQRZy6Pt9tPVyXYvQ
nGOeid6/PkgMG7CvX6PAiyVJPu8vO956WRN5U/5ys1YIPd4hJTmb2DSUy4pppWd72oYKAD4cJGew
C8NxWM6kISE6mUHdNadhODQaeIwPQ7v/nF0GK8+7LBS+tkaZjHNAuYhwoOQyOF40hR1mTVfTPQ2a
WStp3noB6k64SRDQIlula+ErurfFsSydHWJt7KVv9YX05pWSOUfg+7uWstIguZeOGmO9nPyGMGll
vmjkwRh1aXt+jfjWvxrtFQXRCx6zhXPWzU6IAmpPyr3tODCbetyB3xXl4ubCU3cX3/I+mirCTE8m
OI4/jkiNqthZiml+KOOmrRrRDxV2NqS7ut+dj9pbADT8aYUFqegHYyt4ORS+bOwJvzgTnSO7jHvl
pAqflU/HhgPaBm1qSn0SggjWYrLfc/wSX5JOD5DiUzoYiJUWTCAnsfS+/Z1nscu3YNVZrbhtuSCY
Tx2mr6+/SsRJqnYUKdmtL/7pnqQ23OQwvu2CZbHkH0K7h1xGAgu/JlG8Jg2D0I1AbXTA1WthE/2f
eJsEd+OgXMib3uhZ1nzLFxvs8BrSReVUDOS3CxbBrVgfy0JRotRx1iAscdWmSlE5pWw5NsYzGg9g
OkNzP4N1NPhDiIkS07vf5b1yGe85Cb3/pOS0GbEoRHiX8AAqYspYNkIkCYkaxCM68KZtFmw3xx1i
lLkjLQKVn/d/B8jWGDke0t70FcLPqyC1/KvWqYrYw8pUN2Pnqg9/dtg1dSjmrOE2cTLNM/C4FEPb
U0ovVUSGrwRW8iC7uvQLYZ6i8WDkN53M6C+s52OUPhICRUjJ4FTLAD0Vdci3wp0vk6DcbLjiPlzj
6xwZ3Vh5SBY/mpjSLOhazewmRaXR90CpC/izqaOYl0skthjW1Ldc49bO5MCP0ubqHBAXkvv7xlLC
Vtr+IQtY2jzva6SLRNroD1zIg/I/o8Jn/mKRY8cAU29wLfkajLnGz8MRpmmSA8CebWIihUHc65y6
9iyMrSAetS0Y/RBL+M5lNhE9vXc+KzreOJ1SdaiCJ/KYOVHnJiXqzg4zdpMd2ZHeDvLVH0KcAT6U
VH6V05LgipEYkYU4Ig+pocGmUTRbrzsLVhZXR/PIDHmfatXi0aGCtqtjcGQ73Bwr6pGdLyBZJCcw
CUnmKn4Tty/Aq420HrGDp+K2t/BR9SaSnrLTW7ULPPK3mNKY3z+pqlDjcWdMkk6J8SLO7bkQ0pAc
TVUH7RFFQ/5EEbeuL51XESDVg0gICQfaO7xcFLDl5ivFvInHzK/Eu03i3FshHUbzOf+6qCwsbvgx
5i8ipyxX5YE6w+znDCWCwXZu+3oGl8y5O8781vj76eQ5xh8F4Hb+XKgUbGcWhZAB13Dm3Z1CvZfV
7NFmAkTj2SmZG7q+JUilDhP5ZFnB6iTOPcNxssF5cME/jRm8QjQW4mqO/Rqv7OzM0UK7YBmRxE8d
s2hebkd609h5FRsDQy31iyhlYgnelmhm/+nIBSoCjJqKCiPNpQQvxesHplavS/QyJPs9HC1LBw3W
RfHO0PqKY+StvhKS+yjaqBvnBYcuHSxDpKWxP2IqB9Bfk/2lEowBf2y+7oDJ0jzswERu/uFOLZ5O
naB1YL9T7iG/AuupAcySOV9WVy96Sj4QhKS95U4RV/l6di7sZYtavCKWOpJT929SkbKyhxkN5TuH
2RZpu9rCBXG9Mjl3OT1cXUFTGvJKhG6bkBfA131d+s4oB40FSZjnOggOrICU2bnCln9GyyPNZe0v
C/j6uG/9GM9ey2qqv8cl0P9sUalGHjfPQEEObcMAzMkDWGbEti2mrOfwRBVO1/4XyPKrW0YRaV7n
Auu7itw8zE/+Wo21i1MyYrSBmb9mOb+arSp+6s8/LvooHY6IUTR6coLDZVlU2i04NEhgKgur+sAb
1xDUmjTthcpJc8QPhu/BHZ+EvoaVJVBzw7b3zxORQAEYqqx2SzTETl+ojz7KMRmtdFkQNqqBR9Jc
ThOuumLjTYePZx9qG8q+bZ0dtA9uFlkDoENIl0JerYIORsY9qmXK5dgIN3YvZ98hRT88zxDWQWPX
GQB+NUWlIzKV1CJq9tiBcU6R4cZ39M5AruIJmPZhiK15U2h+idS2UjcDtk0i3PsWbqZKhEeYuapL
hkXNTcCoYIwf6AoldPdNy9nS+zDP0fd2WGcp56+E0tAJg1lXeQjMhm6zysWWvyV2yQmuys1MdMMC
yDdn13GfEVelHO57S1NmnrSoFvCBBRc4sMoZzUNiWcPuyv+ZwKdHpojrXRI0Fjr3lZYwHo4IEjVx
08wqbSEJAdu9gvT3hEHZzDjKopC/QJQYDzVdauuUQt6cr0ZQkXWWU9B+bCyidZ5JcgQfbu/69YA+
tAvMrMssnjLUztMmlE4il+eWp9mdpVO3Feb+13TbywBEBqYz+K21C7BiCXc3M+4KiNb9h9r7IEbu
paNMUrZxK6R5+8DEJgF7Oc5UGD2D6TCso1wRjRusYOrycxe3OMXI2/h8OLgr6zPeovDD5B9chc7R
wBEexMqhE0HkN2Xwr//RZqKCqYi5VY0ft4SSfetycJu1V5pRJmwoMTkHQoOheUJxaEElfD5DwCYQ
PPjUHrkhIWd5M00s0T6PFbgTJ8sNvvuQQUVRbIG+FS9zgKEAkXdsgzasg831/mAmBm9/fwKimq2p
sJoTVpexEBKykqP8PHi/v2JJ0l1y0eERTyI647P77/aYTSHC9OJSQ2Lo6Wgekh7sHwJoc5iKjjvE
dysg9Dq62GT9qxdh/E55PIm15XxITY2y8R62vO3BEZZYK/BNtFzEilmJ2GXkcnuIzB5pUU+NImI9
/spQv7HM387gqkaE10PqTpdR04SeyxxbIDg3TWo8hbAca2LeEdsKJlik1/pV+BCatb8rrt0TmG9s
/WBEhDaRu7LNWBj9GjSz9f13cyaZMTMEbXvh+A6ei71a/4QnpPohFwUGWa7RRxG52g83JqwAL0C2
emNftBUrd7BMkcXL+hwb4q74oMbeqLncjWbLeEzbJbjlObv/w2SvgoqLaF4ypb54ajy/em+ElIXg
9gfx34lozO2YehAvTSPP0t1tGIwVyqVOqmOwdQTPTLHMfTs+/PaW8wtNXbPjVNuWztu46eWz6WSd
Loyh9nbsLKVlh/6WEyyrMGv4p4/loMyj+C7ORYQVLJeRey6XeLfYg/OMdYIxb4XC3IuGy+bPz5Er
QivvcB3Uq1SQLR+GffUAFw4ogzdbJRU/mOC41AXbEcLyQwH4Gq6wc5a99I626FDBTj+eQWzIi58Y
gZTjbYRMCUbzDrzxszRnZrnUuHcB/xtR5UkKj/f6vwA9T4GY1H9B3N84oUvUkoYUu8/mC6M0Mmfp
xtgQMmYk3Qb9DYX2J+jCGqJgq5eAKwokuGUiz7nCXvp+f56iJKX/opBmJuBqod8EeahR8KDZq7qz
uF/RmrxNE3/7vTH8IuUSAHnabn0Lr5Aik2r03yLEHc1C8SEPeG8C4Srb4VjMVkZz8nq0VjhPNioy
0ip1vXWgyOvrcPwG4o+wrxckKrdpqpD4U26QkucMaudwL6bQcPdH4un0F1AavWFmNzCB/h/togeT
hQnJyedzNsCqW8Vlls8Vd2/afjgK2QmjNFKeslH9bKv3Gz3L3I+H+ZBoLgR6ThZdUWSEMuJUnHXk
gSROHzTIklhT/NOO3EMIMXx3dCMvP3vp4CiucimTj6+BEtEeLouTqpvVJ12fDMhGZ0HshRQ01KCo
d0OMwtMqN0YRfYvhtrv5Q0yIE3i4lAptFMyq6PDulVFaoRu/QKihP9CstcFg99YJVgsKFY2/26MC
u4uukxRzFrOqu2Je8zQlv669ZqiGXmKzyaBlTwiTmhQMBEmdPRqdmuQI1JgJlflsbRilU42Yh6IV
dQOG2F13XSBe6u1p9eZs0m5vF9nz9aijG1by5bTIS9vCVd0uQhU1WQ1Yk8QExABWPu1fnEzZcmRH
C5E+KoqrsIte/C225fyVwQyTbcv+NuuxWLlVmhvVX6OdiivF7upTmsJcV2X7TauiNV0U6BHgYXco
W0DNTS28o93jrigePn3LHJZgx8y789/06PaouJ82SkCFBpMX6Tr5OeuN4u4CdNvMuTXbTmA3C574
FZxNf2/krYvxgMWVgxgcKNkoDWhzxM78gFAbqXSC6hmvVnyj7Yxjqa1BO2idnIIJGopbV5JKNui9
OKiIsAnkZRLtEiWwCToAjnNH0wDKSX6WtxVJMH48rFLqf5zn9dY8CknccJOnv+XNIQBSUKaIMmEc
3M/wwC/OuvWYwzYTaaoLwICXjjWBwGLxWMhFzP+J64eie3t0hZNaXcAOhmNwNaeNBdM1fklySAO2
FpF5epLLLkhQNHj9eWDDIpO1Pudqnwq74XDzQ3cKiaVUmkb7kWFt49jTP26z5hvszFMCqV+WIaHp
SDBt/35lMX3w07y2HkPwYPCGho4QEek/bTDSlAbUsGpgIlvCKw9nKYISHwK2pQOvWKvCWOJNDnyp
7cewChP/7diKb+7Xcvim8vvDtM7Q5kKmQiJ2DXCJp0rw9WgVSMib53st6Hga0C5wphIT2oQ6CjOT
cLUt+jaQqDU6oV8WTvXPamJ7vw7g+bvCgonEJpgPqlhILTRTjxnMdubXTFPvpFUx7doNGwCMXhlq
KBkOaXNhVlFUNe4tWNAuwcyN1S7KKzXd20rwk7fSgOMFJnTCZq5Ymij5lrecR8T/L5yzfpezqFLz
ZAj0RWgmzTFwe1C3/WCvjdpQrtn7moIj12GslUzD0xHYQnI8YClcjAXL3tVRhC/3ziKDKJP7mKor
PRuRZoV19wecGCFzQUhtQy3GuU/4t+w2pZ59ltJ1by++gTnubVajV029muTjxsbnYJA0FV2K2aWT
XZFuCVCj2wE/MOqJ3IPLzDpOEYRZtgQmvu406CpB4q5XGjUHNtNzNLnxn+gIfKY7sfXFKIp2T3n5
qSvRkhY+JD3DD0KQcjdTDIATaTr/DSZ3hp8jZkRXPx1oY79OMxzH1RxwzPHO0kyXN2D4cOSht6Kq
Tk8z0vAmnzX+d5IcRBMF4pqFgQK4ck9iJeoCh45PrrsUKTnYKgGTkkAhwKHMUjoyY4zzIc2b1Bjl
TaoPu2SpE7OB6sbba2Msh8WEsRnIcMzfLUhsjUn/YsSqVClEvW0ZfVEx8ECgGxIZZf65/nJbjrGv
tyZwS6AiEh0ZloyJt7TWDmIP2TgZTVrmd1GbpmY0alaeSb5xkoxgfCMrp0IM9DnMkd2GIwyCAHW9
aJnJwQOvDeiiiFmO7KHKWpd2b0iDe8ugJIZTt2keEK76U0f1l6c0H8pufm9fFCVyiuF66Mn0XSl/
jsqAeJ5xZaga+XJbjVrrShHfSC3x6gLBs6fvNkLq29axcdpsQ/2bSrvxhvQrh1dhWzw+XUd8QyPw
nTl+MePrWmB39Y+OxTd6IcsJxrNb2EkgBWYi/Pl8OVxbrcQwWpNEqcQF8irOq5q5EkKEBN970sM4
LH373vW4QCP8gEYUgAzjuO7C3yjQKSN76RQFyvEzzJPpJzhZAqkibR53Yn/55+CriYE2ZMId2OpL
Et4z/+3kPP24Ec9VGw8Pvx86JbtcDoMsrxWOYcXZzz7zJupkKd7j13h1NjqxM09UNd0hL48/v8Rx
zauvPM5dLnyWY8Q12r3xGMQzxTfnmOmervSPjzia0zRqHVmv5DYiUJp4Djpvnnj0DwryosUCzNJu
uF16dwJH3xuBH11f3nXuzB4JC8QgcxNnmaf0YMv6BnyE/ZhRKuafbnU0NF6FE1sOY1Kh6IThpDZD
Xz05p3kvlv2D4R/W93JswawTPfQBexw4bRpFV0PfZdA6vlZCRbQAiz6pOpl+zyOC4BKbZ02SZgG0
5Kg8AXFMWn/zBaaPradJlwRwPLgDrIq+sffJfGq9DGJ5QsrDG7ubxDBQfQzNbGLI01PWZgAHhyfG
LKGLtr5ybaUdsRezQs/NNsph2kKVwFE0E2cgj/EvCFzCp1QFtc4bDKpJQrJ9B9P2eki7YpWbtKjw
qLl8kvygpQnGYOAPK6eM6pZaCdA1oPHTgw+E6fbhqdTMnNS/TbzzZ0g1+ZNyhIWpc+sBHMPnysyO
PTBBQ3HabuyKeuxglIXtPHcBleaLuWhf8jMSvGGMqu0wso4pfstAgsnKK9Yt87eUvtONI6H2s3zg
Hzotq0MwODRXnAqgQb7cjotu+FPVWU5g60d9+a6aDX+paB/xzVUe/TGY8ocR+zATjEPR1cIUswPo
q5nZCMVsoRG9DQyyXIGfd5Cm4GKLxKFvn6J44mcfCb0VoGYyxC45BO/prbdMSySIO51s0H/g66im
Z74TKrEeRkzbC0cyAnYBZj0UV6QmOYooNlJ8SDhc1MfEhNQvxxTcA0N1zPSe4oKhKLlhyjL9oV1l
8EZVJI+yi3s1n2g/VsQIDpfNfani76zGK7OR41uNwV+QhsrXP5ZGOickGV7Kd38nMIZ1B0Zb6ufs
VxsTIbpTAVwAzpWv7zWOvpJi8Q49kUYGIjFsj2HbZCCNLlRVpZwEzE+L1Q3tUlCgI5x7is5nsZSi
KCaZQjU6/siiIcuJ8SbYe7SDA4DUbS+3f1vcAdMBFK7gZ0F/WrGlp5bmLd56Nk/+YhGZ7Mo7IZ4m
0zhfRQbBAyXR4P5URrTFUm2SNIst3RBqXhQfLCVAwxSnUExlgnhMxmziltPpMMFZYqYVos6NlP1j
+lmXWsNhQwv2GVWgccWOY3cwcPlu6Dmm20pAwAAUgaRWBpug/rA0hKT/5Ny1SGg/776QU3JGtNm2
RQGStEd2SCvsu3wswmQ4Yr6p9Y9rs30Jt/35uLLhqd5J8riKsD2/poVnjWzLYmqnsbIXwnWcH3jg
ZXFwMPu00mi08r1FetI4P7QRXWvrpcYQQ94Li74StV3oqUNYGooW21eP60PTh2hToqDPlD9hMjCE
ODmXxBbIfNXHwuTo+g7ehZMWCAa/2PwDOSjOWwGHLPm416HOhmrNhjZPVTZGdaOdsX+qM/76KYtD
MCwst2y/lKAR0ytWoxG6WrpfHZTsB+dwbWMto6nw5LUeQh4jB+6P+dZaAh+pXNfSkYBtEyDTLA6M
tPxbKDhUnY8sYWYDx5ss/ogxgSoNnxK1tXyBjFgZmITXJAQXFg24y6xsiG6ouGkMvgnQ7lHqo/NR
9o1tHEuqGlGEp3r51v9UJ1Eh0XXko0KQmcOHzqyPcwufPtuXmkxXimQCf56T4zdTqmAUvRIwnXmD
/dtqKnyaqWik09jmdXcZgjExTDdarOS2u49nTorrwwA2Qzrw6aQ97xFIVuyh0TpWlZ7U+Q73pjr6
azARs1Ov2ovplPpyDZZEXH2C/aT7Ravkful7OFzJ7+tNjVwXiPtSEGAdmVh7rvuc6ZUCXc8tcVVN
utAemhOGGnye98FVb7MlMFJxIRb1AcEj67n3m2ojghL1ZaEONutg0QELsdoG6nQLXRW4YqOSrlf5
+WPBylobgEvv3+V5L62SmX+2c27AVM5bwFeQ2zanmacWF/jRo+s0rKaEdjsyiGG4GvJMIrIB9mTL
z/qp4SZm3aVCOTK2BLgC08f1RItp2XXVkwlQvZP5TFfx5xOBsxijKS9072ROzN/x5SgseWA1pK/m
e9rddk4aiiL1j/UOxnIrv635ex3WxLuOcmTFCDZexwWS70UWqbxdhAIRVQz7/UeMHBNy8bGxrfO4
9KxvGmKKv5UbStw0YDpnr8OWgrxplTf5jnWAm8aoCsGkPAFUE50b7dQ8n09qGPrbBTb3VE7DPwy2
jISh39XMoHwG1KD+Cy5PfU0PkrEVX+trv/XWon/NxnmvFBbuj0dFKONnWf/ivfMn+iPyt6oHhgA4
lToTLOL+uTkai/PVN106AdQTuL8VdlRO1COsyD37xKfmKRoH7CmiSp5CdB2KIaFZ1i9ph3dmJi8Q
xoYhFu4WFw+B94GyArbPJ5M1QdgdXKPBzCj7RV8i/oPuI8PotDJMxHQvPGRZQGgzyqTGbV/J4HTC
L0ZkF+bEIun902BIwfmBUa7xoUG6FQGKy4o5lr1IFFK4QkC+S8Y5KRkODesfBC1G9RJEomRMiEil
ViiM3bPeFKbN9ysmlZvvZClkr3LIfVac++pg1a+1s7jPH/Dc4FnkSPLvpTOw3UVGkoQkGI6vno8z
LZZQBnPIauA+AK89ETn6KF0MCy4wFIUBDZ+6hl8ZH3u8vsWnTpSsiQKa63Hi8BZB8NqX+2g8k6Vf
GRy8tKNSaLgPFCkUoORa3PYtCcJFxH2Gl5q4MNbUkKUIFf2diPTJXXv16A7AY9fWqJ67Ms2VP65H
xRb4E4USecsCHtmvXaX57CxcJQzcAomQ2cNBgzHeYyKQAsMXLfIpBsQFh1dB1RqDnImhbw9z5ZX9
iIvkB07OCC7yrJ2A4PEq+PUgT5/Kao2muHET2ubW9iuqZQAQm0qqFPNVYc9SiIuGEY0EFzix80FZ
TXYXvLKTIobPgOcVuqhGETjow196ktNQUVZpclWosKvMQaAr1b2gQDaBj7meV5xlRGU4LblGNouu
SAF2Fs7A11GeLhxkiCORrazEU/aALaduh3ODC9Jw/PQ5mZJZ+1SkOc8g+NSG8jd+/onPOD6zeYno
OO+n1BAgeoP3t/XjjysQhivxmyZSKs20h5OJr5aOPgvp3k428hVlE9eVY0oo6Swc9v5if7JBBuyM
AUeKWl+QW4MCo2dZSkO60TJk6ZlI7VZWA2VfVN8/Lj9R7kUsqwHfm4NiPowepmF1YLHk+vNBADDv
tpR8RB8bMeknzwgmCE2v55HRNq22JbPx4LHp1paCvOez4xOKTEnTkYkdq0mNWGw05OcyQd9TrcRC
wtMOlo9E7Fq8WpJLngTtQcjSoTC5ULudgSMwXNU0wFyyASQBEkoJN5s6VHadVFr566/ui8xU04Zt
7dS2GYJXDwUXAVXb6uQY6DYRCptaZ+MFzwV6vqAnuumJi0tMAhjd83U1BKvYURD7a8diHOmPOQtP
dL10Dtn7pxtKy8CQBCxq9TGsjtjLyLUTx9Pu9tMd1YBpvuKaLzfAYsKMv5Izak6S7pBg6uOi8oPU
HTXhcMCUpccwqV7LCBe7eqaL8WXMHCvWWbO0DEcR/zvugHfWwaibKEyKiem8BaUkvNy6Uzk5nUAY
AkyIpqlMi8U1XyCBQTy35dz0QSJBGDqKI3R4DJg5Pxe2aDyTOYesWipfCOCUpbAivt4yvR+TTKK8
wiMnMPymhHEuFFw8ZqR+hKEyIlIFhUYABlnhXQ0+4P++IJsV4SjPoLC6OCR//wvFFCLs1PO0dFmx
xb3INzJ7fsPB7YtA83E2L9ylOLgp3LYsQbdfaUBxQTPzawT3zGKDNgY2mt8ZlNjeTmHWzjT9CWTp
DdOwIzj0C+XlKE++VoXa1ftcwwCtUmzOPJGYVC3vOYV4cDGCgxKByG38YNsDr7FQPhtiDvMVesWg
z7FveiPULbk+XgzBBRqRDdLGE6k+TmMGXJqgJ4HLyJHHvjRuDGXJEWWFwWuFHNgoRoQRpSIohdox
MIQTrp8LaEiBkhLLl87H3AlsWNyOfDK3m0XoQg+uVgYby0TlRUBJuNTzvlYqJNA1RkowwWnJ1Epw
czO4c4PV3IbaRXggB71jZULsOJGFFgPCK3yTF5HfvH2dU8B/7QBTLA+VWL2W6ObOPTrGc1j3PzSl
evLLVg9px9gPUbCSifun4so6f6mLYKPBYCNEspn2+K65sJYqO6m9x1Z2IXkarxBH2P5UDvOA8OIk
E0ttqhmHCfNzLH3ihZH4HXcoohCcldUzT3IX2EWZXiurqdJgG0uWbXcoOsCiauwmW3kkK7oke3Pw
k3I2UpbdxftxJ8S7AO7v/GJeJU46fjqd/Uu7xqMD09Gu4Qd3uZIUkOpgBdE3LxaNZvZuWtpTge7g
RUgs1HOkmiacUYXmW8F9Q4pYvhcQ9hPDMAgWuKh913/vBtMnjSuRA5K4UWsiQJ7LJp+JqUQD+xx3
MGfCIQyaXDKDrZEsf2IfMy9kyrxdpFY+IME84i0R5Y3yo++emBYv5zzoMyMZpDnYO7tulbDSV8bn
PFAXRJJk6LZ7IiijeV8V1PZAiAZGGM0xyvaF9EQkW/+uzB7g53bxUrN2qLNPZdw98hjoaNpjzpVM
Oq58XW92t8bEva2AHVaN0cjiDeVIPyTdWODMPDWc2C8rvoxtmE13Gf5jc6QlLWfOFi2dpIq8Jwb/
Q91+049ubDZHSBA+wXPFUdy0aYLQfW/uJ4M3DNblHB215xY1cXCaoUw7uaSdCynLu0bn+XMqmh8K
zQi7ULu63TDcmbYlfotp30jtMxwycyTYgVv+oxOQaCqjj03qi3XM4kM5Cdsz/qiAv/u4DRIbkWbh
xP2aXLF2ydF8luGnuvQQNzSEIcpYp1WgVOZCjKbaX42B3Xqr65Z//gzxKWLXXgFxUC7Ok5XzQrb7
J9apz+L5uOp7gTvxA/uNBxrDNr5mq0WdkeT3r34u6xwgIS2M02VLOvnMyb5eGz3sKXwvB6wGJszP
aLmsJzqL3QZqeF995ZzzC0ciGFRII6Dnu/Zl3DryjHKFH727nDEOz/0MAo/6sOwdNSGWPiBphOAo
tpnEPEoyu7k90xUfOXd0pHcdmR80hOzq37Nd46gxi3+WOJPUFqV4RwUx/EonNAG/HaQjCsG2g1Dt
IvA+fXZ6E9JTNIY6TsX+ifbpX1twOAuxIo+HatgaWcf13NJ0rFLlYqt3YVqumA9tnf8sVp32Zmp6
gy1UE9crBPiqclieEHyRerEf+5wnEX07BBW7AcWs+l+LLSbUAN8Ioeh8wjux1yBSbaVREf06vM9t
C3K3q2QVhIwf0M3j0SbGjy2IhrTLKAKQKZf644u1JlC6Pklh4prNUaB6deBQsVkJqT0a+gF81c1y
ZnI/qjsZOyroxHhrC0qFD/Kmz/jY39ZsJwkqoRVUphaUEbEheHfyU0iD3h3oldNhjgHndITUu7ld
CFVyKHD9jdb5lswXaDiIl2wlgU0oQ2C372NF6SBOqMKlwwbE38YfvApjMxV9JMeNfYdPM5VwrOyT
MktVlkLnC+1yumW/ARzYRj7mFdF3FHgPW/976L7gPwwMd6VwrO/ZOx7IetCRQyXzY4A+CvRowmER
ugNeWHByXninmgZmyReFcF/oUZhNH5hi4VIE7wi2Sy+YXQEDfKxGOF/WLfMotC0rpv2k9f74u4ie
nNvYwaHvzEKJqc5bNcSawE9BD8IrnC8rP8N6rVTcblgZiqNBoDrJbCq9c0bombjbGAKjcGdDSvIU
aOTk8eBK7Lm/BM8q+2dhboRuIfGDzWXkWhrTzWpj981WuxPPxoQoehe7CZRzW/3qOizrQWoC9WHY
3QtuwjVQB9F4B96JfMPuwZV8deJGxAKYcQinu08u3sJiC/Vc8s1GNdtxo8eAAfa2mKZ7vVpjJllf
4tmCyfYqfQytdByL6W2l5Q853DR4ndSd1NDtHoxzzwCL/yy0aHF7UdxVp9KhPcN+xkfxZWHdHiyA
qfmCqSuoIGfckKsicAjcx/YbiEAnQwFy2rNLDxjzAYEKIcgh4NvSROzjUcZftjkhen6WRbb1o78r
s126c2LlxWWdS40T7w6gsXQ7m7oxk29ZEOd70R4HVBxwTqj4FKbv9FQ5aHfBcRrhnsuW5vpsunLM
TPx6RvAdLRMJZa/7ZlSO9TLEyyQJJseDHnaq0ZaqIzrcy+UYtgr8M2IzmF8C4SRa+3J7ZxSyxGdZ
UiB+oaz/Pkj/7sP2mmoSu0Pmgu/ksyvbuPUimWa5OsyuYkiVKld2MdDlIsxLxHmedWuoFvLDDB/f
vo1QC00CWnsCdEQw2yZ5hMcuRTPQG3Cg6b028hiPtrzffsUT4Kdd8QQS8TPD1qxujbvBqhdYgtT/
mPgSO8zT0sWDoPtu1ayyGQwJMEdKo6VrfTGE4IiKrH4f98hRigyBIEhZiRmENaTnjFv53uGiCvku
lBK+KPbpxcN4nxliqU93irj1huwBaPLUJwYC1cMnXcjNVvBcjPM/Nv/2ZmNhNE13+Y+fi1Oy/RuQ
Mn4c5IfayZfRlJw+bgzbX9SKd4CSn5PoLHJ30S4N0Ja+S5lKlFMzFR9B16P7dq+MP2hytpjEBx09
0AiSLr7B3A0wzwF04lUdEi0WZ1fpkhYDqzj1bgF/S48w+b2VfZhkxNqN5hvDm7lwGedchrqxLrFL
uLSK/wzEaq1lAuGRdR1eCt7s790+Xakg69bqLdpC2z+HlsUIaIf5ospw2/udqD4DP4SWTSX53DOi
ZEtJ+Ir1Wh5+C0Zqx0J1ooCZ8jeTHqPgWWDN+AqWmnFJQv38sQocxuUVIJz6SLcnNX8/M84tJGvc
2I19Frj0GJ2HXG2PGFgVD60ZZ+NGcA0N6dcaVA30G1vLUt638fMmgwQ7CqVJIfjDdXA5yJ0ze6y7
JXT0c/a9qXLbIBkhrDi/7E0fjAo2ENWYd+cQyoqungJfAwKLhSlAbys6myAO7x/NIDWAisIA0L/V
YphOM7Ls6SynbCCLk3tNbCMaZm0+76F9WfKtlhlb6gw0sAErzcoPD5/r+lUZINsm2untSyGmm5mE
PYkneGYscMerVv/tzRohi2OO91/wVb/sgymbyhj6QXOv7zklp24D/WzOrG+WAoZF62zEN/7Pc8BY
DyVy7FBHGcwxliMjC5qYFN3CGMwcfLfvWerXAbO3PIhAIJAcwDOMCWV8wgvzjWXATfGKMfzlve+u
XbShiWQPp/8o1o39HMkLXvA9PeS8nP51CJ30w2Y8SgZ75GTsDqcd83Grc3qyElmokkOsryzkzHYI
DbtPXCvq1YPSVxgcszKOaNbQGX6f3d4fCtqFCZY4jgNs/P64P9YpvOgMTIvDeR52PlYseGIb57bq
VeZNUTG2ufDaJUovTrgmZAq1E9gZNOZLNFt93jpsI3Vi+srK+zLw8YA9V/ssg1OVeWB4lR4pFvOZ
WfQLfrdfTu7HDuG/NNfg06+zp1gw35QjlSp26nZKruVH3cgIkcns9iF2KrS6Ux0M2+vR5bkSM6hU
IqiC9j9+U5r5YoMk9pc1tF//fSFKmJSdn9i2UxbdeVh3WJBQlrvFCJS0wpJ99RDV1mDRMNs1AiO5
tAw1VRUNwhqhclhNI7jaarRDP2Ham/CwU4nuO++EfDE9NmZug7rkcDTIpXeKUQ4AR8uxHwzUHhtG
jz0Mgevyz7aA8BFHEbJZRXIvXcMnrBZD++SYWteTNNj5M6t424sTv/oiGqQesbIgksdxIcMWYqrx
46SEAbdBBo3YzRRNMJNAjzxxp+E1UALsp5jd/33xAU+IsmY0331RHiNXUeA22Zwn93nMRiwkhxFc
q9yvdEFndqIyK1BFxTKj3PiEVejqMyMW01Zk62tVMaA4J1mENNkCkgqr9ArKDkkf0cUMvod/Qa1B
Uclwhp53d6IrpXQ76FC8pkJu540qiCWVXauu6r1+HCWa8as8g9Y7Iq5WBGgYlIK26xWJuqj0SELW
pJffxmSRULWrrj5VXakPIMHdsk2c9SCaM9FZM53DJjPiz7ZTuYwc7IU0CORFuZXQ7RFcCGES7nj/
njRE7r+MnybRC5/muNQuJdj54RnSIgAfl5dAAMBTVmpvy5o1/bEfKjulmPwX31vpn+WQAjzhgBtG
wxhG03b6s3pZJZ1w/Q5p3dYD47+PH9nMn2n1dVZK+PuXbYlDW0A5Cidn1xYWT/ZoRN4r4HM1fqCN
UZ5Opu02iHXmECwX29kNp3bmoxfUNf6mflY8miMEXwdB+mSocdKU2sFv8YaXwMCADvELZHVrfjVD
yhi6/toWoTfPYPoSvM6RuuNTykZBtTukVLC7Lyatrt36kehncttkoaAoCCOswAbeQZKfMszlMOyw
a7Ju/SJC71ZhHct6VcPYVJlQGfIzP9QE9VWwS65JEtTYk+Cv7UGu3kBJDMoc68tjQ76bRzBENwjz
hyqbAIIT6S7rabsVjkxc4DCDYBHeRfNmywpdVHHfEVEwd/UaI37LKOAcdJcKye5VwqYnbEgafUBR
uI4CEuUUFkUlM1C51kZMl4jjBI9bHEcjHXDwSFKzJ35FMSfhaUtIdsdm9S2KfLj1cK0+qUpzaYvZ
R7jruZyn02bFQVd1JO+B8yQndpQW2AKvwPE4VN8bcDIs/ul5MIcHGRywKo8XG88XsLMnBRsu5OnE
Z8TU5BN+riRvbRGzEjtwfUJMguCdRMsLsHEI0jvXVK0g8gRGdLrWR0IMA/QWFlqXJWU+jR8QwMSS
YTlO1g3lVMWfA7/QuHB4tmr8EfO0QyXbP6LTndi1FlGud6mUHAKfDlFNfnL6ixOq/493eVAed6tv
xCzh+aRRhO9lQq+XcCWaL2q1XnhWMC0d6KINjxoO1Mh5SDcpsse/HWfoDx4N5ZxqxlerVDoARNQQ
kB7GGIQ4OdlbWvadt3SUBkZFfZDLmngQQSzCnCaMN7QNOWOP+WntD3x6UeFuQPoJnYMBupeg9tpy
4wvMkGx8wifiZHLUExaTguymuXiw/Jnm21MUapjk6xEGe74/K/K5jEFrySArRn+PIUNOKIGPfjGJ
cXQPomjMFxbZ6ZuE758cqg+FNYCWBlipjVpuUhZNlgxgqL0FYTh1uWeSjP6J2G3HpAoWm6N9HBii
N6D+AAJYaQKaYYjyqaUE+ybJeON9XFNLPVgDQuduV04pSz/Py289YC2om/z0VW4sG1xiMYZElHE5
/KZpOyNbQulARR294G6q6sduf4+0rOEIX25WgYwNf13PU2MU2WsFAH4r3IIMkisCmykJ4Y+rYsQv
IbU2VJpKQthgUsI6Hb7TONP+K0QItnwpJdyy7umllFqmsBip++vEetUrCApohR7klKvXm2szG3Y1
YyIfZPKe0NKVFteHjsfct/YsPFjSdKSP2wjBA7ipwaod7ZUWQ68m8M8RZE6GC4J9kB1KZh2MMlBf
N/bMruxKpMZmL/KFvEASV6/UUlpi8hbYUxoTpJz87eHoDPfNNblkeJKcw3LjV446XW6QaMtB2No9
2kEgjFYYN8ywDR+IspN/9SyYK5BQOH8XiypRbEFbaVwtI/E2zvhMOcDfibRa177xWBlvUJiIKgoN
gPTCGs0RXQDQK4QIV53ir81yZPMWw2okoAmD/lX5bX5HO5E6Dny5Lwn+IlozuddAv7U6aO24JrIo
UwyAwI8iNUy7MlG9wv6b6mhRzVRZAKd9R+9JKtrLcrWZW2WHXgePUrmsNMD15UTrYeYM4sfUu62C
9UCzU7SjIOQkkSJTcGsn+xbCDsr2WDYemBOYxsI+XWecqHrDBhW+jQUfIBqZKvLH57GiGZLMYfvY
2oghW+Vs2wQKMKRtegg5PKU5hEmdGx6CmaDk1W9I6xT98DRCGfmJvi892FvGLc+upCY/kSo9ZsUQ
Al2yfksmp36EOgeEFwBmsUux2EVbdiWUaiqF1OpiZmcLJlpeN/vmqjfSiGYIFcWfoesKpN8g9HMA
KxE3lL3zgPd+PoMmzfxiJ/ATbYUzWRYV+9/n4D7yvt5Z9JvvshkYJH1wwiQW55KJyYGpSAg6kdyj
0nTZ8NBlCuCt4YKkFrpHn15aitR0oArxIviFBp+3JW0zS79bwNmkrqT9Czt2NI/ExPGkl5aLNjUE
VLmMX9gvoQ865zaexKMGtHgrwsGKS+hYkR502Bt3UH/FNGE78A8wOkhbPNhBPgtfOI5VQS0pcRF8
/uxZ9NfHjb5hjFtnY6O7fhDRJgtm/0npNIo9ePIRocJ4zG4oiZ+EaySLif1WlBDj0bqHIpUmTQFn
ktXmVr1sEW29OE963mnn5+qXmIui3V5k5OCB2CS48cnVPtSV0XG06Mf9DRyOyPlaVat5c9xmmAc9
5S1QTjpDnB+I8QBZV972ipEgBjRvFFOCfXPLWAC/cW4v+v4ZVKZf3Js1M9LRjydNPDhSo708nfLr
jDlZ+VGkw0tRWsi+vH8IkU2urbfVfDt2kYskQwudd6Jlih8SylRuAJbn02znVEp4B5EPM7rnCPa+
4el1l7P35Pdvp+x12SysXU/Swa7aflqXi5hBCH0a0WNsyWxiixUE6PqSq5lZ32F88QZgfR1B8DjJ
a1uUBXdgo6/yjcWX2uE9/EEE9sGHsA8xN9AP/X4hjw5vxj8WnEAZzpVv7gMB6EscRrmH9M8oalFA
04LAkIjpm4t6YBgEwDiiiNZFJFmiihWdrhrk1n3yQWUbDdks+S7VS8y6LDGx6kj/BbYSCjLPqJlL
vxOxaJ4eqn+IVhNnCDx3Tk+7aEydChgtD1ZE+OUoC0ig3CrkSPIESJJ09pS0Qw22XMz26GgatF+d
6suI+8tQdisVGoIq1BcPT8ytH/ZwJU0Yw8SujRtzn3FJYQYJd6eKvBAQKm4/YwpaNhL2sRRosmIW
Aq5OspMM+KGw8vIZP2GKbJm5CE1rhr43OLZIO7d2ZpW7TeJQiMIy1cOiELuArmklGioFZagnQweE
k69Y1KAWvv7FT3jIy6mW7MjeONSR/HO+kgP5z0TZBdqzbQ+WvUnO9LqwvKP2/Ws1Ur2SwTcmYdzL
m8cjpdGDNG9uhtFBtjfckbFFP7csoBxtR48P5NlnwBDFvqsp1dtHH+2jvOrMCUMUjUhr/yIBmA7B
hEiR6T+OwKb2XFNY3qR7afnlOH/Rfc5GDnJ/RcDpiyY4M0lqBRZm7YAvnxdjvXJf3Q+1mz1wIcwu
lLrVsCAlSdQxBVEhGWEXSJOX/TclWsabmJwByPR9PCJMpSJFuyxjb58vNXYsrd1QHc9Hzhpscp7m
QkM8vjWl1bfO8x/NKO0sQ0KoomYavLTJGKjr41XXLPUFKapnN91d2ELigNv4iIMxmKVFFctvrIdP
XXnOHvjbk0xtS6/w+gcx2WVwke+INNaF/8A8HG4azXR/3ldhV9/43OXhRbxLuIT9pFNHLQ4SHybU
38M6Mdyccg+vWFfECKiMKT1paaNiovr6+w93wVwuUHjbLQkqrPHeZeJPFBRPqhLM3pWoJpwHxkOn
EAATdgawIaoOdaWG0/r3iOkeAYjm2rpLgdzwMfFXIixM1hQf0yQMmPrZ5lWMrTPgvq/C9k/Bh0/r
LU1o1V91fGq1rbq1kPx0gxCe2zb4TR6+GtFU1jYK9DDEPOP80abDCQsUrqSQbuCZFfiPrx+zIMrU
itavrB/6/vfMSQvdy9NxABBwoWc/QRBLlisu0ArmsPhxeTZyPwihwQsTeMN88U+eZ3uy1NiA4B1k
VJTJy+2rY3qgt3NYxIFzRlWfTAQ05o3szUw5k9CvLC5DiweezRFuui+9yTYAj3imWJBu7rGb83sv
YKYZFHHcsWfomC+E35BIfsYZtGFluvTrpPgMv1ZLb0Kq5cE760t9hHURYW944G0nkAhnp85dXEVv
LvO9ucyf4G5gDRRndz+7wz71oNR9k9IDbBghEOJNQ9LzD4HDNzigROeXdug4jdWSjth8u2+4CWli
J/NBNDEVkRzfwA4+gLAZ0p1z5pTG+U1F/wK7hk4cKt97NQy+bIvC/ZzDfla08uquilhbqpeVMtZV
xXrcBk0lgzSyi0VEic7kuQw8SJ9YyEtOPBcpZEsUQB0S42y0BerDJB+9TMgrG1wu9O8NY9/1S5t0
6oX48PkrBt9Xm5qPgpJvydvMqRN/lnv8EwPni1nv5AQCfFm3FaW+UjGM4q+R7TH7ZOwToDp5Lmrc
gcxUgzpuio8Mlrvn5vlANxYxSD4/m91DQdtzQXmgDWNhUMg2jL9kHF+bSIFX+zSumJr+7HcUMMu0
QU8Ec4QpHq0p24L64RrnKiu1L19NgdIJbJuNMAoOYjahLr3jkIaSYYAyCXtCzlvj3XdnWokxlO52
iOXW5kheQ35WxF2Mn9pO6YAtuYyvfae9DSyI9y6t1mCTFQrXsIKP4md338gv6HhlctAHNFH00x+b
S6c5KAJl6UTC3f7PHk+1qbE96F6av5ZjCvCMa5BJDLh7EgC8HuX7ECJ/hzM8Z8qPbFk1NJ1S/wla
FdrsL8iJFhkIG7kyH8GpjnCJCLZHniWifDpL8ymB+XEfP1JZfiJjmX8sbvCZichi+mrTwz2zUZxE
3aO73nj8zQiGfkWNqIIpEMAXhAKgpQsg8glQSrLBwqBXwCTohAXjJWLvZnXVsKpVGsH4sx4J629x
Lko/YczwdLRZFMlBDxKFo4xSBzg39NKuyXf/Go73CsKRdBN5uhRnunTFAOwa6xkyuIkoBy3BJlrb
TJdZSM5h90AnG8qxVeGSQP8YUEEiwhdNdVXKk95gHOn/euKxPBLtBZaPP3gvwRCeWZRUo3JcA6JL
pMNwxiAALwruNC/isQAcVB0Byf9s4urTQkMy94dpYxeiNsBZKtBsg96h2iyYKo8IuI/ZZXnZfT3L
eJ/M1VUBwXG1xd3Z3+qQuGUlo5UZgHo24rmt2Yu3HimSKpXW34U/WyfswcINnR34Pk7d2cXCUxOn
7+kRK8H2QaED1w4eeFoDReMvst7g7Wn6cElCl3M/oyBI2lAziYNLCr8gL3yI/iW5KrpUAQd1ndX3
dd7cmmedr00oDnYVn9gYmDi4gl9aIpwP+RcFnIK4Ktf1FEryu80gDKsZM+hmsw2q6M3HYOdGNtrk
IuMSLzAKngFuozkZl44h008MhYckWolA37rh9Iox09Vh2hoIuGrcUEiNjaD7mNHC+p/fiFVi6lrH
QNlTvhgA0gnU6tZclWM6hLk68gUbiKVbcfyclWeoQVy3gR1L7IM5+bpP3Y4XTDA8KYYU5wdUVD1v
VOdAJ7Y/xLwIpTFHgOYpxsAlro4pUKfFxYrLkpF6zdt5ToF/GfUyiClkgbRlhWNV2ssJD5Wpz3Sl
4IsMSRyDHvB6tZCNG+v5Njp5EA5qO4tO2Cv9XAxsgb8EJ3cF3fj1TFxyx9q5ttXCVUF8R5KNv3Z7
kCR2diIge8GeSEaut73BBqbqD7oR4TIx0qEHVQiznmeZdAD5rQb1J1yd0d9iBOWTIdT6DT8rxEM6
DbhCWrlRfWUGlGc2lE77/7QJznAxdEBiEZdx7O89Z44BygijHHe7xtOcp4nfZBC5Tmw6An07WB6x
OcnDd1dX76ABBt0n2Ap/Sihmk3rIxMHALbqBTsIgajDkH4xxWBa+epK+bd08Q2Yz0DWpG3Zdu2qw
sVj6fs3C6JDNyrSRxMYWYpF1cRV3AnkWwgGMCvfa57VDsXnMAnra5viJdKIwdCIDsBoU8e3xyvWc
CbWs/BUHSzPi6+UA268rtrsAln30lWbfeT/oTyTX4oVtgwLkJ1GrtUPyo2dThndWgfl54YuTAlu4
oXh5MNl/DWSZCqFT4BL5XTHip+e/gi1YI6MkUEhqSlz3L22Zy1Hu1cT36XQm5i9H2q833MugWorj
frp0SkYmoaRBbjclTBKaRaesEnS+6kbi2GVQsBSsxotVBJXJmt2VpGlgkPoF+lb4brwN8Yk/V+we
qjy/XHb4cxkvp0gUmNqz1dpZAaWXtVJivjaeD81apV86/JR62NOrs/bMPmzCF1RrJH2XpmnJEPQ7
rW+mYifKqtQO6NYFM9EStZiBxghvw5ud4OSarhfpPGRv1HIg2FPH/7f3mDqaZSVeMfXF+zOX43oV
rC3d7Tvon/1wy3Vng5wjHAwyEZG5oHAnGTvbhSEp4/3tROvgzqi8e0B2kj12O3kbofjBixSBygqM
B7BTibvD0FkLe94rlK+rJbyJglSgX9BwIxs9JhhFbYdZqLpvJg8XWNfU6js2xKFaHd0cvqTTbMHx
pgP8GFcvoxUZT+gnrYi9GGEvW1oPzRqIxQXjqatj2Zf7G3bwOQUYgkqeDGiRARUwq6V2jmCQ+vQk
Qk0PbLy4G7tqp5XxSgoTB+ypQzVhwVGLG3gF1yc7K2/29nyiLKrJee+Sp78I0RR+BQlIVlxpUZLa
tSWRWEJB2qIITCWIBOr1LM70p6Lyl58hx4E2Uv0hokEheJzSkOtjThOpp6W8gLXEJcTz0gXb6y0e
HZakkJ/O5DCAOsSldFGHjNgty7laUqCiDk1omyaNgtOc1ePLTQ5/m9cVwUQyMruf4v3rsD12UUOp
/x0qIBnjm7NcIUaz24s3oydEQDkt9Rmmq5/MPOw1TPcsNFowWfJKRBjG+eKAxjzjZ9x68/GMRquA
7GMTzSFvImXErXqZ99KN5he9+j4+LZQ62Nx6guOsC0emMyIEHKCQYw1zLGyln8uDYXbU/rYHyuq0
LNHv48gO626NJiEuwZhuAJkWSzK+wzdJQRR3WX3+YJdXpNlTFsy3oMYgFFud+PZok6oY8DoCISlJ
WBj4Thn3Rg0dsra0RdpiMLDQuM+mbmENBR5pMdVMP4Z9ekR/l5Y2RscT2bLXJ+PubG01jLQKaxDe
vRmVlb20qNPxX8bjyP4oCby1K3Ze5HcGDIMOcym9oAC/oY9P9FFJ9v0Oug6J9QQGQ9gkiqPagX/2
ymzEPK4X9xiWoHDXPTyWvp0Qe0kXo3fo9W/Crye6D4mZ7SBPqX7yK/0EpIDZpYyuF+59sqPoByp0
XoyEhQ4Yc0qML8vH7rxnhk5XHD9KDe821SeJW0d8lfQ41eXh0wD18+KD7iTZZet0+AG0KCFIkBdZ
o2ikzBYN0ViwxKELz6DImoHey8anEsdG8v1qufICOrB1oaOTn76/VM8y+84NRYs3bK2ZQzbpV2JM
tUNzB9F0ooLhDTaDr9xvfNTCLnFxUNtkT0HwT+g8ivUpwE3/UOdHSlsXR1Qt5aUAacDE2QS6o1oW
7WYR2S5D4v91EAXeOqsFe9VVCQZjccl/8U+tOGaN9r55N12VpjInnXrQbxwg+bPIiYK7a1ySFXHM
qPnzTqXlYUbyuyUJyj9QxvXz9b9s0AmI2YKxNeJRczf523aGoIi7vX6V5K0+lrYxneMrEf1ZrhaK
evFnz4QoZmNMrNG76zBdt5sTXWBKgoxhog/bt/swipab0KF2l9BdDTf2zlMVCH1Ksa4qEiJWsNpZ
yGlbG1A9nBZBmsEbwE2mqetzhdLQKHCtNde5/dz/eODfs5/2RdYrt0xxKwT/BAOaMbwurnIAf3x/
sUcLjg03HRZ632LYHbgqVt39wNGsdJeeh8Ec0RK6VmCB04NxzahmAHlKooxW9m5W5CGzrqaz27hK
cbZHL69U4a7J95lQHVgKCrSSlVQqOW+bujxu8WuI0XmVcp0Smd3H6HNpqCLt69TJTnJFeKuLPh8Q
BG8s+ZwMwof4C2DC3xY77MLr6F5/08uD3XTe4fmKgOPkEL2C0P/TIA5JORgc/Ov4uJ9QoCp3ullC
i8bKYadYAfAW6GTobNmft1m+wWNHtDdWAw/SAdHJ0WCGYKMOuXnDmh2udpdNvEF4gUOxYlWdFqc8
vxFPgbfIzQKoyBFsJOjCMWQC3rnSVkWahLrKF8tEn4Z6c0UiWztzr8XY0l05gaEsxd4euE4eTuMU
QnPRCHXmOyHZAm+x7ahtrrpB3TbYWBvZmKJk4hffOZ9cdrcEWJV+jNMjpb+GAz01xYY/AJRcUGgH
TliqIJelw5KMtwN4/qF5pYgFU7CHe4050xbuge2dnSM6X3ClbOlggdFuEvKlNoyKRPnu5I9irPhJ
WLG4W1sgXOjMH94MHhcCvGEktrThfXm2f7BySnpMiHkLB2ifEwdWzsHIQ1tJKyEjEF7K4UTr5aQ8
p9fqABQBSSPsfbwPdRpJaVakpOjhc41P+0lhSvgWEg+LE47VaQum2KMJnMfuQRGKWYtJWXAKao8f
5pt2qTDKnfxxwHfRuBIRiy0ItnDxToxY5ciT+ZZcXVil6LMe0Lc6n+eCeoL+dy9YmnjfvLV69yrw
pzaDw0/+rGo6VGnzDDfFIhE0SLrKzgiBwPuIkvdGUOJOWHwTjXiYNPXfkH0zqaTPnIonqJ/aAPYD
fZRKc4KEYkVXSGMRCQtEM5qvyRM6DCODoFgy7Hc1BZI5ItHyVLG++LGrtuXkL5MuWfNLAGSvqOFZ
r5bUP4dmn0MBFONSO9+xcJFM8ke2huNR4z2+DPjslgB2/6XS8hIACLdgKOWKA6nc7ZLwK+x9z9lE
g/FW7ptNA4Hddmma1Vdrcf4SiZRfyfo1lVKhOS7V/oq4aGGt8AI6eSWM+gA7Gp5u6zQDR5pHNSlQ
htv08DRBXXX8RNv37DGifr6qQoOuMwJTqQBZzCilzpo41SPNVr/tnx91GVYeyZ/1hXKgZXs0+AUm
iitq77tBuI3CnjaOGwtGYAw5+GqSosoSihMSeOJleWEWQvGuIRpz4sDUWwm03zCiYpXE3vqdYvNh
SEehYXN3c+N8AltBo9Pu5bnkydKIn8R6jyj4ZpJnYCgOMTAp4i6gQJZe8JcaOLv7wjlTWrKwaGJd
iuif9dmF5ueLo+2VlcMS1e4LCG042BBZYoqubBt6EV4dmir/X3z88kJ8bz0we6DRwl+14whDgPyJ
jD/UsOn8Tc7uRdi5RTRspPWthfasPhMty/6qCj0lTsM8i+siJMar6VU9YagvkeDo3vdDRghPGA06
v3Y+/uGtWzmH7Howa39gy85UidCP5cB5fec8y11/YWSVaaapE3d5hFSigzh7UmesK3nWH5ujSIZe
PNYjOnCL8etR1AqmrdEKSTSWkV0ZpKEJfTURncXh8BYjh4fLpDJGHyOgR1ZYAjxnDBIgh27flPUZ
WzxhX7NxMM32O/e1vrOhukvrRqF+8e1vwXuFYnMoJ2Nk1nmqp5IOmb+PhysDFPFjCUhr2KwE9Kgm
SpyM4pRX/dbvJ2ScDlvfsgkSh8wHURZnauQ+SQ4NWN88B0z/zqL77feqvHMOz5HteSJ0SyA0PZsv
/a7dHGrn1n3I3NJXBS0dR2mHJCSGBkIzuiGjof0dzVJXEiNWqwI6GqUbX4TT4Uerhj+9hlH1Q2JO
kH/AOzDqHbhsxs5LKhKFjYjqkbMdMGV+SM5XCO+ktcECn9Nt3ULHHqQ0XhJXr6/F/fDjeg/L0CyE
sJyDsmWJY0V9hLL9I+WFk/fgHykNLF6Cv5WiJH2DHHVY0duV++f1DlLgm/GKGEfUwz8L9aPCCv3c
6oTlMT66eTvKehgs2NeMG7+71/If9WNo9LDC8Ge/k120GtG8DiVSDDUlf6Le9Jkl4dCCh+MUk/Ll
pBeueIf2LJ41nfUj7lD9RzueJ2NjCL7iyvSoIlKA0uFfkXWPbOnNVsNj1Wt0ptRgfUGZbnXOwxdf
CYzxP9XUiNN58MqO7ooDnu5b/pphJdN7blBVZ1VVdvmk5uq31Geo/syc14ofet8gXCRpMGwKlXiq
eFLveYWNhN1VelghJNwhSO2zNE/AWUWUW+3FqKkUXY3C/P4F2atjfC9F73dJpu7ODo0H8cGzspMH
qN1LB8ESEpJZTtatCU4eVHI379W/EJraSo/j3NvvM5mdmiUxgRtwLiEnSmZCiMgvxf1Bal1WWjys
ldF7KX5UY9Nd2hpslzGY17NDg6tf0+toWW3KpEcXJZt4IObl81wNPCTKVyidO/67lggbuOy9yzK0
KdUPUlm4MdfilVt0pW1OuD39AvPaAyM4rQt872y1vy9PiuET2A2TNsOzrfSmAu9sJFQUbBqpcCoV
DzuGlE1DUSAC0ngNeJK3qttQHFeOu6Zs1D/If6vE71lQNp5rD18E5/cPvaCeRbLW/4opeoX0lgg9
e6BNq3miuvEr8KC/Thry1hZdU2tR+cnB7/3o0oWtQ0LOk2WMlNuqIRfI/8Nw1TccKsSwpaWAaCw0
Of54IT1ijACB5NZiTAR+8TLjzM99S+U19KzpdIaR7FdNhj5FcZYi/e20h6JYUrsa/fMhdA4pvcjc
IsPs7ECxLiQ5w3DBtYuisKmwoDZp5RrNwzbkHBQwC2LFKVLJQBMYEAqwzvc4eR2LUcMnFPsMRn5S
ETvA4l4twxkuBKiz63FdVdn2ce8vdp6zxcgUbpO3olaN4Yq/Zh62JC/1Rex15J1+5F3lg3yJN+EM
fyMeHKjuBCKie/ZNIcgISVb9WUzzMoL3B26B+ZsTGDkWrY1D40orQBfDG1Z58Hf/eaX3WovIpoXd
NteZgbLIPmoxDglDniWQi4do4n+jwJonC0Y9PaahQECUxvXWWk4K6KE2LRUYC4x3nGPx0EGjwYnN
8B7lIX0e4zNVbXNai3Prll88spJtGlzOLX04d7we8NICgysEM7BMqMZwbziQeNySHQ45sSVQeo7B
7ee8+S1zzaFs7FNlBxS+DlzU0Ow5CedMbLj5BQW/bzDUZrKp/l8GzWtLqX4unjWi47A3aLK6xooT
QlicpGAQIOvtVEP3BI1V88NuwAHlQLxUT2hs2/9OCKy0XfH+ghThTBMGih+q/UfH6YWSbNDf4I0z
F84R3JYr6tatbhASre9NyxA5dxAKYlkU9XMhvb755BmdCnxJeA0hHsHAm8n1cqckx6XSuVUbKqo/
Welz4vLctD6EkKD6c27aZyLwAQjrveY4r6CvcjsHlmhx+MFq6sCwdEfNwfDWWl2FH5xMmhhdYsNN
vNgbd9nORBleoBjC3SZ32ihyavq5OSPoWFqSYWL5auQCI1GNLGumTxMG+cH6IIuAv8PZpbSmJ/t+
Ca/vDLpZitkuuwSyLpiG1KmW5BD8YupGtAFxetR0Br8SKlt2l6kSUCUWeOzgwLl3XicrDTNhm1D9
jhrU3bzEcwBvFdEj7F0+hr+eP6kr2bHpoOcPyotL/IUPabeH0ubPxkJB49WG9WInvNyckypd5GTD
/3TRNFVbzV/UqxPP6wMX4C9GpgYf27g//ALUadT4de7ehe3EScGgSXxY8QHiuG+D1QxmMl9AV8v4
maRuYfXT3KQ34I+FhLx/mNHJ+rcrlE3ORrLZ4fziFwkSSCLzd3M1IU1FDIra7SzEQxMPYJT3We5+
glT3RH0RSU/37Klmc79a4ekNdqF35vlE+xOAjUFD44jrfxRuUNcBHsfS/2xqpIqrD8ypkjdpuvtO
E1xkE+w9gOn2XZeeLWRbo4hCNWdEzAZGEttpqovYmGyykZrKFTXqGaFiXrqzYxj3p0ijuyAwoOSz
+a1Ykr8UZzWd6SPczvnYOcVx/NItTZU2qyL2VOwz1pj9JpEpYuq428SiKBGh6Uc85511aA4blu+g
iEEyOrZvt3k3F78dHkf0sYThozAmVyp6ULRKakh3nMDDKOUxrwvSqi71i4PhdhMqpsNBuLAuuM3/
+LYS/xohrqNFl0EWMIOeMdXOUAx3GWkjBxfyWgvXAmjB3cM13j6WbYHY8cuBYSvzOkBWFOAO3LZV
x8FoDHmG3H17EKCFUrGrPK9bPYXZBWsvBbMOD6/HfnTeGBVg5ivG/NmpFyv2tS4pmk2ovGhgRvhr
7iry6LpOw4mkRP3Ns2ffvTLJbEQrLMJKzCfbLBLfzeVsyEXFsuEsKDfs4r4YzGpW6h2ZTBYSYCXS
nXI8tPSDHgsL8QuTYFBt7LaTVtNSlUZtYulh6jFlwE1n1bRx4rLI00TA+STIm959S1BDAzNHjQkK
r1yOHRniQQlJlG9U0RShVsohzsQKKTXwyhW360Vm/vOoaam1atOQaq0XUjB+R7GXqsS3tVOGdEdQ
D6OGVe/u0Mb/1roCo1S0O+I94A2bRs3mSoEjMd8XhgSivV4+9YpgxGyEoMBxGPbXvV/UcVWHt1Mo
68/XeVTsxhnw6W6CkAvtBksiSMB7zKzz6T8VGB5SHMlwsE27ZQ9ihpTRL4n9abe/GVL7+EUkfVL+
2vp6aya65VoQHKvnEQr0LGVYQaAw+Cdvsk/tKo8jE8oetcS6kWamksWhs/vVCYeZebn2ju2HRWSk
v0hNl8mRGU4NJwoFKKb5BgIBkUhWTpuNMtztQEoKnZpXkcZfFS7pZjzdw+AdCfeCplGmUkR48Jtf
+NQ0RO1jJ9IoYWf1VWv0oON45fPZlYy7yPw18OYx6OtZu/+wdh9liWV3Pgqu2G4pMa2iyCL25sww
2QLZsYznkKOfKgnPQPEtDjD7UnYw33Gx2d13j+htjyRx6kTKh694mzwvoJLy2BnOdh391pKFs+K5
lKGcSYLl6JBhI3Pw+n1Ll61PdP2u1TS5tyPm9pHN20/rOEFAECX/W6PrCDL1tr42t/Df6PBW7eNf
aDSmbvP6b1bwqs0Lr9WhnQvgF3T5lTUvyXeRsihM0vpAXOcTNaFd9RFucLRvynmRePgc1CnVxqHz
zS7ftFUEvIh+QssnIi087VD6z5uf66xMDXUbsGLTDJVg4lU3bFZNQt4uH1a7Yg2DraGzN6Zr0DDI
/covY9cosJvKcIg7PzlTldDfiEzt3mtMcehfMdnJgj1OphqYEGkCASreTarC4oX3be+EJiToyq68
m3c0sTaeyzsaCOJnJbcj3afFWLtxP4DhX+VPlJdv5eFlHosVUQhhrwaUlSFLig9Dmpykn5ZnRW6H
Ct7YPrOXWlBceS2UMaXd2QBcagiqQrq79ULquxEscGum0X2BAIRC3PjtW8K/H5zDLyhcYuYq0/VF
jDnXaPFeueBg60Xv/yVFxBfyAxJu9AJL/8D+7QgLKrj2qYXnEfJMMugHIns55ctYN2ffU41FE1+B
zxNqpDWG5XXbCliwCBFA1iqqbbfBy+Uf4WzcjDakbclath9nJro2w80xe4OFOoblr6LUlPd1p2sN
sBak/XDOjlFjjCDKZ16slIWg7R6mk9lRI7/gkywRCQ7Ng5VyXoTu9qcrPj3Y+xtGiJ3kR7Cnl50P
2lysi/g6r0keABM6/qhXEYl1hKuUkxaDYDF6r2nA/2sAk+3vYD8orFBNQ+93sXL9nWkN5BHTGJqp
D174ErW+3Ik8IKsUATx2GsRpvyB6GW5s3Ywaik/QbHXhyqYlUtjb7xOkzScuLWaGOEiA9t6/h/Vk
5fjgg7LlUqnx2MAP7/6hGwgm23zQ+BDGWtu6xtSMwp58F4GT+F/u0XPjdrG+KTkaA6ZSHdEhzSEW
PQlWHEZ4vwoaVBkCqbyGmWKAqkIkSe2bqM2m310SSiO8f4cKb2eC6N5msBAOLzrsVYSB3h35eeVd
dHPsZlSR+AghOr7pSdhsKYV/j902uQ5sVq899DwSjCwupfzLWJa9qynCUSBJknqqBKULLJjAkikN
XxHom2U8IzSjkGQ0uBRBUZcrqFwAzb5fBPdhtPbEvPjbHNM15nUarcgZHmyw72hrnO0TSYUp7oDU
TCAVJ69uu1UQLHJX+GqHx9XFKX1K8VCSNjMCNXH0yc483rQxDu9Sv6dt/pF5vqVHGlwYZM+pBlvU
I7TMh42JSfIseloi4c1JJ1/Z3ojb3lDt9q95+qvcmdYAGE/CI3qh0PdBygBk7Y35Ip5lLnsBhCh9
QjB0yg7bBEid7YzGxbSZYdwxF+NCBUT6+/KFpJYBJwopeNiuugEVNMFm11Aj0HIOb3kF0QPTHEmM
B9emqEDaPR2XavkmlCUzHXQC3LnK8CumxeUJmlxMO/0PDDOHDt7WlJr4Xs4AFoYAUobloMLuQk2I
sI9jzjH//YM2HNNzeT1yChSaBTeAI3vhVGdNZg0zSAQzhLte9DUi7C4wwH8FGvkPh8Y1tkxx1pN2
BG4VwTPK6dgE9FAgP+9Q0aNdTk4tMbhXRLlHqNNfQO608jqTHUsjpeovV5EqTQluvzRwHq8Pk88T
wutwbqnBcq/f3y6pBT6tlvP4xuwGMmkjCTxhXQMRxooxd3Ccexgu+9ehlzs68QBw0BfRzwPKSpA6
LfWLitbYodwedhF/GvDduuGtcjz+datD/sBAuGD3sLYKmHcfxlOp8KV1gKszJubIuAzqIGO8KmpX
mGRDM3ORZoVXoLXAFHNetWWB/AlRhXFk+JSaFZtmTUjUYNbcnHWiSpDxHS9IvPho0GDr26w1Ng96
o4gdMNdxKqjVyquXg8oHozt5ljnh9vJAVQi9R5Y2/bBfasvWZRGDt+/hZJr4ID377OJaaGy9kceS
wwP/qFp9+jtG17n3J3ILe1qoDvG0XxhrSFLBCdmOwT0zgtDXR/fZ2GaK0rtqsvcMNi7EonixD/aw
hRKRJn8V84FK1tVmCqJdmWfBy2UuKWcYVyYzIQg51u0eIE0DZR14FutCDlmToWgrdoQkBsxnXbCu
QyZdauXaTYSDOmEbHvWDZPpo9jn72f9i30IBFz1ssKWa12h2ezJGTSR6FiA+Weh61l3vRg6G38xN
UPmVapNP8J62nwyMpfDdZtAPxTmG3B3NBkzi3kP6pUPHEGYaw0t+edRioVFNxTcKW7syKXLbYSFO
+XRoZAtoBBA3C8mIidAH2UNGaFzqecJ1vkGEQUcSVfJs7iSjDNCZUJmrj48xdkjKqygXx47bQz+G
r7sJP7qrriRiR1FcvfTZBZfnKFFCn6C+AAjM8ceSbQPGFk5cNnOZEfSLcWnl7hXtOB0nKsxveiQY
TwueHTsFHcPUp3KSvRYAiqps0BXLCvucKUUQGxK10cwpH3S9BUoZPhyhIf0GcO9vfHLYUFmy2Eil
kQSw06EnF/Xd9V1tGTDo9AXviqG3dETiTykDLyW0qVKNUWuc0wPv2NlfIVqY4RqwsL80rEl9UgKt
vjd5Oc7//VUgnOyGxvGFXwOjOetRHBcVHFlW+L1qXQ+MYcRrYQzBxZDW8uZPCJR5KTF8G0fAMv+f
C7xhbiuBOhy+kMZKSdXjuSV28HpNTTXn80s8Bx4TLg4YVNZvJXaB5fJdleokiZpw74Z30r9PV/ey
a43Nzml9gso/xGKBEpMeeYDcoJl8/IYTKU7dup2sseG+VnquDlbxZri0yoWA4fjk892guK+0g6bT
Gxe9wKHhbw2cvBOYDkeguyWYTjusu+lGiqD1UCD4sku+WeOv9N4okkO/UvAm2PZJWobBfcT7aAXS
yCpiMF0ib1c/g5t7rM5f7cKMzLosJDldOihARAMfWyUJSAOIDI55xwR28SIfBD5a4XwaBOuOh2iE
7t2uAmwnd2EXt0yE1Hy5CiSOmOItZtkQsLmeOGMtEHn5sPLDkk8fvbJlleF6fsbe08yTWVgmPPHm
5xuFRTSZwRabBLKrBL/B/iVb3ShyHKK8EvCLxe0AMFFHKEOCykSjlrxpAE9v3pXGL/Jwq7JiyAFq
+4ZzNpjSY/1toHq3aWcSm72jKFE5Ayk5wM5qmC/mmFEPvQoD+qf/G1ZmiERccq3aHpUn3PGrLCdz
f87+7a6rPVvmKkwu2Xlz9IA2lbMhUiEfmoZGKiXpdoeZ/K/J2A0nBVbmxh/WXPLyYT7VWPhYCpx7
mYV8Fbh3CLQ5fa6cGqKWEPICx8klaUMgORz88mCQRQoIaWyBEYC5dSBjF2+J4pMQkI77sCuGGC4k
eqwd+plhWGlJGX4SKpRziijX5AYO4g4J1Zdyb0auq3zSdRi38RW4qpwgSi2Qz4eavBP2+N/5p2GP
/fN6wTJOznjEyWMy2eqO4QaxDeUJr5O+RSFvFwpRjHxzGvg2qHzzeNQLvinY8UKKOAwpFRl4OdC/
Rv2zHPR7q8O24wVDMcV6fRoDAoaY2jZku6SPlS4LPGrlwU69ZMgIfeJpVDTQJ4hpNaxTTcnDqHWS
i2f8pu9mPGGnghaDDVJWrTTRcVyO7t3Yk7+GqAAv4BkBtbcslzbfttdO/bGy33Bd6NNItrY5hEEL
wgKTVi/OZW0yi02jkEkFH7ZxQMVP3OR2tfFsEoToilwhILPMn/XFRH7uhe3ZVcsRG82Z1eDSrA2n
810MwvYXYbJlPRJqOD1gevGonI3/1mjOPL2h7HQad5PuAOMTIEU9kGJQYmAIGaBd+J9lO7wsUitl
4vXZmTbODZDz8Y1aYboQwaEiIW4TnoMhX9uJc2GeTNQ4RC9+lQhVP9mXpqMxqcyoauk/elrnTH86
HtJSWMf6geergY4N/TG7o9Z14kwWWr8MIBKIhzY9Kj0kh2KO/eCbFy2ktMPCiHHv7CsRiOyrZNsP
2NuJJeduC1iLXKGUTP/yuPxCiaA17yMEhfC/lhp5VMppPaMS5cSbG9AAiBln/pqz3pysYEN6NxO1
iULJKmX1EtVpydD2+TMBL1/XqMCK8Ar0JtbI4DiqNSS9c1Yta0qFMapnQQm2tL5GHqHPK9ZGCOjO
4iZZ58+xs/TnEoaKC7xU4IpaQv9NGUXdlOBeeYpuEHbuBhkGypiyVFNfOPpGd93pL/U7suvFirTl
Tin24ojjOY2AdGHOlQK0Jzsa+b+PhulfGGTGTBZkC0RxIZnV1AmQzSa3nGnKMEVu4voSTLOM954W
kK2Nq5uZXReBbHOjedamQzNhvuMf5VaNq+a5KV5ToW8dk4RcWYOqlM8utLGcHG4j6aJsSAA2WUha
iGhKvM+DfGeikHyWrK0ZFl2bTdteBNoEK8GylyQSBAqfoCazi2QbLQ+RDB4P5sKVnkaB6qvKM+kD
yw2U7eqT2ZNLvU8uItCh7wm/19nRPAWI1DgWDr/f1Y5RqYdZRSFge3ocBlbjhTMw6GLIyflUCXHd
GRXZRLGeqHDvsJMSSnVkguP9O2EmKpJ7hko536sxlgBhMEEt9HHPds8WkUQFsr5CEOmv99ArCyPw
spICdatVAWfhy5YF2gFbvAW9cDU3fcQ4lma5vMAybCrqg91N3XL+B6JjqWVN/aynbK8GlRxAeHhc
HEYY0wj0Mp56uKcV2KKAXRBGO5HXUHXU4Y0Cek+dFzrIKwWAjUdeV/mhv+xUNIqagtzEM/tyAnOj
XsFn1z69Q0dwoorlvmTWDeMMqF8Mzf9Au7QwP+Fr4Nw4y2DWEQ/OdhsY8wFAHEy89CbcAEvMXiVJ
mLc6S7MX63NBCiOIEGQLTo9TmLYKZQSOkMBWf+gzzX9B78UHbBJNljZgn1bPdadUCmMbivozudq7
aQ8IR0lc7qDZSQd34Q1/lEofYVO9KlNUyu0PF0GQH0bC+GPj3CEPv3sXAZ2NUpm9OnBOajql6ilB
mH5GLLzFPkQeIVceqwH0PN/IFKBiawNpWPY63spnOezRSfE7/YJzwSeH879jFrXnLCdTVQzbkuCY
uypFzxM2ycLmtsnoV1K2i5VcE9Yp0TjBXy2tZbxHYQQ9mlyQ0gVfswyQvt/d8+A0K9NEX7+lJwxz
rdP3wQwbQqxu+4oh3wHf8CKUjVjDGohLzRJ4GI5VB3IyoGRF9aTlG2qo7W46V8tssvngOEl8/5he
lGsBT+NmWCZ+9QJfsHBJc5Nwwi4oe/gcxixYh/xdN7vFfK8HVmxc1Mkkub0yDC7Vn7xop76bH/WC
YuI/6cYQklQ2/c58M/y8Guim5sruO0EvPevk8jayTxDA0upVVmFQI+0PT3lyzZ/I49xeZ20WIPWi
APR+QvwVdSHRrfI7Er4v9cT4zB/yIQGmOKh2SM+ueoyArQKq7DXcsyBwQ1Or0pKs9ToCB6Oz5dbD
tw4Jze1x6Phi4OtTg/GZxyXKtbQOKeNY61CHgsI4Wgh4BFRMz20pww+UT8CbfbOW/s9Bzf9fDCCE
wEI0USwMtfcgSuXoBfi0CA5jg6c8OQmmkXhMZ05yI9hUGgwwH1leSMa7GbzxhQEworGkTee/Wk2I
loUxRJX2daJVAnD3YQf4YOfWYXf7Qgl2wDOJ9mRe1jtV4tyEL820eVnFSY8bd78wamSySClEaMJF
KHWe7favHJMgH9o7Alb306crCJY41vKUM14jpe5DtavCE+zcNui50gS/ttqckSO2H2GXsjUYwV1+
SrjON/DUn/904DrvhFs2vZ4jvy33c3IYMqsCnFo7PKkhethe9Bltw1DVsoHkNRsNBPOR3idAODJj
bGaMe6prJGcbQ2LQzV1j7/SX9NrWg7gKPXb7yoq9R13EJFtuu7yU4gW/8/8t21RcmUmnoeZ+YPmX
Y8ffzwYFmtr7TCn8k9idfyWo8mNnFx/duOuSTU2CmgSnJ/ss1J+nQYrDH0u4Cuy0sFS9Xrw+zJRy
tQB9yGX/9tiRwmqt0VjjM6hYzqjBzQ82r4Ne5LAvZd7bgybO+5G3zkbEIEemleaqKUeqAwTkf5aL
BLxJDsmX0x8Vsc06bwFs7IaZO+MSy5mz4U24PY8ojxf/6rlTOdDpNdd7v3u8iu8E8h17jD2mUcwR
0dnTjyrTEF0OaIzQI00GNe/WHim51rsM5ArtqcqQyo7XSgffHDbGQYoEcGW522jdaE8zh75wS9PA
+PWGv0FZBhTafscapSHrWZBbd4UnVn0PQc1lfYb3d8E1u7elRr2Mbyf0Loe6yI4oB1yHNToBPrw7
2Z62octBN3Bbnhm3dlu30KHI2dHxoWxE4pD9H4ZDz89kffFgf9lFgQa/GnzWGn22izofRU2czKf3
OFeqUqdxtbBiTEyXTs8ZECnXOPbjrpwlPlm4A1y3jMAutD8hW4y1JJSOPaKcL72+iq64myVbYq8j
mwCCBzImzcu7YPaS/dFkqUBlH1m8Eba1qqZ4XJSkspU+7gnNGGGDcU3h3QK7k7hGVK1lMiAmi5TW
lxwWw815rORXKIGbWxeaxWvXlm9XYqmXFd5L5yxjUB4d11BjE5xGe3DgZw7GYhj562pCrswxMTUx
7x4ZECxOJ/caCVWiwgaSnhT8hTeKXPoomRdiLmzICUj+iqBRT6ZbCnDqp3JawQlUExIIAw8vXcQd
q78KxTj/D8sMzLYD031FnQddOmWY461Tf2hF7y8GVwODaMlw8+cFbsJiXh54bAXXZC0mp39UAdQk
m1A9KxBYaRm0oZ3v3V4wzf5RzK7VBrBTnvRXthRkjqyWjkxOGbWjoXBY1An/40hMhnf+mXqwW8rN
sCwoq3yYEP8oTUDICY7lbvJpcl5LfVt1/zcYIiew3qJKpersor4wedAUtUNu/LalRGHSo5BT44Vw
ICu94s0HBFHHLv1vrRvVo+uoBcf4+kbTDRH6+C51FH7QESYRecJ9fzUsUIZNIsg+S49o6+cTnTp/
Ri6MJ2kBfVfWoe5uamVSzZF7OOxOeMJNGyOzsGocKNOjnnWgCxC5Zwj5kPN5w6RG7u8GZKyq4Wq0
NXJIgNAdpw49Y2MFH4gheI242XdMEPkbWxom5Sx8HyiRZQnOCVW55F/QOXVFzmpZivMFZcKhH1GZ
t6V3Tkrm/0kX36liHl3TYTur6QVQO9OL6NXCOnmPzDxA7wMqzguEAiwSKX/otrJp1QYzZlmv7hC7
631Bo+bWa6CnDRw5usVWbq3kwwXNBwuFpfj3OOf/VTc3U2REUy7B8aCrkR/IPLqQNw6sU5hkAFY6
Ent6eoXTJ+7qRLZVGuI1MutthWDyaedjnMtK6RL/jJuhNtgGDvbNiDxCqHrZ2NDyKHYgfL44q+Rt
HLR7nfeCuf0p9ZnzMMhN0BqZ93QnyiEIqS3ObzYIfPm0ocoI669APY4KsmeYDMmsP+IPFG6GziXV
6Bf7sEuJDRKlKtpYQTZ6Z16YktZrygw9v6XqN9rUZc1FQoNLse/d4FuiLQVV6AE8zPGOFC9+TYyf
B7J4y6AOV9KoPRr1zAsSB2IeWREaKWPytabivjtuBEvl6imSXYmMskJFAPLEFPZwUkmsXDBDMOE7
S5fRKGYB9d7ZUG3lAogQKql5ow9ZPBWEib+v3/nkoOG4ihMg1rCI/LT51TplAMcRHBdzB09AUNCN
2ukfj3hOzD/MXRYxHLgxT9hk6Ha4rtzCp4N9LhtXt7z5Z7hnCj/JGMQtLGLU6sDyxnwIcC5yEDZo
JwK3wjArf8FsQyrPZ8/RdoMBv1jW5364MRspTSkNZMFbQI6nygxY2JCCnu+nm4Ib9OoptIk3q6rL
cS1txsex35s8gi0BtST3YtcbiTJrV1fQllgWv+dVQffxLJFw7xRX+t8T3hYnapd/g8UH2Dv1dzxH
5B7qevAy3R6PKX7Qqt/NLyfC+cxZe9UsjaaQV7VW+sojgAxcyqp992DAXGihjEo9Hn8wKqMKt3/6
TCRYNPwKLn7vxVeBXn9K7VvmYgsRHjIvipX3yWOYw1tdtNa2bzQMoxV/QAZ4mKZDh4JDYm1miBYo
2lingzXzOpfZX6zAXREbGjXO0zMnqC4kcnsaZbWBCDpHlT2aaEkVobjth6STPW4lk4j5tMINWZrq
mFWJXKgLJFhDFRHsyRokMUimiENhSQsw4jA9OCb0c+cGdCWqqbZFjPFZD0wOQUd5zaspt3GDiQP3
8LsUqxDokAhSK7ZTKCVmchKAOprwkY6Ff8wJltPFZJC0pFNz6PELBeXFMjPkgt/DCNR7Qn67rCha
3eOLb5pGgG74w5B5bdNxHI5S8ROU3En7Va69DE0S1KS0Km90NXq9gRO6Uq/nFShp+eYUY+z4fepf
E8IQvAX43r+TlPdBOczVUPaCbbG4kIkXZ7dlj5U1TjTkr0lCOf1838wVu5UVeVvz/gmVJEKwwniv
BAR8nugkHlXy3tKv7QttTPBOxjmo5DUOM1CThrPSQDWU6dZ47fBjsBVi0pquwSHWQK15OPdvtwfQ
ON/D0CLOYf1OXoHUrPc4RUANUAMr6KhFspPehZBifLi4AmM32GRHqXbPJ3HO2E9XgNobUiG6vH7/
MjLX8S03PPlw3/mD1W/KzcZPagOoIgdq5vZgDPVSs7hASei/GuoWm4s5hyVRtseVfkUMmns0PAFB
WBjLtScDmK9fbur10ece6EaWdB/Gi1VdsCQ+yoVqy3iqPB6S2ovHPqlb4v76DyGccshwampvO6NG
u0Rhot44O3kznNg84ugCbJQ7J2DRpIJr4edniIlYKnyDk74qkh+CVQ4A8lrwZ4y/2QvutvfU3kA7
2LmdIMo62GoxXM85RsEaf6XuL1yVmX4Y6niJ0xBEsvrL7pIqKwJqCGDRVGjk/0kQuADngWQ7Kd+h
DEfBFiVP+EEjerbPp7rxah+rHxp3g9dSVJGyjkaiN7pIW+bSTV/x7+yHHQDpqnnjQuLnV/tJbOwN
/VoJ1lO3GSR/AybiaG82VlkgJe21T1uaLOu9+HKHIQIQPfBbZsYA0zh1MxCOesfXiJuPGsL5WanE
lzbFjnNJyZkoIMUyCoYdsGn526kR92QbZpNsFJjnf71lIp2bK9mNevPTrKvvAFITmgXy9mTD//BA
kAfFa1BC7NPLkq2HcayIXgDAxIBwCPvaAcpbnRS5mLwhLqHdkhe/NIXRA1k2zXqJvzqyke6/iruf
0w1gAglQJ3dB56RMjsZy9rBqUR4md5MJEICk7SD1pV8O01L7dhFbMVPGIrqoB3El6lU5AxW8lUzL
0/eZLuXc6PcswEM9FRI8ZMjFDljnW9nVkB8ofpk3mPVHagB1vTJzrPDtBZZeOBROnOmUvq1bchkn
66drXh4qw1kf+GmZKaOL5cVZiwXANn9F5UBFK5qeUao3US4K7WwGiu+8xFPT+cT8syouwnxDLCUQ
rGWO7sq1hrUg9m6AC/uOetTkZFIcwoRNjSAtKC9uMd2inLCysE1FQxLO5GmNAAEcJF6g65KPSX6K
E6xDqEWeL8q8clBmbmfwlVuuqtJi/qHR1SBYcBnmSMc94Hun+7Dnl6L+0e0DXoD6mH+X2nB340eV
JY9g+UlXolgol5+ebiC8Uc8noW4bjR6GmiZDy3FbV1Noef7IkqDP/o6vZflXlNDQ6GMU8BOjFo1c
31yd1oXeANrebJIi7I56yRK9PJmJcKrHplTSA19Odd8o5QiuwfMLdetJbjEidLtOVBJyMz9/Qz2x
y2vXs/IdUlpPcY6b6ZR1v8eecRvb0WVJzGsYSmSvNKmjLw9s6sTJacEg8EEuFqRwp7H+kawQuM+U
LHXjKOQC2+6baZhV9oY9s2A+Q8Jq+N30leMk4JVCpZ2wL5QhN7A4kswp9uRAixSt+Ke3riWXYoYq
hHmZDQR18oCI9k4la7c8d6aogPnKwSBtSRbvDOgtnrZgPhE5aECktq4Kcq9sHgr1A1hLRsvCoGcx
Z7fnykMRvFQVADxJ0yhMydDMzohOwXq15IDudn1bO5OhMLEWVlD/aVIHfX3OVksaCW9go40v0wf0
fbewPnr6feN34fDfrM/IsRX4fz4FN5iHP+zTnDZ9/+hBPuf14AR7v9u3NehZpc5ZPI1M/lo0XfGK
xhU1SLWzF9WaJKle1+2sWhzPxe5bj9no/7peVXVTyv3QCR4DNOgV0AoRmi8hfMBFxzjnkVNzSBlc
9S++zzF2WMXrwXkGJZ/3rhU4gpb57maVd+GvV+F4yHQ4g9Aw6xXEGtisAzi2fOl1Nym+wphUjjxB
4eQjgubGUmskU63n7MWgnUOin+EYKKB2/njL55f9HZYFuy8qbDlsrFoMta2Ql8aiwVAZz3yJxXTX
DJtveTlUU54ceq2oQ1htrJ2DGIxsm5g3UTJvdFB7Liv4i1exP6Dggx4FidJcRXKpVAKUsl86PPFy
LDl8jwu6tHPxpR+GiGwgm8EhHH/6Bzx68GsNchfQnKFB7O5HhyxWhpSxPzvIK3CTL0sN0ntJWVzY
a+8OKU43kaeegcPDwSBOOpbIimUtgIUDMn0SpnfM09mrLW3rkKp2Vn8LXqCEQvQFm9tLGn5a/8mp
hdn1XAyd3K0MOXAotgEdZV+8SzG3OQoHXBi7BnmZRgDe12MYAorA/vQF4/7nsMAyeNmDc6XMmTAZ
09F/SU1dtwKLSVPAQi9UQZIYnHyCLL0O8OceLqQE5g+b3KGZzQRnzEqDi3Ytl2HtC7R4auzS+mbU
ou03t+Q1AM+QVD+NZA1NnqTThbPlUy+yLFwkLbAtJ4wso/1drbvs22le8bzJsL7f9s3P9gcaSLHW
Gvu6uoQ4VeL98xjmp5xzMej5pNNmtSkLoaIVcNGyOxg10asWaZCsCQXTj+rPbmVV8ZJi5BZCVRiK
MNNRUm+DHg5fRkFeBvuMEHhuhlvGCfy1K+ek3DcNgcDjtIGHd6B65yJwgYtwmrAoJzj7S2uy8foS
vrDvUVsGNw7FjEEBYLq3yat9nIJLFxlAG6pmJgy1UiHQcYNAz5Niz/TTbmy0JYHL2i7vnz/jqiuS
owPwYs6gmN0tzOaD93E+eLxvppL0bHMCoxTmmNcTZ/2OHod0XTllTROC/EjXLR1lL+llG3eMm+T/
n78dwYnwch+xcs8rPryAsGISnDTNBexoA7/Pb93SxQGt8d5fCJp92diaNKl2WeTbcvEOsaRKhkBx
nfZPzrznLbPDOFg5CZjzBoJs5D0ELa1Wheb75/woPpIMUGcjogSf7oFU+6Qdo+UD+/Jl/bUf1/qr
5OqQojZwCcEETieK4Z9Jpk9WSjx+N5jZiLVSLG8yuQdAf2LVMR+v/7oZz/R3rGqq6YmRHhFxbE9m
Ue8y8QZnoV9wxo0RgFXSDaNWGHnk9VuUfJSWEoP3ZyPPp/tzMSb7N3YN82/BaSG+tkfAv7kOb0ut
/5FZoagY5B/1oliCx/QxDHh49lZuKbmEIaNxwWNIXCcM6yUvlBLBfvmVj876fEd32U88MnGLedar
3sEU0Bm7b/nDFvZ5iCeLydjNkY8LlAJIo494bHDO8f3iyctrcLCvrvQI+s3G0f+he/ELMfoPkCHv
wDerQ4hrLSNDG/A1qD7aeiT06sadEW9n0WAhdt7+tUplw/kTxAnGsVyiM03CLrEGqnGBr7JAblQ7
kZ8JOtFyzzJ0azyisdGnkqnHxMPJhY//QdRKSLGABwtxgvhhRmVTEGjY2JQHb2AJz0VbXsr4MqCy
85AyXYBejG0CmN/h3mnASVSXFhaYbYPNBe8aI93zqxVq5gvIeSULslX3o9IaiGqqblachsVCrajm
1QgFEOONgQthAOK4stVeB1EZ2cV5PSAmi/c4lGa6skLhuIwrXiwcEiwtUR0a5P4mTh64YNW72cxW
RYGp3+tziRAKw28etHH/59/92oXtWDJWAp3pcmPfflqi5lZE2HboNuy+xqrXw6THyr0jsU6rfgrJ
Vo+OyKTodEaBXFzDYiAP501/LLRqSOpuZzXQKE9C9+n+KhLxvxmD6QF/+qKfzvbUW8uIWz5umAWq
b7Ai4dcHxHDxxJZwd+B/cC5Y9qo14kL74d3gn9G8qjJrPG9ICyHa8XZaxz2zwUP3vB5BZm/JPQ5m
j9TRTFBBDHw28qyAe+zNLyOwkN40L3l8h+bVJpu0WtkTH+ESucwGjc5+RPcGSnkfPn4GMXFRQEB0
7SFCuBT6SN9I1GxXeOWAQe2sKzXMIcCKZgRn21SrGY4a7QGyvgHbvUO6d/n8vlBOFLO5mtbvdFPz
uqg4vvpeeOcGtb/Ol7MoKedJffMhaJkO7LIE9nMtJz5VFIUJ315FvTDJeGsO1ptC8j6bqO0dnFGb
yjSDeFX4CDeslezLR1KuWO32f+8elac9GRa7l0714xAAyGIVE0aVIPNfvvVQ9uvMy/vdZODzqV+i
SkJ6xeLb4mHe74+yBQtwEqqLJ+zcWrE40nBUh8PpLSXYuFVcf8VS4xBKdBBxLoeP7asg+L2smFSz
nICZ7o2FSJRizQtNYFsdy45WW/D1zFC/0l0xge5Y3IOtFeRuY4PfQgbKT3LfqiHrSxwuzyQI+pyR
xe73btG0abezca3ESeAPiyVA0CBRMx08Ge7HWRCpX/QxGfDqMkV8cbG4EAnJhS/nIViNbWmNFlOd
zia3Pe5aJJfXQSxHwruVtf1GSU4iVcGNB4A/b3zcoal9viBL94UWjk2JAkhb0Us8smNx+cNMQcD9
cnGIDp3ywOUiLbDREtsp/CK5I1gNZtVTLHYRkvxS7m+BGpGnw8sPRtffLAHGBNZxdIOAVqaoo5Wf
tvV+onaH0Q2lq71zQ4QhtzMIaRQ/Axyiu8wr/YHNeQ3TaBIPzKYEs42bg5baps/2PTzdn98PB81l
Zd5b9eM38C+lvLZiWxkVENGklp7hKJbzZS+6beM3Ym9GOTCG6TQiz5ZKZX03QUNQQFas5C068uMy
9rHWdczmHgk/MbOWCZfs1An/1r+1R6nMY7wqNfE2BnWuQbBhv9H5UZ/m5Cl4xneN1Ju+TCuzGM2V
gYSkssi22CWVrJj+N6LTF5C6QzWbHs/OdQRBp43mvoE9VoSBkO3zX4bY/smOMBuuMW+ce/jSNzgV
zwAlzIcZf+3MyjW0oHG+Sg6lY4dLaWOU5geyHMYjr+7h8Jd9ou2hltiFbfOZ7VNYDI2bO+Cf2SHf
ng5dpSErOcgztdwWNU8ZrR7YgirAnvzXoByGgfk5tSEoDUVWDTa3c5xZ5bW4rb2i2bLBcSf7smw2
C7Rcbo0nqwfUCaShpPP5C0y1O58kd54J7t6+V/GA93O1W3qO6ZDhWTZV05AjTcYcDxfOqtE9mQVk
MomxNh4Rj9ZoD2/6nC4/U/lliXNR5DMZSCKpiFp225EUF1jRdvHCPO4mdtVYsyZTcA+mzmUEN1UE
HGnzh/nUPYSenzp1LPV6tWHD+P2I0M/JIhN6BOosIURJpm+8/17iyF0ApPWIJ2KF6p25jScFp8xx
I+coSE+P4cDnWFb8O8+YcHhVLdYu/UNlOAxfgsMk1dnFNOBtKxNAjCKe8dpUIm2dv9ZZmssdGN+4
xvRk0Yxbo8TAE5TrpsnZaYKShsksPnmjFRdknUhurYscNAD+HWfaWAcgksFvT9KR6l0Gz0eVBv7c
PwyY/ZvqxNuSqjD2KswkBsoqp+dTv7KXCWqlN8KXQ1wEB7ROZWYyxLowoIj/Yxiym4bA4io13tC3
2bptfQKKXC9wIJIHqs04es2evu2NpscpUDfKgrQdfZetlFd3qM7sbQTFJxPeDM35BXENZWi3V0Ei
c/96xFzz0JBM1mpSR+dy9ZKBGeO+29DhSUSYlxKpMZUJNCf7f2MBXksaGdG8FYADIr9ylhCIeB6N
qqUBQYkneG5NMemsX1yF8tFPBidIGQvLhofEXqEy2f3QUiXI7JqvcSNcOYWCJJcUWjur24Ho6ga1
MusKgA9JpxwuIn4kTizlHA+7JYUDh5BoibrhVXqzIpKy8km3V0RILLN+LokzC0d2ow1PpRnYv2pb
3xNwIWl2V52M3F5AbiosYMMzAPrWxhKh8Ox04uP2M0d5PjucM/6cH8cZyQSX1DPp4jbyHxvADJ0u
sOLAUEAQJJzFBdmOuEz/+ptHxWyyV+MFUh8JIXms7DKy2rynA5t+8hALSah1fT+xTRiyRYShd8py
TCi6X+Q6AzdX6623XRm2xyQ6FJCKEiXeAp94GY2B4U5izBTdyRJEPZdFrMJo7tMrYY1ZCB8455lH
WEdBIAH0Sn4TZvk4D38vX7O/4SVZm/nCkO/MWYN82ePOE97otoL9Ha0/tJqgP1WjxgPuK/pwxbXB
PyTA9ktMvetapr3NJZ5LId2XfS88CnsHNWJYdoWEmG3cvi8S78fF/jW1iHgXKrpFCPX7bY/rgp1O
HoZi5rpgDVb1NiufNYTVMVj3lhyNwuoOtFs1ZWIqyq0UySLcmGTGHhMqMUoL0I/hRztDGXaW/ba+
+pSsG6t2B/ilMKj2n8+8szre/raFWoLGhXrKZyIyWtB/rI+3TJuunl21e0eoqwEiKmXvRvY1NGGB
VxW2S0JIrxFU5aRLCjXloTsEpCz/5fWswUInCixWEUOTY8cRhyMygjsrRTbLp5yyH/SXZeKS1tRh
VjKsbOUoXYCsnPQ78q7X1GhaI8+mZasQohVWU0HfRd2ILSE1ATDGU0oUhhMO3zc1j9RVHV57zAe7
NAxHuOwecDkdg9bvrrupHItKwjqpnk8YU5GLAmlhBeg00gnMPyolnNs+LxSqVVaiQRcNNoBosO21
+ZYaf9HuExTSk+wDlanw3xj1zaFie8qzZmn4mBL3VSMztFY1+4HhGT5X/JiYvCxIEO6hgw2M3jrS
1nCXg4xzMyWSpGDBsxyYxPZJXyDl2i5vFszhMD6+Q0aKACd0gP/Bvlxa+aXmlQy5Gj9Jg7RtgGqf
GxeIq33jbHw0mZrzGn9ioEnU+rihJwUvhcXpDyRLoS3SprcKqEnUVnBcXa3QuKMjdqHwMyhsXI8a
+Q7YNMrbzoHWWHX3Kw5x/pp5zTZRz3HrM8ZiBt6CaSW6jJhtMynKggel4sTIQxpkIVldyn1Rnmn9
8RbsxeVs4/HJfOvndaAd3x9K3MsGWAlvMtgemH3xfzYh4aStXiXKNSopflVdklw8KI6eOHiDAYgt
byGYWKWJ77WXe6j/eE9sHzuF0agQoQdJknsvhU+mUR1R5Alq8rAM9+0LUj6uRMWbhre343NqyyWM
Z/kN7vRPwKnBrw1XI1ljUWAkz1qTvk7j5xVh6TjVExplS5PNpD+k0WfdVpHCq7Sy1R2vw/08l4wq
fjy6bjz49agKDhwZEKfiaW+n9xviPCbteT45uwWzRzEa0W+LEfSv4hHK/uYiF+4lelh5LpwjHfyK
EllWtIWmDZJpdonXOeGzKuNlQcUN3Q5E9Vprthqv68DS9MwXeBriW38jlk6HOCdEQDoOfaEoHRIt
mpIKKWWtI0Eh1uLTbLdjuFNBr9JmqMO/xzH1xUc0M2e1NKwuuMJc0Hcyo7Ch5rfogftTR5p6ti+s
q1n+6yJ63NwmwMvvXD5wNTeUGkGNE8eLZ9PR/LcgbsaxlVnJ6zXc4SJQNX6WQl2VcukH2lTU9HyQ
1E4EmnlRgugckUKMny07O4ql72OdZuL2nvWv3L0fMfJsQhmGniJS1ImzHg+oqKyiRCNiGAlJejN1
jQkesbTB+6vItzo2BNVFH2RM3ukB0ovE7ji+25VK605AOq2ZdCkUvYbsRx/loydFIrktFVRjhGJz
CBQWXUDAiSSxblCXYLsUDWMoNe9vmFDmJ5vJmrq/j17517vG8q/4rqMxQ4a7KgBMWONFDDCf3cLE
LXDxWrWas0mKI6B5XV8BMHvaDqucGFxDkjBllTsrc1+/PvZ4P5/YsPMX3dL57EBjn54U3Qhmdocs
7jkmA58BVXHTkmjmMhgY21r9k70QCKY329uzn7MgQNNGy11m9dNPjyZTJy5iF2q/ZJxE2h3b7sAL
ArYoXXtiqJ/nbk9u7hxOcxDLt7l8taDFelPs1S7QPRvwjQTP7Rr7dzJNcoUE3AeyuLXX1CX3EaKQ
Wn3vuW2sshCoLQ41soe9rrmsixXNFvA6LRC3MQ2TN+TSwNJZxj8m7N0GEn53wgcH7jaIy7QFzuWp
HO4GLfNbzVgHVNiPWHBePOSt6cOH4yIyo1MAGnsnH2SQ1c/zyeMZjdTNB4njiXXlQ/6JxOPBdOqq
js3DsumXVZHPVJxUmYKGi1Jj8/4DcqupFWvu8BuWMi3B7Oq82hAGcJTVotGJPMVPsq84OzlcfJE/
gj0WZHKD8I5Jww/0ONuiRFHcORKfKjgzY7inBG8vwhxMJ7Q2Qft+Y8QTiZAhobbS8wBnYMXmwGGs
P6WKrB0O7+WuD+gub9FbPHYZMz0zq6SsHpBbqJVVuZQ1W/oWiMte5SRCd5YzAKzeM+05XgQRP1SL
zEVGRGUZ2y2LrLnk4mIPPqbjqT5sNIftaUsRF+RnYQMUOjBKchTeCUMepw+edjNP1zyX10XUeFIE
nYSS0HFZdteeHo5Ca6sWeT5y5AErHTQ6BICKijpB6JJu2wwuQnSEcsMhtROLg2R4z3a6lsCLLq/z
yXCHi1gPeeoOHzP1b1fskSQ8jfiUJmmKAoXgMQ5l7a9mFjsCW7Sz72CwtWcI3je3GiHhbIbfslmy
hJZgTnM0PKcnsmOK4ChTRqg/8Ik9LPrBmuNLeeQUOJRKs5ccxhzN2x92BkbGGYl4Ji7pUYTvNWdV
UFOh/bhcPNcRgxqmZ9ZRn4bQzq39XkLqfM7RcMoudALWfUiHQE+JTKdn9VrJIXasLfwnweXK6D19
OGv4LF2JX2BLYyTVX26K3zSwnMcdH0YvJ7BPmAzT8eJqtJYJK0ZK3MlPUNKIrbmOUbtiaZWlNQWB
0kDA/cTLkjaJ1sQXMBpj73LxKqm5fRXJxxkv0q+BKAuqBcTyv6LisO/UvIsY3tgNf2IVGixvE8H3
L3tVS2M7DT0cbG4XMXZVDbbo2BqQT8ovX1B0Gqeu6xZKWnWaw2XzZYc2vuA/JTDZ+uvEMlniUNUE
cS0L1+tGjtR5K1rqffiHB2JD25Fem+sslwtaOv8nPh45SFlK5rIUM0k5go+mJHGD7/DJWxDnjkpa
W8X6fxDXRuVzcRcmdTJraPDHXH0M934GN0YQuK4rAwcufJWs+aEB/p2SF82kpL6j+7V77nOiJSmB
BQ3d0IHghIMEWnTcMFJuQRqoJV/t/1bHR1LE95j1+077qbJb3ryHla/yYOAS9zlOQnxm24JMKcsN
M5uH3RG+C0HkyblQzHnlEL6K5BoPqvDmUR/XHviyDwxLG13aytlqyrQzZ+d187CsOIBFZ6dNumoq
Mm9WKDWANSXOPOLpH9okqqRT/hrn7mqCwGH9QbrBDIE2DohHJGz0j0Ox8DtMTmhFGj5Idti+gzEX
+ehGmH57DXeOwan7V128r1UszvkkfJ11A66reR2fG8Fj65aQvWzKCMYYW9iCmzWL77HUMigVVzJu
KOxBzxu+RHHmyufnTBZ+hHO29ghKMbdy+2a48CWTlDW0QpVLzAHNoQXCfpF9RjR1l/6f7Jsf7x9n
8sJM4sx1aOAMih14gQFKpSLUrzUq+2iHopees5oMDd/fPHa0o452KhX5EM9gkkG0t87UiQ12G7c9
AxAnI+GtIFTZDRPjlcUBU4sBn31quh6URN1fSHdNRbdJYF02cXzivm4FsXaJddsg57dyUKPBAAdi
CcBPOX9Q329yDF2Qs9BKWRtk1yaYAUwTdgNWMsEWJu2oPGUZyhI1uCuTdCKKCdlESHvk3EsoEfPc
OLuS8X5Dlg8XzMEGEw//VoCdhQ6eC3pcH7V1P6EVx+FJ5/GeAx2JWDTmJsrwW2BzVMBB819VC2vO
AYq6/MPgVC8HrPMCWbrEC3p2aruc8OAdgIf5u0gIoZZfaVpJB+p3ZTZMd0vrhSql/QHZJFuezlR5
iwzps3eoFVwUWzF9LD5fiKM9E/OKrYf0o16/OThWOGPNuRfqTlonGbEMj0YgaSgWZ8HOloQ1sirR
zxIAnyJMGASjvbrz8qynVd41c+1aOvupNUjwIEWsh2CQTnBLSAT8TO1RGUBr+pwQJlyAnRDRj+At
OVzdrusXYSGSPzbZzys5Uk2ZffgUvDQynVvySY51Evbyoo7qHQUIbmojsxT9Z6bkJzPYg9ebysgv
AVl7neSTsol4b4mYy5M+lLi9PNN6nie8uDi+JmKIR7xsw0r4aqsBlAS6KS+jndD3kK6U2UIWfy9O
/kaoov2SUV3kz6J2r4grj6pKwh86o8Uv80ghF0Et10Y1sF0KS9jjmc6R/ZK6mWTbiqOGBPfB/iJC
3JENjW/ZpYBYLhshZSRkanO/9og1do9xqtn4P9CHjAI3lMKc9569xdyJTLp7CPRVWGzLovIYMBtr
SGFzRSAggIGZ26rGk6ipdtkxk5ooh3TfIghC4avAgF6XTBSzcBcst2z48DWQInCXaudvNkmay5tH
s2xcwqt2D74Okq3M7OiARGX0MtOrPt9I4XBPg7z2EkPtgXPOjjBvfO5FC8MN4+QXLBNbFxWprWL9
jhNp74d1kbIvFbABljqnMh6Tk3pgOiGQUNevP7jP1VoqvaEm89lBHhO28V3t56w5zQNjhFqM/8np
wDp3CM1x7rmQqRHkRICwhur5wAXnWfkQuzgyk12yoiDaHdCkf16f/aNblM6012eiDMv7MV6hQa9R
oTpEhZOan54CXKGlN6M38HWRMfixR6OxH3W21nXdbT/2FaXUsOflNhumdWUhtBLohjaC8/KMtjhN
o543HtUajp41/xzd4xqmdxwdIebzkZVKZHzF6DV4P9sEaMNGLLZObxp7FisN9xZ1bE/0RAPcfFgr
nwmjYq6M27+q/1rdxuv5XghRj5Cbflp6V/c0X6ln6y8eV+bwe0dqgUq3b+or/dCOxGg1AEHNj0jh
Ba2IoKXRtjZCrim7c041hHv/K5u5tCZthivq5yVE9rkDUT4fS3K2NeZavye8WlojDwdF1dwjUCQ3
q/eVWAnjy+GpTaST5zk5POj0fRvNlj6FnkOABCUDspgvu9cFXtcVG1l5PYcNXfCwIbrnbsRy18Q8
A57ulmPVwy1rkVMnxr4ebzN8PDWeIjuGlwQt1P8gDccIMAUcSxOdxxj3I9v9TCjN2ERqtjfq0qtn
UcTxAV2JnnFlZyWdCK6Bt4Y23iEZvZmEmOlRxNFk6twHZYfKVS6GUypcNURWg0nJPb3ItS1gRJMZ
lcLhibRwWMVzJs+9Ww7rcQmkoNAWWOj8UJeZnMWhbfulwEByXkN4eJb0cajtLlAipgnOlRdIU+TT
MrWOAwO9tOpkrSV5wq3xG7NwDQEtsnvLAgeIRfNwo6e8E4+8m3pszEFltg+U6HAQNKLPoUtEE40A
hGMkbT4OuGEYfYRdcWs83a67Tu7QZY5lFvqzQ/CEm+FfGb44RKb0b2cXr193FhS5grF4Y94hxCZQ
VA2MX1AlGEs42za6WZhghiwxa3cKjAYm+dt+F1SF4NqHuAoqbXDbp30jy63OL23uAyMxhUJTObzn
8czHa9OWT/fQcBPIKvK78QtsL9V63Jc6Q/rdM94GkN75r+eS+nui0ShuD5lki9h/RGzpHAmj+zBj
RJTovTffg9F8toWsaIDPX+XeSq/Dkg2mmxr/EWuT7Qt/hh5YZwzEsy69DfS5KqngHqxc3TfPtmPY
Of6Jo3Ggi7usGcG+6Q7CpCuIvJVAyDEjru6kBKkAgxJuGxu4fyIi3ASlEJgYfdMPTZQlJ+v9Nv32
cXDRFXlEizVHN7q0jmELcLAcZY1yMx920NJxRM1+dd+mhqsc+o4ve22WaHuUMZtt092+eFaV6a0Y
HO07UzaU9Wb5Hya36LqniZgWWZvbIUnoLMdtQnw2hB76bIipFOOZ1UxTomd5F7J+LDVaDZJqXOlN
A2uqq5Rs8m7U/r6yvyP8zjQZ3oKYoxOyvHx6HTiwTNfwLf9qrNdtiXkJhPoSt+UZudxmXu2ktGVH
SLW7p1oU8X4vLMINnW9xBNKAVdAIfohn+aCrr4P/S8k16FkxCduCLHNXXqy6AVhL+zOrrVObCkFW
3foUHU0X8NPAk4DOngQc84n+RNJd7X0m/6fcaFSHyFo3QSg6u4UmDltAYw4YpbX0lfOPKrVMtkKa
x2Dyp8Hl9gacwGIWcoGSl5epTHO1ec2GgZD2ahRYIvIAXvNR41suvtw8oEqDsOQMHaakuWvuOPdr
hTfg4Cf0iZ/041MA/wDEFsL4HiHesbiqyV71PNf5o2h+InLrWqL7lBarDyCJdks/gNM/3QE66xY1
EzgISdiWY8ef3nEMrtOo95kZN8miusd3uNSHMwKLvXTM1JSbwzFs41M7LILQ8RpG+J8zviNplucV
P0z8mgp8RBXkHpqMFf7/5UEHhHH3jiilQA2eKKxmErjUDfHAPyi1RHXb6mSMcazcZfrCYYwOqmwO
iUsYcW5T7WZmv5YTnj66cFvZkxWa5MDqLz1O/xu23pUjWZrzdueiC0YqT4tI/Bm6FMpS1+6e1HgX
BltbzigxdKQxty5cDqu7adEE4FS/9AHwwiDtoHS2S8c5afWSVkt+KEhG+uzpNImTPvqoxljyY/xH
wqhmT3WwAmus/lNug7yi5eVdDBZhlv412mYbIQEKe0+fgylXCK6dpgKdpc4ZexQCuplvAJNS8Q8R
RXtGzkgnZy1MtFNR4j+wcvLpzdsoRt7FveYu7FeO2cM41J2j0IJwEuJQKfPzjTMRdyC9vmCEDTtt
3loxdMrv9NSwxF9SUKUZ9mcrb4cdMxi4a2HNIWVIXQbZnvEHkdE5ESqJQyK+sq1YiiowE1voqS5r
n2QiRrZBtRRKuVcom9Fa8zBcELBIX37iDOE5lA44iR8U3cc5EuC30TxOMxzxsc+kCHf6LpXn11Yj
LjldQmzhkEBlNOAyPmuIyQ22Dza2LL0UxDdg0rxpy05N5bAE2U1SliKWEsdVKPIwKtOrkYso50CR
y5VCTrfvFd97DJxOSNpI9HQNu0l4mRbM/Yo9oNPOSK7EY8iG2TYQMvU34RB7W1DFZjX7ivluyER1
md2UCkrrJMI7CRNQfEpXfCeAOzclQV1osx6GabjxOeLpR++B3ernBqMMRElTzWRnZlsLA17l56g0
u1r7L3pfkk7noc+oNvzlrWczX1nkUKPwC6M4KZinLGXDOxJJuNi3tbywmkUvDqigr+hsqBDYrlSW
PYAH18gpP+PTuKDMLQvP8Zy8snkg01SNfhP2D/VYPwNzM2ifA2N+nG4sUsNAKF2gK/tQqTOdwMye
J9icLfkAc+3lLKP2TcNAagmxoAcaH+DG13z2jQ0Y1Zv9dQ2a+sIs82qKZBjmNFB5mT3DAw699tCt
7fL+wS9pCXluOIJ0mHF0hy74ISyXgd1f3cXf/5K296MWyAdoCfvsNbjT0IaFYUaoD32UNUrCOLPr
RVV/yWsalqPKdMdqU9XB8b1SlANprn3osixhbnXDXttpvbFo8A1pPSsvg89vIn/248cv8RT5Xw57
II7qI6Q0WdISTpC+GVqHey2wDMTg6D2OHq/GbsruFQ0ZxgL9Cr9pthAKAZEeteSXS1GOiqnvzPIF
8pPsJoyGNLbBgqUzk6k+/MSX4i4H06E016zvJGmDBixyyUlfXXZs532qcfq6TcP1FGdSZ28wf7bu
a6foewdgxOWyVvUU5hiqud18FydSa+xoRiBtuQEMVL6D73hkkEga7/xUgN+WbtRRtwVV1+/O/2eP
0/Ly6SrxiWiWK2CvG56PZSX60rQGIGsst0vEWpcMdYyN8CdraRCZmt9GSClU6EDhClGJ6pMELH5a
k6dIEB1UDE71hZgtOBZK99s3xorgoMeAD+RuJbbQ8Ez8B1vv39cbW6dYbKZb3tU6GmgmTJlwg8zh
TQNQwQExfy3BkGFUnjLre2Lp2SP7vYuVhi4cPxM4AKKcrxxIalSb5aRuwT7pDcoICt7v2+ol/weX
rcrMRLj3MWamyLRImmY/YKBvC4O3dSHnJhrfF1nRmXqLRk80pAxXUeZOzZqX9zLh9dWVWTV0TNT7
kmN8wSR5SAZe1Dt0rW6ZOpfJpI3l5JZIhlwAi7Rz4zLfn1zw79CxSkm+xYzV0U846jdgrXaI9o1V
xswmS2J4xsU6BjCB9hfAnZJa3JCZLAu34S3br4DQe2MaDGQh1x4nD+b1quWd7eqUPE3NMV1n0CxH
KW5pkrBfx6C6VMYYz1ege9sJmRSLqTBtLjz5SNxac6xM79NWMzHSIbgduqZmaejFDHO04KC3GGcH
ZG7eQebP1koSIfaOTQf1fWIo48bhm3DRia3EUkg9u/HiDaUA+VOsblVV3peSdV/XGsQPiWVNcUMA
FXJq8v69/JQB0SkxH1YsFD+Xo90DYC4N2fxZK2lLPaF6QlFSlMxLDrrBStb9SvXBXmmxaz33Svbu
kZ/6KJFNPYLoxE095NVlZwfF0fqeTz+zJSD/EHnTkdx4YG431W9K0Qa0w2wGi/oaMQ6u+W3Y5ywe
WVfIEmkjimFL5H9u8Q/4kClbywY6RpPuL37yHq8a8vGRvjDXP4gGVWFOM5lD9Jo3ZX/9Rq5m+dIt
aN/+kO/qVHzzRYkMDBlkOWl/xh07QhyQM+OzPvIbpIENkEYqyDcNnntdaMl9FvZwDFgtSsvNjTwA
JWpYwlZDrO5oD9cUG0VMPF9YlO77YrHFEOtDAaSlLJqykO9JZI9djKL4msjUOx/qPdBCDpd4AVnE
ya3DEjMdtJ+T4eyyvkky0xYDUoyVvN1UPDVuK3Ro4sjOqQ55JV7qDnpxXNxU26t3Y3cZrmgLSsUi
psWRPexZRX9LKdZ6qanSPgz5eXbC74pz5I69I0+8o0Av+akycMHkMSt4pnj0G2+DXSytL3N4Qcjj
AIJ/K+k+3SsoAVMs7V3BYpEOMenTtRIJ7L1eqo3OaTypOKEdFyMmujL6yVg9UhEzJ+8NrBlkK954
9Uc1W6erMzAyPIAdGqtMXUa6XEoVAA1/r8biFzjbckYoAb3jDm2Gw7ubZfdOfAbvvftgJsuk0fVd
UGHYxA5ba1Xs7t3e+9J0rQmhiXVjHCU8C2EzHjpvp3B3TmtN9DepYJcZyrluOiC559481OOIFsVg
hLbG/4JTk3FfrpeA7TPg2EdyyHNiPciWGbvu+pW5lLOWhw9BGd2YyH17w69N5M9TfSpoA4BNCO5Q
ZBdJTevCRdOIpmswxYH5hHx3hT/aj4BQUBowGPVqWctEN33OhR0rGtteTqkJ6eX0zxQckDQHaogY
Ny3kXGrEvJT5PcgQjHk+6ikuxY+V/c4kLiuGh/hvp23KGrLmV0pLv2t8PsKhvoiGBGDMFB5Vj5oP
YOb0j0imymgITWiliKQWokCAAyxsJuOfkKaPytY+FV6VAwythwH35iPPN1TAUkYPgz7a+whi2KjE
WMabQP/8rvTZq0XQLMLNEXYNlUShgoAvwe7GF2QN3seeTWLxt6aOvS9m+WXO8DSqAc2BdTCvbsBG
kcxzXIwJLxvMR8QcEg3JSLxiEfQa475Sg78bTJh5eTxQ7d+z4FIupdRKo1X/f+PQcp3kY0hH3RXE
GbGl2FXKEEUEPcTOrQWl3tq+MsL3ow4KKdMWDeAFGbqnNcUvDAuBZ6c4cvO7tTe7bJUvGeA/sl+o
S+OAYlw+tyI+4SrHbv4N/fJidC7O97wuPvp4xsdBhI8Hk9/uOn3Onr/VE9mhYOKLGlDB7WMHiP9k
2wApSAdoLhBwNq1ikp2SntY8Ev8y2oTOFUtlPO8zsYieNzf1SSulxSdduPlJklmqso4WuwkN+f5J
w7f0CYvEwTa85CU5USoEfOKmV/Oj/Q1C+V2f63Q4bOhhQi9v4pF8Mcm873LR2d77ZAm0f42Ecn81
LeVrSC+xOOnrzN0Q5UGHSxq4PsxmqXfrhiAJwnwIvzcnDa22eZnBNXxcxRxnL9XxTxuHxwSjpusF
t0OP5z5x+WRX3zdVfBidiKldEfm6Rzv2/Nsz/hIhzNowlnUAZgAZ2svJTnTTmFd0g7xKZm85O2ln
FuMMOc4rKBGMF4RL+dyrTWet+TtErKGpSHNu4zqGaSHVo098iA0IKrq8i4D1OSftqmemSKuK5+Nx
WLURA6DhcmlHTy3HKWeY4F57GdN1GoI8bAEsCy/X/G3gIgtEpkTBhtxkUtqV7lN9VaZKjsliaskw
O3F+eGHwIeNbSXVYLu2IdZLtDCMZ/kM9SAVntdzptTsSD1yQOGMzK5U+v7eMSJ2whi8k54Gc3ngF
6OOKRZpJTgFKYCm5DKq+rTizxB2V/82SU72fEy7YVvRr1ivt9ako46cOoB4RESC2vSweHiwtbuGp
I/x/hJCoxr+BEohjdhhUunzDfAXukY7UOmiZ4biStULfOKeU21pnPUohVWII/zSOtRh6l30D4eho
xbXxVk0G/4IyALw7ARrkX6gBPku8EVpbf/6zqPAC4df7nVSv9MxEn5vFQhqcyqtd5Fu5x8e5bE0/
lIT3u/aN0ZwuIa7SvUbkFQjRvR87huKOtFP8V92tErmknknyOGyj/kukpnYTG36qAapNE2un9Av0
VcX3lLe0JsMRtJpELZ7bIfLr5dxQstCZ1Ez1TbnoumGh9D5cmAlZYQYRASWxV/6aEUOybYK8n2pv
AsuiPqY3S+oug1C5h4QtA8lsP+GsF6vT7q3caQtgpyT+zxmG9CMgLRAmwmwMkRZk/Rg6p+1KenRf
JdlGc/yixfKZ+PbV/F9e/OuURast3Gpnvd59S3ktKtDkLey6k3WpgdbZ2KfAL1HyU7ruqRvrddKY
tISxcWub7veOaTOOK6tH91JFWkO13gl6JeJMMOPGSuG3Fh5zeWcpQRKibFx15OqBPFsclABoRypo
efvIVTlKFas+XAjiDN/5zfnR0lKlS8HHTCDPab6R29qQTc/vq7zaUTjPr9cW/tAYYu8DVjNBuat1
Wjwb1p97bR1XH68ei36j8minYdLVYaK+mPl48kD7n06JKerKV364kc+Em5MkTv2BQ3TwER+wtPeC
wIIDQgq8L4e5EsOg9o1tDhwybEsruUgpqc+2YJmsIS2oUGM4DZVcX/yMOCXsunmidNB65kZ5qvV/
bC0lrGVuHLGocBFCQ9a/2KBKb/CopivOmJbyFYGJ8+yMfeWNLV/mUjfcvmNBZjnQjY3NoINXJB1m
CI6HsYwGzQBwro0B/VHesx/LWjoEBaoY9jvoM6BgjVUV6srQFCtEAtymEWzO5dDZn701C//OXBkV
wOAwAUb5OiXHrpkvg2fo9p4UvOnTt28GjFuSg1ekB4vSO7fLL5Yek4y/METVBrQhmVMwKOEwJFpO
lUNGdB5shysZHOCnWNRqZc/Z9Qt3SmSkYagOPFSpyAyWu0c4ZnDDzVBtQXAZ1PQ9MSgS6UJsFSbP
5RgNKo0Pe8OosvNn1hxILFMw8Y0fH5XYq9QhVUhk8g4sifDr6dCOjKgF1Skvtra8mxXmMtiqp1jj
b2hCGovm3Ak2t61Z74MIbKos+b0FvR3L6rqz+YuxlNDCmuONzDdzin4WunnPUT7eLbW9uf9dTarB
jmIUvs6giTj1xmOXTLT2tjcUgnTeRkQmWHLG+wbZZ+kWlaXs68SZaHmKJ8Ps/xu1ixROMV0T+5Vw
ZIka4jX/HsnKxsGV7wj53+hvCV/xWEtXZle1rzJuDRMs6qSB+Jq/oj0o8YjPwOdWLYACRisgnXnR
OWE8mcdvXlJh/0VFHRpQDrMHbGjdA6NBzsNSyjlzXHMoJyZQP89DIz9iryAUhIoKJg/R640j22Xr
SGfoYrDUVyLQbpPWWHLLGBH4mNQps/MlR8WsqRWtRGhNppBbyfg562TQvOq9AlaCMcVBPXv2OZbG
iVJM135D1attNwnnkE+x2nbUNQ0RsB61Hg/atvvsebpYGgfz0CG0F2Ol8mq9fZM6QxxANipWCrg3
mZQ0/kD4hgcECaog2XJacEuvFhrhBOkihOk/98DeCCvzQB9KTDfnNwgW3YC20swtJ9pTCPLZGkHp
XG3InPyokjetOQoon0q6ZM9UfnN7TIqJufGb066uefDhTun52sy7jJoV6ZyYnXhSt0A5yQ1K76cN
QFMKXdeohWv0rGDn2oNdIg+7p52olcsh3lqpLb+cG0sBrTgLOy4tTIROkcGQY/L7RJr30uIS2gmP
w4z/tOGZW+s/XIojcGYOsWPrUhBJiRhTV6HYKdNKMiqnb50mvA4ao3Yz9fa20ZWz3gLT9Mnl4Tfw
1FG5BZyX5vfGa3SVdMUrIurc5jkneXuEFTbYy1y6T/hiu3CYGF/bksE3JToWZkOJDg4Cf0NGdauc
16HOUSmRIDj5hpZce68ApAh9tIxuqueP2YhprDAKRLVJG3efXiGoEMYrz71iq/8wW84/QOZzcbzV
kIjbGPGQPs99ph+H6ZSBVVwwwousXWFjCQ/xwGo89Dj7P0Drd/u8Rr2JzJJZ2bgGubvmRIbULIfq
Rci3lQicd9N0Abgsc/KbM2CuDXmP5YK1/xPpY99txef+czvM0RdaKgPdZqNZYOgbcZA2FanFR1lu
NF4i/q7pp+bQaS+rp+wRnZ0QCXfS2oudTlMPeV7C8WjcqZy5KDHmDq3b0tO40uOSd6LnBhK8JcDH
exhnt5Z8pif4pJqgTS5fjez9zLBkGW2ijoVqqn6cNjFIBTT7xAnLu1QjYLR8l9b5grN/fKhAcxkp
NygG+Bxy+NHWHdcZhJs9SZwjCdfUCgcxt653M81cXgLmg4lJHV/SdWDI3bYa24KnsjJKPLaV974m
cu1EuzP5wg3bm/VzT1PFNnK94me25s6TytffPJJjYHfn7zIRAZpAzf9oYR3QLnNaTnnexjf5A5Sp
JF3QwZtDfqXgAZsx3mQI+NY+4T34qgTcAe91wMKzHpsgrWPUJKm7E3UDWiNlCXB0IlQ3HLomK0ws
L8Fs/RfkkBI1Texm/4d+v+0YwKieXw//a9VsBmhDvF6f1VBPQnugWpmV4cbLR1OP9ShlX3+1FZPH
jgQ7JqviAFUFA+di+vEfAH/TLe+sBDq+9Bx1mnytyyqhfZYQnJGnsX/LKsAX8kSR2SEc+qKypr3p
jbdf+v+seiHr2JK/QUxrVwWNTz/q+vhsKvrcVs4SABv7bAnh4lG/vHJeyuPypFs5CZL1ouQ8Ww9o
YdgPu8od5ZBH5FiCkhCtecbBSNJeByI7bzy6iUijy++p/MTY/DGHI8G4Wm99l+feal/xab5M5qI0
SpvAFwyD1/l2M83Nl6UxUrYMPCzKKyJRZmhXqOKeb8shx/cjCmMKRo3oygw2oaj0HTRKorGrBxye
z7ydm6MF0I1LzJTBrecnh0AONPR5xzFZ5hR6vkkA7gSsv0FJOUMHAWjIsvTWkkzLapZmim/a34of
7T/XeI97KnptS+XqvhWZPpeNr3j3Ag0/3hCwmvHp8OcBXxVVWeCbDfIDF84tKRqxi3mtmex6xAqn
PLpCd7OOWVdlbvfEoPYwNl8dRf4GrLAlw/mHMVuE4brIggCKKxAGWovHHAbTCkN9VfYMQKGV9grg
1+CIGL4tBXSJWI24gmGWoLPhNNyNSyxDsvi8lj4mVixFICFtg6V+tutkD0QP9RFmUf/FjTk2EWel
efDry2iOo1EUMx86qMVXcoXYHZjCWzQlJhe95ev8Nx9Tdl5qMkzfblDJRM5O7kMLYnBNM1/vbKjL
qjCLC4nx83helKgrDIRqiGXoohU6S2NVCyUFvr3WsR/+nHhTKAqLjs/jTQNIixrkhXKJ/7TigXyE
H6TfRk45wUKBFeDCXQaUwbWR/g0Ss88NzAc7f2WwSQcyN+yVt1hCfbSIqkOHtk/ClRnVmRWd7iDb
9L4EZHIj/rog07MWZUDzvinxbatCO3mj7B8nR4na81R7vSGWLFuWzEp6g7uOoDtRvMDnVxkDDWY3
QQ85IYv2BKYDD2EuqjCOk4iHS4Njo/WXv2yIvc9z2H/SFltfeNY/KzuNdr3Ij3oe3N0BsfF0Bs1b
uBvi5Fv2R+ViVhNBZIWwnNNXayutfMaw4G4TsBGvduZVgQLgmX9IeROl33N05HbgAl9Km+ERZDdN
4EbjTgt/ZvVM9MRzla/S5U7xca377ENf31CU52AZcZsPi4mnZakANePMD5VgpmIeEJGo2nyxQ+66
K/M/kBDwYt3xXLCDHt6cV3XfVylbYln98pBpcKBzViRhJeQoeoV+0fyK2KJzqfCtChRZLhPPPN1Y
ES7ayep1JVEg8LKroxy2zdNq5aSD68B/rVe6y8TA5pprCYnixVlJkP8+zT1vIDbefMhV24l8ve8Q
honNDtfacI12bUBaasJxpqm3hUj8qCFSoYsDW3GCSvc9OgPLI32B/I1kJaX8lbAxXZzvMw/sGxWP
R8GkaGoDjnuHmZiW+d48/qoA0q1mVNX2bXBKzBa2G4VI4QGW1iTvG7BDZ01GUa46pKC/SVfM43GU
XfYnpcNO052t/xQLDvHan6eeVUhiPu37zJ9vTRiz6hxh7Tyi1+IPiiVTIz/1oSTdzLwKfdUBmPQR
qHyW3YtJY7Jt6KDZrqc8FrbNxuB9EM6wPIekBnoZoJnI+ccX/H6KkpAg2qrbVKV2fiL9gpgtkEPK
DNn5xIE/zFiprIG7u8QPaxa/s5DiMITByT7naJN/cgNy27t3FAflBWAMgOPX2s+Yr1MNcE/fLQLW
S8eCJbGNjX35gZS3xKnlxunhZtcZU6/cXMm1iOzk9YW1V+/CXYlSjxxkWgQ/d8p0ZUpoL5dH1Mva
SQOv+LrQMCPMsGvwS/KJe6GmgrEFmoiTD1KaLJuDw6DaMtbL5VNOHrfVXs+/2MOfbmTp+HLhpt7c
RPB+W0o0l6EeKbyHnSJye9LDhwppcG8gV2mb+FEFzC4RAaZ/pOHmSO4RFXtRxu57b+Su7JqOsHgX
LKJ4U5NBt9u0PUHiIyW6ldZ5MojVi/hYX3663ocDcS+KhXxeI3Xqzu5VeO6CBQjiWyGM38U4l5J9
eb6zOoYlGLDAY3nfT0kYvU+dF85DtUzqkLGR0hmKLRVfoJKQdU1fATQG3xjD+ZzhlMhSlh84rhJ0
OzhgTVnKg7oWkR1pGTC0jcPB/T1yfUzMlTpzQJWG2LYwLLEu4LRyByIq1TRqbY7l+sgMV1+S+R+1
SKH1tXsEfioyAUeQlmndBw+AIwiFoUYv6QIL1IRecuwzV2sdm9Lv9QDr1u5Kka+xMS13qQMZ4N1b
TDY8Ilpy95P+WTnCvf1QWp3qTeutLWReeiWkjS6a079EIbOVajhLnE9q3wfRUMr2/apixoauRSmT
vtwIma78aMm1Q3y55BrKPVp84E2G0NXotsh5AlQe6YPehE6kEigPGc2Gr53LUSbmYqcZb14l05pp
p1xV/WYTQXbDTKzYvINS1852CG1Gy10yylrxFdMRQoZlNzCMV7spm8kwIsnpegM16XPs1RragzDs
+O0NbPTLbiP8IpAhcB6TKTXNvJ2C6rPoTXR+ZF3mAScDyYY8itwdohjxiCZFSzrehYApXtXB6eic
J2+2tir31Az4vFxhjK5i1JXGi+8YelsVMb/+rLckBBpt24ZaruzlLbaFPn49Sa6ErOEIdMnvE61k
mxvQoHhr3kV5ATgsZIjPxxT7Up8BKkClex0YSNrOXBOF8QhyK3ZmSyh6meqVZqL6FVtUXTCrXFdD
6DpRKkeiakvUUg184kwLGaSV6HzZGKyG2y9/Vx7umwg003MlXDu/M1Euz5GGuhLA2P0rHstr2EAp
vVG1IhzjzL5uAwKRyXcDfVO9xBswnR6iimsoo/8WcFYb+v8fiREYS/SZLe6Sqtj7jcxEU3h7ZB85
AZ0Dvc8HUpQpLwQVkmQRNREhCVwjDGyp+wtfK+5/5n6Mf2daONZBI3yirf6j3A3WNMUAABVK/G5v
frEFBUjwwnr+Fb8rVxcEoMGz7BGHu/AX4WZ4zOYXpaRcKZUq7KikZ/5Mi1yrAmBg0aMlxyQtXCue
JCoDP15XgQfshqnoTFYXVzAVJDUO5Hh1IAI/PgMfHgGB5ntuYDn5V/L9AG4zrDaPr4OixWUo5Gus
ZXPnLnLUOIII/EjC3kPR6XLoRIVxi35H527AJOVum2jMnVFLh3ftaIXXpy24x0oMOV8PMmdWLEu6
TyBXH/lj3ogs38HMwEyZfoucx496fKH/qgYFizOw9vQdeYqHblY+YRKR2+tv8T7AhNSs23ZT7Wa0
L3g+wZWTB2fJSi6pw4LuwP+RfIyHrc11GqqTCPjS6mvD+KlIsEmJyHLaewLmOkIiH2Ma+a53oWSM
irJPBw/k2tqxhieWE29anGZVZ5/+ujK2d1JrJB8TyJoLJpP7uj3tSa56kUahgx+Vj6tnZJsqFaEf
v6OK/MsjChCe8+s0mdeUgko2aMoqzBl+IeuN6q9/CJhs02UNmC6BJCUrlftzDwix16k67uiSqjvm
JyElEDJg1RbYu+fcbS4ConT+QiXoqYEEa9ZwTYGehg8NRXGX9babJWdds62fVAwi19TgkT+LRaYD
ozC9CmrpMxNYKiv29wV5HBAAunefTE0VcgFWAsTkhpEte1uYvF2/CznQE+gRxk5sHK1KKsiBCLyi
kWM/1C9y6ke2ky0FYPiDUFgVPMqHo38yslCrXQRNDnF1QHqfWgsvfkGvnLpvk8UaCDy6P5MKpxFx
+tV5qMXQA64IOkFpK0lZ+LY2/4rS3WtWbd04x3KfwYfPC4X+6aJqKA2myt0l4DKRLVqYM63ujTik
KyOMaM+wR+9zk1B0F38kuHYxr46/Lw/9qv90eleBUXXCvB0utfccpeV0imbO8Yfx1lNo+1Bdclq+
yE21wzTCdRiQCqKjXC9BJv2JzgIgrIj5/NZmLhCnDKSRuXMj+wDAxU9a5pu9qFV7EcCeoH0TDG6x
pvAlWUu8B0eArrCT9vAaCKiBEPJsDCnNdlfngqtSL46wPSqC/kJEbvSCJcDgBCqI0em9kQVu+Om1
WyL1/5qccGrq9uCfHxs+DBTvPr4tOj7WeeVlNB8kuaGl3nCdIuy77l+QWQwA/D2Dc4ChsV5X3UX6
f94ZD+e15cPdxFHdWyumlL4dBV+5V7/s4AhwAZtNX7Ler/dCmOfqzwRjdDZSotu1y+H8s+TkWn+r
wnDJBQ1p+06AvhBRolD4LsYmZOI/wg9h2qlx0J5PTlyu1zRsaeKeE9JjaJvzu8bZE9ndy5pmcIet
Fygq75uSXWBJrsVZuUGKoxXpwUZwN19XWF4rwiFnETi+t/BqnO6uZmSEt3f9py6GGFRAAyFxCFUF
qwAmMPTObiwK74JpJwmyHaqil8Q/8wcCTJLnWUx7ofhXr6y0Y+SoC1dkcN1jCldH5ly770i66/1w
0vWpOvi4lWSN0mu1nreJtbh+GctjJol48ad3akp2CsofM1gQLSo2oVHsm7/kCjBMLeB5+c39GHmh
UrxxAlo2jaGfGFCU3AykzyJOTSTn8CVeyMjxEHrZA6rrxSE5n4TszkO5A+hfjAYQbGy68Nt1fSJ7
7lxtfXjSjxV36v+AQAU+OeLfS4mbH7oUhs71QjdguwCaz72P9FzKqUT0uR9S+463CdsUbWKVdKuf
Q9oxzX8Df5QuhPyrhtxUnoNgPpNZOpC+9KmZSUu/qsvaxRa/Cl99ZRjKjvKnVJ9Gp8NFKu+pwrpF
XIIywmpkpD0zxeZ4EHUhYK+fz3E8q+RDuJiVh0ok0CW/dfl8aeToxd94/51gbl4Jm7nrisR7G2rz
XSv/P+GYj8SukHjaEnq8nI/Ii62LB570GoN7IpWk6h6jKCSzYYHK1VszzEhIVb9NmbpjCjGjpp8v
WhXzfxWZtiDVHZTOWK6/6gZj9O6WbF7pApywv0uJWNbP7q19C1Zl8ecUFaKdAqpA+mT2mNin25B4
Y+c5dZGZMjdYcgznb4dGOWSUgbM6tES12DAkKy/g6wNou4JR7Y3Igi7TC2rim+fExfKixGrY3T9L
QkznAoeWQTXgM1S1wwKC7SJwHzlhn840sCE1WlJAnknqJ7EVn3pBBE8AjOT3B7v0FRe/tXDzV0wx
u7LwiOKLTSbbvaMLxMXbkFV+gyzFerRvvRAxIMvSqd5BQ1JNQkdS3ODSoch5pKuMs2SHvMDQpowX
zQXHSGCqYDxKUadckGlp/a9siYlLt79uMT3wIfMQCT3yCsHHg2ZJSt1TwZu4htsUZySsX86WOCZl
BN890BIQKTYBkn2CmTixpVCNaaAUErDjwi4aSo3vi6OH5iwiT6d8y3Wgh+wQCCp4yE9Ybi7CGFyR
m0LE8aN7x/3vh2D5jB8vBS8mnWmMz+J4BY3DWvCVF5YbztbUy8ydwZD/GSCw5TqU3VeuW2q2mQFu
vm+v2EBkMguupdIKK3AxhpnRH+KdPrWkOCuQ0Jlb8yTKLAXMYw8tXBBajUChTXM9eTjXJ0Xkf94S
z8rq1ftEv3YHK1OFnH1BL098BsScApI7IlsVswStedtmr+wTr55c5VLJG2jbRxE7bOiiw2A9c2hh
HQp5UYrV5oIiuJC67z1+gub3TqVCNfiPinlVJThXnYw7Dj6xc8dcdw/4JaILu090voNCjmWO3ZzX
TWqxv5xTU9XgaTJ8ecbfgf0H+ToT0Ij9+WQOsRlWueOGonwUEmqK00NuhDGoRR0utDwlg/WqhVjV
sqfhX5eJr7hB7XopThWtyyKJeQSMjtd7t1ZisFV3mAPEfejdZ9I3/SPt09+2LptJ+6mhKnpGd0aN
NafEfpF+wUijf3snmkx0V9JqRrrJW1QTQEy81RMXykoAHLLL17U8GZTI1CJmj4Lnmy3VW69hn5EY
Ifp7K3cvqNSwbjtETeS6mXHGrr852KzGPsGNw4KAjgzlaBs9JO9mfo52WjWSJUl5Fjd5t4mu49aI
CrkKIrAxg1dj6SOBqYudg229GRZqd/S0TfyvSGsad0bcCvQSOyAxVzr44wZPaxi18texxFkKy6J+
DE0NUvG3J6vFLYBWIViKaaWGLbLt10KcUnJVL+vj9hztuaf3MoMjyKC3L6BtBhcOs6sXbdZY13hp
Fuw719eG/Q/AIlLe7eStbGRztab9DD38yG3PV/6R2Lp6CPBEtkM/3vRZRF+SPns9lh2/YD3eAqnv
oz4m1W+3hdh7OwgMBZAcuOfz7tdntfAsCCRmoO84ervNCg13SiF+p/wRdpeLcH3TyvL7V+5b4CD5
BuwY0ufyWLLZuijXSIqYF0qCNZS0LudpJ2/D9I/5AedWFt+JcTMsNhWG65tZ84xXyr+bjtJVPxQx
HUKBvFWRZfqGER9THHcu4nFeSJFfxL7G93Jp9KKTYexC4a0+dsu4/oNIMV+R7MTGiwKthoXTVk4L
dJ0z51nvFT7r/mw2ARi0AdVZVsqOTPygZXbwhmNmIXc2e4v/WD45TCVjx1QgGqSQH7HG/58qtYI0
HxC38NWE4PF+xfW4uUEkuLEKQMqO94qO9DTvFvHsGuQBRzvryYyUwSJwNFmcEUzMrpa9ij8wquFi
F3ZRS5E87SpUNzdMZwypWiKx15VfomNBvRsa1ZVLb4+qrLTqDB4ryQ3MZMdLn+uCfFylQU7/d65y
8vnMqZ5cJHjhfRP7HxFACQTlL+bUk0l6cgxQ04UDisDM12Ph5ONgG5tQbf+QfxcHvo/zziMFtjXO
EF2mRxNzWuzEJSqfZu3C9+ZyY1oJWDp8F9MMWdwBQ1/EKnjd/vnDpoIPvCapjeHTJTjy4UiztXNG
Gk6hE+go1hzb3eY9Vq/Y9HPMxTfB9Ce3ftiqT63h0K8om6bgxVwYE3cr7mKRMapDAHarsc1t8UPq
n4N+SQQoRMOQ+ZCGe3Nvo34bw6GUEaVxbos61PDGtYEoZcwOqSk5fY7IAlhuzuCcDdiXmtJNPFvY
4XLvtSaN2hA/FwRjjQwKsuBkGh5QX4a6ZtasOcAE44IcxgvSMXsjEAJwL1n7bErdnkkjAEAYwFxG
aNp6sRWBDxBKl7PK/1sQYZtdbdpRsf74pqwU88FEb4wm+J40sRkDg/DGzaA6OrEI9s1B4bJmf+JE
5O7k9mNK7yu0inU/WVAH+ecYTZjO5AJwC7I6+Xiftkq3uxSCkZ3RYPg2LonfWArt4GiXfdkL9dXO
rfI2r24cx10WTglNDjFXy2+qSL464InV8g9i66Frtz92UMbpe35WKat7UZ7P/ICbmUHTTzAZd0ni
SN+cfjFF/QvvdaIVCWUz8MuQt7DmD9KgJF09eO9N5cn/U0p8J9nv2eOx3W7/GRGxoqIdh8hzOzdL
qkr9aV2EBi1EmYKzi65q9bFgIUZjI/rGXiMAPPASo49pv1To3YHr24b6/kjlJkNQ+UP8m/vyn3Ax
O5wepG7zw5RwgF2ougftBEuWsp7Xakk4heLxeq7xTvY3x7Dsw99BZAScUIcxnzB1Q30loHiPnV7B
ZmGLSeATmcoDyRreYj9X7b6TOu9vTPBHe3x4VvavLy72N3hFoLINlshGcGpHT/ShExyDOVocoRlp
UmpfvAQO8Uu/hIV/Ml589MiMR2rOw0N8Rj1xQnN3GYFVA0DS+wfIzzfeh2iIWr1YizEyCShKByXB
+Dr5R2ZDRgH3wDRTvdsZ3jyQmtyfTeGJA7V5eLt+Rp9AF8AS3/orvrGp1J/0FXDrOfXHPPVucHBH
BvzFxvTAXAZJ8MzYeeCvvSRMs3TPafkN8pGcEp8kmVDvXxU8C+IrYBW8deGkNqm3i4SSyL9zehTH
NmSRiws9ZKdi2KITITkRNHk1lVwR+6oZVpUpt8pgkl9NbBoobtl5ffx7IjnkJ/Te6vFoXhODT2jS
4Ayf03dWejZaJi3jSpw+fPd085jZlR7rkayulrPESSMoOPaF1f6aJNKBrDFfjt33ktvfp3Cr0Gva
EkZWUPltWVGdN4YFwJqTKlAzOatSBOdF87JlOYD1C1X42DCgClEGnbopVgMI8dw+bwH+At4tAvFL
LeLBG4qxg8G10hc0EglMFlP+pHW0CL7tIVwPkXgik1nioICl2jaZHwfNMO7SpxWZTERB9F/LN4tp
8NUyZ4TciIzp+FiHYBp115BBf9t0CRr3d/yGY+M++Nk2Cy9YwHx/rIr74HKKn8t5argJPTGntDHu
/w6diqEGtJObUdED3LXSh2E/lp4/TsHhSfSTWrL3+XwdLg/65RV5w+Vo206zwJxh5J6GquNsdTJP
JOwwiamixhelqsrQrjiI+chlFLS4prqRs5uFcHV3FxsVXVugKw/7sTKb3zx9g3aXKrldUpBYH7vs
quKKORBeiigmH6CEznEhxx78GFl0s33yh1xx24v8mvuelqHiiZGAwGZwlJKihzWP4LTSt4+yyw9L
+Ia2Z0UhESSzRvYqEqC2FsUMZzhI+RzRZz8zqWbQ3k3TDTNKEuBdm86RML4t+BGQukuE+UhpnCxI
Yoz/Kg9Z21EVYKk8gwKmjWeuxhb8DNdZrr9I/EV47Ieh6pLJDiPSwnO2HkYIt25lf4pCh50zjMQL
StSd4iUM0z/sjKoGE1UaFx/dyHu0YhbguzQi7ziduOfAiX9Hz9c4QelcTdKaH/LlTbhOZEN16Ujj
+o7AI2eQ/yQq+IrB5EOMKaBjGV1dEPTnewK5YH0XhYtEB5MJAPE0OZwYaYIQnbXzfv8cuCFWLlTS
Tq/w1GCLtonv/3bZyuPzCJKgVlYC0VpPzth+5PNdR1LZOqnpDkkXDVEkYTnVnULe1w1MpOR/Pqez
Yfpv769vF8vfcdw4ytGpUFWq0tlLlePM/01/2Rz87nfOhLYh1fPtxdZxsqypTJ+sMx/3xx9sTTbo
rerddBisHxW0lJ4jOfNB5z9Q5Pk8N0BCfJDrdVmRAsM5VIbzDR0hs7DQzKL7VaPHQHNAlh9RzdOt
Kl/UG4MMl6BGjMhEqdPeLyP+qqBsIWY5rLw1fzWY70nOK1yMbsSdQlKAtKmYuB/zT5jhfYgYlP4h
/QNe/hw2WUAGv7KiC0lUTgH3DdcjsgW19lxrX8EUxGtOTWKhPYH9XY1Du81pfZz8jKfIPtYDKHn3
2fxsHwh5isbjQVJhc+auxgT6PffmMJSA3Da/TevY3y5pVEY8f1C0qNTDCwp5H7fc1z84fqpk8fpB
o2FYugNbNC0jtM2VopR6CtpeWerRu9CtebPF+676n1z3WjkE9Bg3resxjT4CXqai9vlHmMU7AbwJ
VPSLn4FYtgl8CgtPkhnbl9xNT7X2iOn4ZNCaOKUUYrBkPt5V3596cNUPXG2iIiUmY1QXQXV8dYM2
tRzo5nJHPuWv8/bMC2clsRc45l4L4Xg+qnOo/oze0eHTVN+UtHhXXxI2pe/7gFCEp4Dgn3a/vD+D
I0+aki9dcagY4fRcgkxerEpb4hGwaQDqc08nMRErUvPUdNiN+ChCHETc3U33v5Rg4hrK0F2KzfTs
VIaaP14WgdjRmm8Kb4v8XYOGFErzKUmhMvjCZBBXPZfPEInWz81zCOWVdS+2u7TzjNFfLFK3dE7x
3oLq9KoRaG04bck4nHJsQVEKDvwlSCh8f8fzYamyLkUbPfnN5zIdwZyV5CsFOaTDIwdnsZv28fe8
kBrfIYzubNiMldN8rhPb+u2kdGN35+VebjH+nipy0nk0uxBa9+yV2UHiFPouF/WtTRWILlPy8o3x
+TagmBUEPuQGpeXLakcHZAv3P+kOWHQzSrJWmszTpN2CwWP5hp0RXi1bT8RPRbB+63Pp/MsWw46D
XV7F5xe6PiM4+V3z0ZeEZhe0yNue6s1wl+rPOkBE5R+56ApUl3tXX9YGV4qqsGgzUIsPI67OA4HD
1JBDJdcuk2nTVSZ6gqq0yCi1jO0jVyUZIPnoKG08LIY2cfPDYfu4rXpzbdqLryF78mRFUhxH11z/
0T/1vvgXFJmj9hHKiBdeOCG6GKD+g+h9RxdiakDk4jb7nnH8sCMj2B7aUqC9QWCWSyyINxS5T6EJ
du9LY+NobN9pCzY0pIa+65qf+v4+5va8HeIzLnSAFFjeoLcgonl2GbxGJZX+k3X2SZud5z01JdPh
TN04PTuQjZgQDirlZjx4n1VZt0dmK0Ns5fPuq1X+z0+7OXnvsANJV9oiGiqfLksfOWz6SLA4tgaF
kNKXssOPsLrpi1zs5vWT/Oh4NShBuCwarTZLljZeDfP9bbVg8VvjiLpePDUBF1fhh/qam/5GTMoH
Cq/2Cz2qPp1nNG6DIfAE3KI+isMLWxPt2uzRqNLX5nGflvsySeauP2jH+LLl43/KrY2TO16nepG9
sUgAiMFb3SGwoHO/D/OZ7HLtAWtQ1q2ySJnbqXvAyuWoZMhglJs/jaQqnFQZt0hHX72fjIPYIaIK
L48RDXBMMbyOvKizvHvZLYVe4FdyVa0m4NG6lf+NVHlCZJqMWJlIBY8EDyFMqZlVvX+W2wNRC2wz
hLXKw6rCeRwr7zAKStFRbbM3reR5s6qZWKP9RyNykxKYpqylZVT5JrM7G/RsB+1n15CHplu45aZX
4sENGHFvogAXo7/34ai0MMetQeXhKRxZOZAtSeQRYqAmnGhD2J2YaMu6RO2nMn0CwSlcgZ6oLNDD
QsM6VnPkNHq7QjBMPpLnGEXBvMTRJntKfhDBDMxLPaJ0O9iB0arFNNAr8fld7G9AWp0xu4Ky7Tgi
yzGUDvO4X0olLEGOwnpxiqynGMfttElZOh2Npbb9Md3PW9VA+fDcHStdkpzBPOxJ/cUknGBg+civ
sksUS0guXwIq2kl9+HbX1PsP42cr6/OSjJRTg5yneBll0n67zG55Gwj4oYpQYJR2CAtVDR0IQiJD
4aytxzIJ5ih79GSDVJn2hvhzm0MGTxufKvmv/ZQdPDntIZIq/aHMK9LsPN9XKycMZ3m5sZuyTmQQ
9rJKklPALPjJD1iPfc1V5ooJVYKWUI4sYKTnXioJ2UpyEHBw8qXsGCDo+P59gN+nRbCVR1KCab9T
PiZApZyvwbSgylGCp1cgbYaSlLJ2YnKsq3/f6iAQKR/CqN3Jt6dPhoamS9JbjOnoVwoS59IdBUl1
Atp1GD4Goz1Pn8Dqmd2rMhcaI4cS02s5hxVjt+Q9Fo3MUqjJnvK7fsK2dce1ZFP6pNlVe59mutJ0
zTZK/1J6kCLNdy9XpE7bYTgNg0ByAu+9Gma/+1zmfUepjS3VTA4LZzAUOFV/UwN2DFbvxpRtugYX
FpgmrUe2cBPIb8Nul4KzLu+EmUSP4x1SKZh+SWo6p74tr3i8dnaQ+iHRYuJUO45HOp9QobWqwIt2
+iFqhI/vpL/HZjEAiP4aczf5jeymbEzuP2Eol0cDmwCVCzP7+UpLHtGxDMmFYz4k/kvNIQveoaS/
4te0h9ChR3TeM+iL0M9HDxf9MZd1q9VxaJwE7TCIO1K430pgphdl2Cqu68CJywQWrClClErHYg80
PYe8xDTH4qTwGpN+c5pj5C2U8lrdcKW9sde08++hL198+1NVfX+AppbHLQw0SsqAvrmPLNFlB8Q0
ee4mD1ymt1usYy3mBfFHi7ZDzKi+NRDZX8MjN9Hm6ApLk3duX3tWHDYEoVe9GqHG+oWqPdui0Gu5
Q2HSvfxNmuSaEAzW0qB00YxWnLdtIZJLhnigdz1muAB03eF/2cOd2r7cyexZ7k9N1EIP0OkL0BMa
YKdVPc87o1eaRaFExYt2v7p6u8ZlMVBYyqKFN57KRpmp3D8OpsEVh+4NJ7ipJ4M2sJ4tw0TYHE/O
ownJRYRQLTXSHV/QwSz2a41Gwq4QWRkL8e7Y4rgjF3FyNyiAm5fWIjngGbQO0+sZ2bPZfpf0rLvc
cGeIOT1/bKn/D1pe16vWmCtMyaxktaSY7NMep99UCOSmpnQFTybffyPP3sxkMlbuxzS3F/lbHddM
nQd1roZb5ANKM9P3p7PPc2arHDz2VZabzjSg/fEMT/hMA5PxcH/YhkBX/SPN/7vncolLIEKImuax
u96xjpPk7snUT/ozJjJIlpCQndQIf8UgJcgkPy/ClMfEpQ0n+dvNainwVe852RTiLQMVFnBPSrkl
x22ajD9coPAWwiIR/TSny75cvYi+GmD40/xtp6ETpmujtycSYlgcv7HiRrmaDJSl3Bm6ju0f/vsF
/LksedqampEfWB7jZH4CjSFx0HllbKByOTyfR2sJWdJF3X3rQS/enE7w1QCzkw5GvWUts9EDK2sr
nM4JsJKyKagLWzJ3DSADZagMKM2JtDL32F6Y6UtMKxCWB1w/P/joF4FTqPHNc0yP5VeQkFAGA4ah
6xugXhqLcT96RYt9PL0Kett5MH6P41ocxC9bNCLwyPIS2Sdoi5NVVG2iygdAzl3FJR5tukctfWh+
h4MzPl0u/RRFwL6nQ3H8DBCwSuW8wbDlu4ea9igq3rW5qpdrFVprQv+Hyc1aT1Oz3b6R2RJ3xuu7
Ml2XmxDblihJXUsBc0k6z+q8qjlfoni0MkmwzFeiYBox+/16qMVI7bQHmZTKpSrPtcEavHP+BmnC
WvZoWWwmqwhKrBNOBtjhGsRH39RZpqRhNsjjxSoABScVxd8mFihwwgzwXT4ua2DTtInKE971xc8z
/WcWdrGMJdo0bHGTMINWnvxTQ2Oec8Z4upHFFPfjNeY98G1k9+4G32omp+f/oHTTdyg9m+VbmRLT
8eyb5phBQMhoDgcmXcoIZAGXPgbrdEif1m+BDZ+qJfMjlHmpQyxcB5iva9UAPVFPANxIB2X5bIGz
8Fj3WhY/PjiqYnOKOvVRAtoGONr4cp5I7NagtgBQwTqFEOX36VTl8z+EJEwXtxsO1AO8cYlNLgcw
yVcww7isXGTUEpWTOJe64J5mDsZXPS6Fjt3Eo95J3u21cEI4Gu4rRytefI1/eS1q4l6lzNNXkAOC
YgN0aS40H+5/fJV/iBsd0ZUGFmk0Ln1Wx49W8QdD9hMA7Rl3wV05s3ZJYtuZmczjuA9+jFcm7t+R
UbESjh4GaJlcRXX3Xer4GQumzqj1i8B6Pqfw9Z9zElDz6SXG0pBnAScoYrmqUcvZ4IgkSLibPhAU
kVB4jp09d7BQl54h5bM8MLqN4LBHZHKdPv/BaR+XetlrM/PxGsgTT/03pyNqv1y1LFdAmhpLDGD4
1Qjm7SWqcrJiJtBHZKUBz3m9nwV9mE3yw9i3V/PJvd8e81RJXDtVW5V8nQFsFEDkG1hYu2JJgIXV
JiU+g3d0izI7BafiL7h+sVLOLJ8IlRDEjI+/Gorl6Vq2VtzVaGvbRK76cBYHBZjp/xPnZHrYgfgd
Bq5v2spRjI8yusTmN0voeN9RKKUYvTTErtISpdTh+iarCJfMlOG5vVNWs78bE2QJh5Y8gTiThsAS
/1cdoF+1jxrFssqcc7gCUsa6uioRhYF2ozFnQAgYbJNRmw6/wA0szDltGBdGjYfzPLVZzlkUQhXS
5BUGsfuV2vRVfD1y7/PMB01flEqUfVyKJY2KJq/YhsvrwqXQmXWy8dwMqvg55ZHl1GjscPnjqVY7
8U1jyhB0IDZgX8F6DcDLpuS+3WjVbBkZxI5L11a/NgDh7SL4gfBI5Iv0LObKExwXJK17Xb2KgVv0
HPDvoycOUUZoDm1Gk9Pk2QEKvTDanZ+iIfrel1x75qHl9xcGh/EWOdX/LGvs++GOqPmbN/r/W0hJ
Yo8ViyR1mViG0xHkYmc8zdi9yuj5FupPgnZeMEoAFqa+q4dx2xAm/58bo2iPLucQ3G73IEcSgOUw
FX5XCqnoI3w+G6amIlikToU4ulYQSl/ZIAIuPD0ZpyQBe5ZHS3cAQbus1GtgTOmBPkXJFBLzKjJF
pATZvUmAvb51AF7/SxP6XQ+p/rx/LrYXaN84Zg0ljLmrMn5tJUYF7gKazU0eeqOb/LHje35ZKvv2
kNt8uoksGvoQm+7N/kXUodpAFNTPJnL/wcam8VTzmUuU8gKNPEsXMlejdQPtmB5kw4VRtAjgRyaa
uEJVU/PV1wZbgO7nZPobntwn2iVWMJOJXZL+uS6Sif4g+EcxuQu/XkzLKmCnMXCCghyEtkL5Qp7u
3yz5umlJMQIRseFFmPizgxPBSW+3b3ck3ciVzZsTG3mswzevxFXSqfeJJ6oO+0eDS7fgY2pqqo54
fnFfm7UUg69FBWOLdQXV6SNwYj7fu+9uYNZnHPRGPSV6/bAm7osBXx6dASH0R8gmg4+yAkl3jLu0
RuUIFWqEtBxEEQ9JjXu5H+0p3FQd9krpYU85KhI7L86VabwVJiFZTXQQGUqDr8K089VPVcQi2Rg+
9cbD8Z17mE/5Pmt+kGm4u4+8F8t17LQ/l2w/Qh0ObcU4c/UQWZPrW39TgmEmAMBNKipeB2RURG1C
2p0VqcUQrQgQH31qqYHovcCE0g2higKyZ21UnTX+XV+zRU8MvrEwa1zLWyaCZyLABP8XOgvt1yq+
iFO+Jc1mUnruJ7MkO9eh9FTzcdeJFUkqw8dEJiG4lKo7zHvVfclzzeu2ozaXFDeKfPJF6RhWskpW
3D5eT7cOdKTbAKsiFHG7Xte7GFGcPCevYJC+mpMVLnMKQSnjWJXLMOIUhituEKUFGTtv1hQepvVz
dAa+AO/7wvbUd0sHARVJl23IHDtgul126UJccMH/wgVeSxUusKKaxK7VmZShJaICRNnm+mr82sf5
OUhpJACcRK6IMMmVQjjISLSwPAh5PfkS3JFaNUciyP7+3DDQ35Dd6VmIkrssT/dl1b8CghOX2xwr
yV49M2R7u3ObvxnRaO36F1kBhoi3y+MU+fXipCxnvGksJqaaixv3TqNIEx06h77jqrWLp49NU6E9
JMBVm3J/FKYdlNDbG359yHTPCnQ4YskK9HtOm6xCLF7xSszPmTYLohNEw5PHHT/U1lvG1EleV4RW
NjOp0l8d0esLTS5XiJwucvml9ZSZQvJUUeuZ3YPcWDX5j/frSt0WY5vp7Eb8M24PJ5QvX3mpxigu
HI8Jy30c1hbm+LXdBPWQcRncExqX/tD0w6VchoqdDe9zWznNUPeE6OJfMpHQUKzqptoPvc0yDABu
H3QBM5Bk6Rz/uENkv9QtFl4bDVRXwwHC65kHmgPtOf3ABZJWeMnWPYmFxJrwJ9HJxu79C8budMmV
FTY6SE4onndYd2xDll19AZxO5ekl5P3ORqNHjYtGYQ4O059SwKiYW1uAz8C/lOclt9T2zD+bIflZ
oNECsTchYb6wh/d1IWrFZYojhl3slitB17x4WBhm3fOsp52096wDSYv3U4L6p2AKCABFicE833lW
XvD/+Hed0/3eu1+Z9mtyMrvMo5jRlhOuP6+UkHKtpQtBGYY75DsHTXp77mJ+jGt8bB0OlMO7YJu0
X+UNUSkiNEIyqgrNSP5sAng5rAAW7LgTJ1Ayg8JFfqSPdnChKNnpovfkHs2Sr3X+bHbzy6VoD9kv
DW/sqg5asElndddPolQvteNlvDNSdmeut5OSyIOfc2Q8vDo4h41b5KRZXAg1h/8QqZOzlSJm1uDn
xJ+TMyhEiKQ8nyM2lNozh48II/W1on2NLkRBu95ioS40TsqkfFTObJsm2H6DH+wNa6FqaBfwXLGd
QR5UQ1ZB5P74Z0iPwjIjaRSHa4v7q7sOZPGIAG2XVbhZ65/Yes6dXSNhRW48wl8togYJqxX5TD5P
o6Dh4OCHu+prKk6rDxLBHfk/rVVMhwncizEuSha4lNqcUIidD+XSm7cg3HehXv4Akor7vVTLQF1N
NNeM3ti6UVgs0s2lfuWvSzUG11d5YH3/dLxIqX+lBqUduTT8J5P9HtCHqKwVoKrPjOQpWVTZqMoR
V9guFFpaojfOK850wA/9TCMfNq7T20MPC1zVEFCJ53vOCnDmfzwuaqqki6sRCNGG8eCuN7xyqJVP
80QOQyJywDoX76WksAIxGalRzFzfH6ht8ntsov9Y818Ic6vlAkV5Ce9YOy53r9aICsPr/E9ocLdj
RWOqy3Iq6fxhTuPtoN1tUqinmtvGhSdBduLQs+Y21K5cPZI7jTUkSmxOvBSyKsxtF+uI8pT8woGN
HRLmKil+SvKYje48lNMgSZTHXyGW/lGDiSHsCqbSwysSCX9dvu1AVafCTbbWhQLMbv2+7cvwml2t
ALMSM6HVW37HJnt0SkycMsYS7KjoiqQ+GVtbKBbRusCE1SqiwHUK7QKer27z1kU1ki2R6kX7vptW
Kg0CsrujH5UxHgMNZ+8lHUzj8WECXlta5ILULhBmsFFgCWJap7q0Ubr6LWdD7VyPXr0t82Xih68f
c40TZ5ocX5cT58i/+l7A0r637LKeJYyMrEdBJCcllVR46cfFn3BaBG0tLp3XWQ2YaxfnfpzzU35L
D2OdiKduT2rrxSiXsECNl+/jBozgkXozrU+UAhqJ2d4CJClrCHEBqRDIoaFNJtZbacgZYFt2vFcN
WBFzKErzKhnrYuueWsL6nOrgvO24ziByBAqtB49ybGcoUOB8JQXVBB44hJGNW+ItJX/CG5c/M8s1
TUdnxJeus/q9O7glUgJ7BJ1NvHYcCeo67PQXOAcFwq9aVBbwK+q0if8EkqZ3RX2YWmILqhd1U4IJ
30obWm5iACtMqkAJeFz71rL3c7gqIZtaw81c+VsCr8FGSlcBTHu9tuF1iOb7KSzyJb2HLkxHjKn2
3Kot7LTz82UANkRblwYKzyUQrtRBgsMGdI9DsxvqpDFgSn2DgG3ZK2pbB2aGXh+gsELdSIBm/etE
zZMezLyBNtQUorvrnfWJz57KLy2nxZvUSHBggTnzQgVpPT2Jx7JSWZ00VqWJoxLNHAxN38GET7KL
f1rb6iv4//347HBChm0TJXevx1IsVnh7QHKMtD4kws115EVqALnYvRjM6Obpfr7JnAEHe5kBUW5o
9nPkVlk3qUDF6Mww+FqWsJUHD4Em4rgtqlH0ImEeSYZnZLC4+ZDdKe8yVIvpq/Ky1/I/QqPnSDm4
VpgyE5Srwj8fpK38QrEvKsi8XbHGpMjUM8XJX2IR7TLGZPa0ymGV7Pbu2pnjbeieHJKzzuLYRx6w
rKR7q88kHx/r10ONCDYKkScn6TNHnP27P/C3lVumB0thPTPTblv876EoR7uezKVE0ut2wZ562x7p
SHwX6q3e9zUVevTajertblJQx6/d2zLfRcRuBXVcvIvl69JGov+FaTthSOXjIq/et3MtnI5o6Ov/
6SelIIIU/NbtnfcPdEGqB11chopXyBZqh7L62zv48rHuByGWHOAm+OL1yTLVVCM4cdjDl3pAWDPF
QhSenAZBoCMDyRswKfJjd3dqT34IkghnTMiE9cyZqDHlnyvLtHP9UM9QynFV0AU49T5pGya6WxkH
ttQXx5/LnHZ/ivU9Lo2e0f8XuBSf0rNVHykDlk0cBp4Jf0HECQjF+/n3IqLx1ReQidnQO5oh3tFS
wERWMO0NtuanlXQJk103miPX9r/8XD+ZPFeDfFQ+SiBRJr39J7YrPHgmdRG725LjI6zLo5qsrRdK
ZkA0HnKogd4MfPMXDPMA0E/c2FmTFXwjAsTrXQ6ZDuzNf5nv9nyXb9glCEqpbjDo5nPTmY0vPzRo
X0uCLJUkj+QLHt/jPRhPNECjtwb41HNq1VAeZJJEvdpNNs92iWJKFepb3/Vd6+Yf3XXdRGa3s7Gg
Qc4HGQgyWnGmm6DDJqmuDZGweUoA0sXtJjRIInnH2f39lCiKvKDfaPIpiObDjIvyr2NTpCgLpgEK
ASSSYhkjQGSGDJO1vQE66c8OoJRzFXpDmdR1blsY9okG4UAeAKzxEdk7wi2QiV+o4vL4P177o7fh
1vNynsnXNj3KuwudWSALReFwt+eCIpQX1qajG+TfnqJmNbdsAL6iMCrd0lDvQWWZNCb/jqvswqyE
LZahvyrE0MecH1iXA3n/Q6al3L9jajG9Flg8jnW7izWBU/OMWOJTB4oSZlj3Fx3waydwr7Uc3MrG
g8NuBLnJOoRNy4RB2BAnJI+0U6MFwD8XNjeIipEJGq+mGV4lx2kD7fmUfs9gFE4PTe4Z4sd9bqC3
I4L4mT+hi7tA8bXfltQjoWPKwvnp7mN9LZ4aJQsr/FTwtXThOIA0W1/pWAfRmWhCE6PZL4tOESOo
ARGhAUoTyjN1FzYkozm9IT/jRCAL4kGATsPIHG5aPdBaf6fiqHa0kT7ZgdfXt6qfuOImZWx4bKh6
WLu/DlfymVepBlDuFYYK1zsZgVba3o4I4rrPX7pe71x86SvglCffL+tdHi/tlWjxttvjJMONlqy1
ZkONUrv7dFv3C9iFICoOx55sIA/flJGmsi/ClNJNT9txxiS/YJj0ltptcXj5ZpEv6BY5pQLNZY3j
YdujfR/2jjnSZk5pfErKXyFYKdW014ceR0JvcIcdEH1IZDJnkCx6MiEDgI1BPhXCf2alGNOWG2kP
OpdnjO6gvObkCp4XC84cjzjlva/YNaP/3fEp57PjAaC8/FDkgOjWGJ5ZJvqGJ5z59dlkRQ0EuM6d
RRGb6XB9y5aedVgfdzd4HFIV70XN15hAN1L4zoAECjDbK6DXTtFKT+/LLV75kVNzrrlvNAjQP4sJ
bSX2FfUMHcFYsSg4frqcoaYWraTmquiI0tSnwJt9m9VX3HAUKTUvNPqK+ztIv3ga5KXm4m6tKAKB
uduVa8h4PQt11uWUIp4rUpVRD2VkvOGSBl/YZPgTuJYTzabEoA8E3k2abXgVL4qKKS+1N5i/lk7k
eRO/MKJwJzd01HYAGrVNi44DAEjQRKxoiXxrgGnt306A337NiX0geWUIy7i07nICGSrGw8wPIjU0
JkvvboNjiA2GOH1mgPUphzilWMnl/KPe9RqoBGKarDQwfyGu7+8pGNvZL/NWA/kJTy/sodXR+S3E
COQqXERbaGwsbarBLg78atIHRLqlmqx8hjXmBzAl9vqtoJkUEi7p9XisMDPR13BmF+Olmw0hHhFE
mMbQ2jnnmrV1IqX3qXUhI9LDo5JQN5sAlyYYqUevOO/aw82jnXhM2cLJPm96ISYugFAMN8AJeA/i
OrwHdaxMjWXcsBaL2W7KBk+/GMZX4p+Gkm0D3izxoRgZVXF7gfbEkScZOWMEm/8aaXJsL+CnSvhe
UelIraxaKT5lB/oasZ2K6KeJLk6kv+BMskuHmRKrw9XRW1WR/UNivlTmUd/+1wtpymx1qWf4uIir
AfhHeKRFDOakKRN/68pWndsTGfG+iJ11u8mD1DncJi9eIFM3PbUD2iko5WPGpapdKPK13wWWZnjt
MCtY7TBU09GAOAFfDk1NOl1jZA6GNu3zGSesZZbktVt4w6LoIJEpd6WJXzM6Qw0WbLDehpNjCSg0
3h4BJeWXaVxsmsBpXGIVYoXaet63y796Czex0uo+ZaKdBJsh/pP1iDEb7gGwq7cxF85lC7hNYzWI
aALASZ4PlM1aGLUJffGATKqQuUaTMvnZ7YJm9ofH0TMJe/DB/7w61CltRfYTWazoGHPtvBSo0NAg
ZexFWiOeVNre29BHDJv+okodJAWGmEv9QgLzg6tSYgYp4R2DG8Hk71TkrSqec4IHalNk2+Rz6dai
IX23yiF7HeL7fm5KyYHWMdFWqCG4UkbJVrPmLB2jCogsn0QZo1ODTlom8AMfe4me0OZIx7f9ymcy
qLKU/q1/RtDCB0cC1KvD/07bLLUfWL/NdBrsNnnf9YfQNFiFTUEGkJY3ECek3NWxeeXson/4Q9HQ
FT3CP+EE6K9Qn6KwK8pUTTY/BmwQjgJ2Q+Eydhhg81iI0S1Ry+ikau94749/xMSNAXmsfkNDHRCD
hmD9OqsmmE6+YNGuP85eTO/eNeYwu6jJGXL3bY+iYCcBlKYdliqggsdUM99Nik8zF4lzXjn6+V3k
9qhF5LkZek0qBsi+rMbolvZKWrtHNtBdgAr4o7yAtQGlC/uxuk/Ql8XcVxA2oZMmqDI2ipw3///c
plal3EnixH14dck53dBfkn3J5rZ3VYf+4W4nDUmhlfI7OZAgEcwAwTZYr7bWcvjgQWT7sMQmWkRx
WFuWj5iEbjZPL1xFQfRj7FffDc4zNdQK7fTT9ZfSOmnW59txpEIFP5gpsCBIGWFM6exp4z9fuP4j
BZTwPuaqSCJGXjiFFXhuvVN5Xac5hCi/cJ40ANuE0Co2RoJPojjsVNNWeWonfVHsF1H/tLp1pxpj
GUbw47+FtNIAGjFSjG2raklLPPREb7oXe5/TYZb00dFIYZ9Lk8N8nplvBV0wS1AU02aLhWk7dUna
yTguOHRxsF942q4eXOOf0bzd11g8ckC1hpcHINucOWKxjXpo2p+p2mhDGC5lbDzZm4TBrAWekVze
Fx4gRPmFY/Z0zQ39cCB6vMxDW4ql4Z0Ree7XGJcoZ9xeF+bnrMRuGWql0Z9/nSHV6V5UdHwt1H1u
Jqd0x4jKQnoitxqYBQwua4n5NT4er93vDK3Unb1Lv2OaSrIWnCVDWNu4UPfS0pEzTkyISiTRTkAN
Oisq+Z+QgDCvAKOeIlzfkeNdsGYi+53B5KvPZtGibLbnBqKOoSnmq2kiFXm1Gw0u1uGVYoyWCGhp
0g+cG1RgzkmExHLATPN1Torg55LQ30IhYztcPHbC/Vxw7biv+b0cjFlfEIsdjOHzt7PMrc+VxXm2
RSDI3GyBFYLj6St5I7Jft2FETruHfb+msbzNSkkaN8iGln+d7/DwbKWcO3f5x/cMnWfMx4ZZohn8
qYnDBTQXLabvdkoGpXE4z1TlucF1vx9skH7M/VvkqWLhBrnJdQhwBm7zJ1Yg7KU+x0tvmWF97VN7
dFRxvlMIop6TMJG9M7e/vZSyGT2tZSuCVdvM6pdOc1vHq+i9Ruvp+JZ3np9ivQotkwt+plx5SGhb
DueCx6JCC8VQ1w9T6vwbQs8ioC6ieWrHty4Ops2eYtBd+/wo6mz77MwbfRv6M6haQaGsNrjjXuCJ
WBdpoVntyUOr7oejGp67jT9z4NPpYEBMlX/1uTPZIYD10iLIu3afmLcd5hxOLuysxLv3u+MjYLr+
aEYLZ2FTVzCzPNA/g4QGvJjIpBNj4Pc/+5i5Vl8XDkAj6dGQXreHHKs9KfY+w8bDgawUC2sKDxea
JiDhbZez+cAsJVOkHilC2hvVGb0OXmvhSdD+zPZQtweS2j00U2CBqKGO+Kf7dDKoZuKqoyQazbZ/
GbJAUTUAyY53ITMVrMTfbSb9wN6p5EI68FfskZwy1RS3Ne+exnzSf1YQBnuceUhIYME0zifCFitY
7uBwuXF9dQLrgeBXw/p/NplnIH0SJnbJfG3mgLqA7kPKGrVuzWpJvw2Gq7piyqGnkE6z8IB3u7NN
DQRBDby84TIBLRPjzxfXn+5xIKVMOc0AEss9lEIjPwEtrZ4pwGpR3acXrAAfdNgRAO6Qind14FuU
bPG/C0tXRKmWPNeD3T7JhiR8YScOJpAAhjqPJNmwxKMuGsQ+Ukm4zEYKyF97bQaoYkGX2/fMh9qT
HCoUJbWBDLHIUWiEiGrK9+gkNM59s6vrxBVpblVOVErVdvbghNmCfkV08kQHst0YEMaFbAWkQ8By
cV0g6pLLJsT0uUGtRYWRnhsyZHU0WI3rmIorc9YTRtd8KehUcWhQGwDaEAsNSt7rXc+gpolPGoyX
iyMAb1eRsJ8RKDFi0sAr3XOT2zYCgpYHla4gxrQdS2ZdfAVBdSgwDjTOPO1h2vf9cwNMcZIkfl1O
bwZM6wfV5aintDpcSzfjmMarcQs9cuv9edehGFb/djb43u5dfw+lYmCT02Rw+BhW+eMRCZSbOvUn
4YzNIcLaWUIFboEZO7eJm9xh7Rr9XtK1xIvj8GUcH/MuTn4hPSjDCiY6YmVVvJeizhoI6re6TFFm
hPfkElXsaJcpTE7SWLKr85zmhw60XfSilHAT8/MyZm/1pY7X3efKAitbkpMOZsMeFiE01PiElazm
HN6pC4G/HtuhAFgq26IYj7TSKHp+w7Ya1kupH8lZiL/t6RgEubHE6WyJrNxQl7A7pbn5d/1fW3/L
NfsSQ6wv+G9UPTzFXekS1mxcROcl03dSQkaHhUW7pkWq8v0DlT3wITp+VFofAeKOdXKnJg/Bmdja
JRlw62oqDZUFdSY52AvPJA1sq5ZnbOt78E0OzCpgrSGPxZGwowhYkkMN9sTePO795/5a61q8sYoy
4zxKBBrZKLpqR+P+O9OF+HXCYZR+KWO+5GOVFs1V+/H8f8c26TxdggKGy5zXVYrqd/bb2USPc59E
kYq782gLZNTLKWNmTRtjwHuw6TnCBB1uT2F1GEBCZgAeJMLkJgAXDbnUIU+zPVz32xJvpCz5LCnt
2xGpA0XDcs5seo2IADX45u4CooomIYYzfYLTo5YWmPYLvfncK37jM000L8JCrlIh+ws6guEzZb10
rXfYgD9mACeFtY2YgSkOSX1F/MjofQfZsv99Pvq+0qso7cT2fRazbhLK0YvMqyUK0iuKxgr+Pe1g
SM7unVqwY/LUkCzRq19K5WgmN+Sukf70JNgVvPFRChFMWj+lQ+6wPnZEFQEUWugu3HeRFTsHgT2d
IzjKJDHqdwxsyjfC5DU5bq71Ch+pwv9+I0W040ct3yU0FHAxTXO3mdpNRK8nFfz86Pcv7MbdB7pe
tBu51MyOnQWi8QLS9zOUw1jh4vmTcps0w9aLhKHB5qr+JTHQ+e+xn5T6albRmEAiV9xX8qp+bVg5
j0Qb/rBtHlitu6YwQ+87tqvNVfk29tRuGEAeFXFjCDkhI5wKdEqi4/iQQKqhRETcHd3QcrJ25d95
jqc7hCAiW80Db7uJTbet3WuHD9212wkba6Q8yi87mF/uqt8AokCUktG+hthpHLCC5DbOJpT8FQO3
rh4AxQZ1QFWoIJ8Risc+AHfB9i1GHD0OkU94dmxgKBYSjou2QENcFbh4iVSo5phAqIDZMssIAeJ6
QtIksC5mJq7yzeUaoJ7ChXjYxpxGYT7345wrsjyOQuzFJ3HgDHmI/gEGSxxRSiwnsnkgp6DHpPF6
PyfbZdGtArZQVfk53VOWSheWyjOo8roLTd5ZVgHX8SkSJb1vnr5HO50n+l1Nhw4bCmkyM0znfuN1
DwYhR+y4zukMIQhj2qy1+e+ufZA/YsFVfsWoPmnU69GicnYCJTvueJD1TePnAELKtDJO1i+a+JX5
fnB8T6rWHgzJzDboYiz1dS0yrZScZC+Wdn4jlv2wSQGNznxOpm5w1xAkBhQBO3iAJ8xxECjU7gML
8ydCOp9hK61VGW7k1HQZEZQ6eeVfAZ5dfbujMkDLI6iRtuj2O3ZBWXm91MHGSTxPb2S11LW+6Gmz
ot4dmFOsOPBZdOh9StZFveQxekDOa2xBDUZ3+pF4mSf1rNsDwvTcgHbz5nyIPCEnSYgjjkFcXKnw
pc1z4fZCkhDiPEG/Tr+CLFEMevRyfyQqurcAwr5mdCZniZfun996Z851GRmfASVO5gSxl/91rvqT
lirPdDzMJFAhKDnL6asuG7332EY3D7bAF3KRPDZVYtLu4Vsjom3r76EZNpoDAL8y9KLdhCeeGzGh
JNnQpIv5gcFUZYoUoBAZpwPYkQze0BpcAy4ZiOsbSpY4jdpss0J2+AJVVV9Cia0UvhjZhk5Y3Itd
jPQ/SCZIPRd9no+BJ78jwpNOKBWWDKeMJY8KJHSy9oIz6Xf7UkyfzMNrjwqvdwnrEJkH6RukyAnP
vzPqw8STG/XMrLIAsz2sxM6z+tZpcMlNCUIYJI8AW6hB29snYWwn6fi/GF6hyye6D0E6QiUA8Jql
8YPmyH8+YX+0lwwxK0LJim1RkqY/YVeL0eDYrbzPnH5z5C2MW/jKv+1Z39hj4vHjC4KT2NG2iGMK
LnwtDIURr3/qrc72lJJG+1F7tlKgOFIRUROwdXw4HVBMPGeaFqg4UDlvoJqwtg0daZ2KWlLf02ze
2ylqR2sYVxPufVQNLJ3bOCezfTdobBO1EepRuKh5J7WuNzMK9mG9fQoPFQSDAPIhMvPT0e6pbGrj
6kwju1w3pcvQxAf7fRojXYB7G45OWG1jwEb343gtzH/Y2+M8lIBRWt6kNYVfCL+wWRozZkTuWXjq
XimRA4Q4BroDjf71UN7Q8EHidU05ep3IHM0gQGfi/13vAb8dm0tOetZO3ZzENHm1+L6XZNNI/3s6
ZsHLllA++OJBjQb7N5EhrwgHAXf8elpuxjnshD4kR8/odbQC6hSph1pFFFIcN+H68nXnfUM7DYeK
NXF2zp4Im5OQpJejt7i7nMkJkPNZ6LUNuURuZETTin94BvDdqPv3B86bnyOnCWQj3IP7Bzx+RrHp
k3ImlhlQRC8Rrq8W7Xdyg6u7rb9Rm/iEyJ0kLorfTXMY8TubycHn8eSUUUPjW1D+ITm26nz2hXA7
Ih9U53/etaJSTJfY1VvlOjvgtdZif5uCKcLx0484ZMe5e/RnPFUoBmSMHrDblTulQb1No0j07nI4
StrT3JzLpPuaqS3Z0Sdm40xA90U4knlIUHw+e/avapUXZWOhCbl1aiOoRM76zf+F8UqLPI9qsGmt
KSEynNNFtykYRS/QYrP2GTGcs0DyGq37MOYZldP8iIqDJKZ1YyG2EmOCfDNf5aLD7uxcTQ91CSYI
yfiuc8Krzl3GgECpIpSzadngNzAd0oR3FxnrGtRnNLzr/XcWKwNhtIcG5i4ej2mpfP+AMr0ikpx/
kwgwfMfjJ12CzoXBmmvXV+mM0tJeWUUV4Y5g4mobwqW7UEBHJZPbHnVo0HlwGtGbAq8NIjOySaBM
lGK4KfSOyTDXCdjILoRJ5I6wCcZvxoIBYidcar8yFEDvD03JXFqmyCZ4lFpXycqNhcH1jrtcZKV1
HBoMuKD3uH1k2xYUC6XXOpSTReUajl8TyroJCGyMNCa8NqN7zGEUJYnZTcWzezPTGvhnVhuJ0ft/
M/0p6eaNQLng7GamcLgFOrz3d5hG5AucXKJikmBwuBrweCaHGE4/a3FqT+wmTTHcF2fTJar+1Anw
Tqbj/G/s351Q9bQfcJT0IzUk3Ga8JD8xIXGGdyecCuUFPARJQ02PpTsWLGKvysCJrIHFU0WYvwaG
zdsqyRMmpUspGbtdAAV5RNb7n/4uf+bfdI7IiKdK0kmlvdTE7LiVSeW5wfCWK4gZADgwJjyge19+
XxrGM0L+CodMeLA5GEySQwryxReMpJDyOPwaHcp4Heyryuu88X3BTj3VGwRiRLWhdCY6mekveUYy
7oJ09kAkgN9R5sFa1rtVWyZu7NunH1mWaGpN+dH+wH3rULfyFOl/QL9fpZb5YkbpQFNm/Orair4N
0emZVTZ+JO0OYX5lejF/82NuLbJNHs/yJji1I2JHJnai6CZRCSm6FyH99th56UNTvb93BDW/VCpO
WFQav3MePSoz6zBUBI54u9Sx36s9HcpmiX1SS+VBicHx1DjLdIpULcj/mXwh17XvnA0dkakuYTD9
zDVkZM/1NLnEpbCEGeGXQxsETBIVD2d0xo7KCpFToS7DSGydJlP/bFTQ+NaDwgUhdPtMKOlN9nDv
hUT106OZQIWynyUIHuXvujOQom5Rv1ilWj16LS97mG+UlASYj8p64FEtcVlxDB/kSUuVbEYi2mSl
BqIQ2K7FNTn36OaXkA/R65hus7P9czowgdjXlfOZdYx1ee0CJFfiDUEFCNBVw2WDlGI88LwCVSn4
ekl8L0gbfQD4mg2eBN0CYTtQGYB6WOVcdMFlmuU7eSMjb0RBkvtfKBJN0Dlsfzyw00I5v/saVaJm
FDA0hBzjj9zhyGBGHJQ0DjJzTikyHB1sHEsySrIr/ZthFHVUpXkSGn5M8DOUwRWSc4donNzyfxru
jbG5rmM1M/ljuh7IMo4Hmy8Oc3QeL//WcxohU+OAM5yPIa1eJY5V36cdTkQyV7Qaqz6bpghrYZSm
GYBD/ARn97z1VElrZ/iMu9vDLxm3GYCJel8rA7ExDk/aSsEoOHeK8LqRcQYT6bFu/9rjjDEpEcb1
LkinECtkcJ8H4fsnvKLjDWFtHLhGlEwEVG6MotpS4o42+wKdBkGj2byNia/Flt8g8ysyHFi3FRnO
Zoylnlp8zuYTQU86guEKo/b8Q1IbWmVB58dmtno26sg1qhUSVwj/fyia/EwN/iAkDdKTg734TXXo
rdl0k6moYOet1ZYYALDdQShIWhY593vpQei5suLU2TXMYzuu32ojbASURXxGnLKr6F6vh8B9/Cui
l0qHGcbskCPhP4Yjd5yGZpjW5EWuCbxnoeJA4528rsiGLq6hobRnnZ46CTKmJrq8ogelPw9yPOaD
le9BjzMTZacUrlJktkL9RRqYkDcAaMsLRItvJ4qdGy6l5wa72IxehE3CHZALz7fNG/6NsPdoDrju
7sOaHjc4ewIQ1R59Tmc6pIepObHYQv2QfLlFI5tk//ElJ99oMUeds74CT/e6CLSXFCXqQ2kpd947
l1EsdeHYLa0ps4F5ZyX72iRV2uJ2h9tD3uJ7M2I3dV6FhtLcOovkh9mO5KljQDltYHKpHRGGxqAJ
Fdm76tG8SbBWIG5R5fFc8HVD+IbqwsAXb5YZGzgyd5mqrsrBsVXFt+5nYiGmsfDxafwrDR1rV4be
JG9SnilRI4OTKKPo8GxHgsVxAeOoQjzsQGZmrwVlDE9L7IKnvl+bC8ok1HlN5Le2VuNEXbCyqG22
NyoL7DK0fyn5UqxiZqbRg0+j7B6tH37qsRr3BHK4KTibj6nqc0qOP/zgiYfctAPl6eA5kX5xHt/k
iSYRhKbJm5gKmG/pQOkQ9sTXEYqEOTE7kMl9rqf88lDvUYDyQlM5UOsA8dXvwm5vYGoSd3EZWpPw
NUz3MYrByQeFPKMvi8gmMUJK2EN9+tdBoXT6YhZ2C0kMvL7zyH7r3egA7/NI0EpKgxuPLW28BSxi
Qi3gbpG1gzk278osEGHR5FgW2tYpSTyl2i+0O2VH63fSy3gWvEWIoC5gtNrUbdVbxUki8vpwnqc9
Ys8LMAwfx979fTmP+PM6IEuT0iKpbVZV1Lkit3vAIG36Uzw99pbUQ1P+LmQTPwM71GGBOdnRXDjG
64aZ/x42LLQ8NQzpoGzgdYXHreMBC/irYzGn7pbUkNiN8faumOExzrJjo1wr7dyy9fN9fdfpENsG
j3WilDc1fLi1nl2BlxOfYITZlZ14zq0ytkR+5+DVHd4Y2XrKPw4R8RlnrsJGaDjxCLerSsl2V/3B
bkQLY4MX4gdix+ZccebeAndD/7H+dsoW8EDB8nuVmOOMd7MpZVNj+VYDAGF+Uc5lueSdq32TigjP
0RIEI2AyU4kmP3+sRqtEP/iO1qZ+2/Mb7BbOtqT98rPxN/7PJLF3pTD42gASST4w7rasWXnNMbRS
DWOmdDP5IHhXH+6LtxjcUWJ0FqpUHGwyL1SEq3C0zjVxUipCpJIeaM3D9SLBfyEdDVqjKIbVKR/7
1etSsrPn4ylS7GMYAcR9bv5elx3s0O+thXbnwwjS37g9oyMpFDkMKi9ujBt3F/EMo7eWoOpHHaqq
dhCGftH/UfSxYBQRltXhtE/mVOA2fLnmY6nQo/QZE2VrqOp9rgaK/fQCrDXwkhFNIYrqJFvf4vum
cfnwTzREvz//m/d/xU7mBmwyr06CeQ+LDB5f5pAld9Ipr+pdcVypAii0e8t7fhXKgc7M1oNrnL4D
kwQGvh/w+q56qY7eJPDwHuetNnwfLxz2DDm3kmT1pgqMxvTcvgxp1ZuBSpLh58hetUWep9cBDatB
3sXmgiWhG4K2FQwc+TN6I30Sb5mh8O9Ohw45Uc/0l4F2p1WU7xnVukb8RqVr0WRaj/2qwilYF95P
eLjg/NxI4t27dwCOBd5bGmPnHvs3+iINSoD7ilHvuC8C4xovyQ/8aiOFdqq4+0eXDP7GZ4uBHBW+
lslZJZinJ94rz8zWSK8k7oDyi/mbW0r8VAEx/rdoCDpRfuSKRzfv4eEDIeC/J6gGI9p+H6wybGIO
sLsbkIuf2dSsoCiOP7RwfLRM0w0gwPelB3gSMStLiHMmzcDL3Q2H22Dy/7w74ZmT5oEve2/ywEkR
31aLS+/7B1XMAwpFiDto8zbwiwAci77n6YTwlikDT0w9Ahcthn33eVAo+8lr5sCdXx+X5LP2agXG
7C/Cf0Wp0OBdZQcN70SKOO5sMj86I8h9Zs4KMyHyVvjeoIGu0jT7zjDTRD0xzlFQi2X89wOoOCsA
35MAaEi+qSglqGfXIt1jy2hkWSZFcJXZ833DQM8Xzye2POo3TgrgfH9gJ8Z4+rTdfxmHFFMChnPm
YRRSbepHj3w2rrQezVIM3H48wRUfGYEVFsBCUz3bY1/9K2j9g1mOWzQZQ6lFU5NMqTf0eLd7ZhtU
C0+s7L8E2PefymUc+9esGRYHD2Wx+D4o53OwBXq9sNI/+XT2C93iMWciU9zIGpc/I29ZNFXreb9F
FeuO2WuKi2pQrUeelh1Uzh4hhneysYOSm5TLVmpqd0pJ3v12BRZo/78xkakvPjj6UBNQn4ZdtBcz
/K+eAK5E9lBfMl0nC0NvG6nk1RU+Wha8fzPh0CKXf628BEHrlVKwnOhnr2BDJtKVmCLffEe8myWx
czxedY8paLdeeAWnT1TdV87x0bNiH6z20neWoSOMYjR8dMnGdzYfFE9rAdl8IcLOX4fJkdgg3wXO
eNUaZ01+F6LT+qWFFwi8A2VTKh+Kuq1ggpJbLLY2ncCWpG8Z7FeH/MUrehrl4vIUF/gc12kDoHgE
uvAlm9oiB+mW6JmvbdI5HccOIeu9X372Ahg9YsON9ldoLaogp5fn53YAtzQ1+E0yvbNQWgzm5mQs
L4EQ8eoEMcJeWyrpG6eXJGUqSa3RadHzSvxOtVPtL6m0Q79SMXpOklsTOE5zU+Wdr8mi+AhW5AG9
WHjRBN8kA5AzT/CY0KGCXSn35Hh55ueoV/KMBQBileHL51qip7Eartp/9txbVhcXLSyqjloQ98/V
kWBg5+vbbBh8rbjTBoIzuiiSefugAjSIk4YlImfOG6e2lU/21eiItcOQYTiBCYiWru+SDAloZPdu
GgGoHntC3KQTL+48orbnB59qyjsfHb/DGUI69cNmovKMTaHQ6djmFtgAznA5mZYqFWQjSGAbCfgx
r/gr8qo24Y0AQFTA9ZBEL1ENxj1mW6MyhJgKhmZ/s/gecCOoQXidTdTPVT1Ya2PDwD+kYfVFondT
fqZ+JFuo0z+ae8MIl9gwdi4lr3i4wRO9wjtjNCgnzsUUN5gdhkPG0tQpCp0oFN+PkR79nUF6toy/
tr2B20Pupdq5bZVNSFMPtvoMPoZlxC7QVRQJvUUy5XRc05io9NIP7uPFW5ogNi9BuGJz22LgpB/T
Ky5FlsY2hDQUXvBh6G4dvnNbJnxf8qTWck5YqPYCFlDVFDgRtRujEOtrr8MSSGAJLTPRe1mrtQGN
0EqfrlqBjnGZaUxt+u2FLJmrJWRyAC339RaZrcv8n0Ztda5Ek/xWlT/xUONsuuUJP9KIEc3n6Jew
hATrkZdOPlBgVrjlighe1REq7VVG0+uHyAnChbXek14/5zIy8W7al+/9eRrRLtq+Q+UMO+Q0q1YX
cBXnyAJ8ip+l2PGAuf4Eg5nJGa9ILsNkmJUEEH44BksnsmFTBO/sZiRZnORh3ii1xReYU2Te6OQA
je4VRwQfEO9YDULsEcpxjuxouvREVxLJrQXZmyO7qKKKu3Riig+D5lfIzv0h6UMUadUQe/TALeQq
3uwlzJLFQZqnEOoj0EuF91X2oz7BPqsa06n0eXlC9NYMrfhoeo5s9qmh9h0mzyvyobfQbUb5L55s
WlYfePV8Ofliuq/RmXCnwpNquxJuLxTNDdn1VsN9o+NmmM47E/35yJ7PagLyHQWiIo1Jy8eNBxRO
8A9AOXO9gGukTycnese9vfA2P/gt8pvlEJT5IMZyFzqqE8qEK6LjN3mQPfWC8/BQzxLXUKyhCrjl
si0oVnHPkz0+a6A1rxOfQ/9rnJMCdR33AErNFwJCbnVrgMual+oIn4rob4HH9R8xCSEKQvvYl4iV
dKUwREg91DsRHBXl2qkULDEpzAKLAk2mp5vXX1vpHke1vGWSo8CTW+cacOQ0PvZpblZOMU0omExn
7+E6pOHAFIy03r9rk0bIdOH1zZrGTIBo0zk0RPsvU5bCqXec/WpIs6jTqtuWruMqXme23r/qeQuS
vi0A5x0CwyJwhLfInUFgpfTsK/i0JglN+4NTagTyAHiEL6OeiriZB999PbuK3rMEmg9aTqcpt9pO
A4ZTpIw8M0CiUJhfiWYKuSZqeQQu73fSI3++he/4UbDQzJueYnI+OxyRKIszuCAxnfcVmaZ48FCF
DX4L/lJ4nJEmC9NbNhEjtn1dVU4K5/n/vaGEWxKzakJSUv6w65dhPPEAc9zbJIzOwHL/DcbziSV0
C9iB4VsPApfsaa1PkJqw9Cm2AQFkaC1g7kKnipMSOARV7YOXwQu1XkUBDDHr8Z6FwDNDlx6S5MNn
B7B6kL2j4v20ut/xPzxsjitfugRLqN16OwAkxkioXAfuArdG0L6QCSJR1azv2gYIhIW9cC8wpuXE
Ir3JBnRHaVnhFc5AZ3r1JYSV9k+LiCZnKfp6D/RRZQf5thYGztqvH2WmVKbA0KEpbYK+QvulZu4D
QWVjttR316Wi+vu+3/yAFNC7d8TN03syDDoUNh0VNzuFWNvMF2+4bY7U90h8Z1L8ntxMQfOZ//e3
bhv1dDnWZNp1kFkQOGxCMggMWa9yLuq7XRM4+zTOH1fjSshMvdMiOZApCEAlRY6MZ8sweCzFIpdu
GafGd7E5/TwynqczCEhm8bAWp4UG7baU2Kl7oz9T29vHjauksf7F9AH1tLDAO/8GiUQEyssspFph
zjYZn47S7RKTD2nxAXaRsFgKrPgVctTbP3PwXWbJiuiNmVvRTX1xqQmhj8jhoNssJE8IiiYmo+MM
FXpmaj54PHbOi0l0phoLzVESIRIyy/PK293C1DTumkNeH/Hh21N3spxPK5eT8UOhf8nwNNe/XSAI
46a2fBNZdrm3eEI308G9VZVW1CdtbhsA2yMxMSoOyD16hYeh41byaWinKSYi4UDq9NFnuE6utfvJ
mZuHY3CBb+mcDuYj8MmEdtLZs7yfC5c1uiiZBGmgKf2PycWTtaeo15VvuHApL8ffWWiduFAp/fNx
gqGuGg6xjgWcNuhnRQn72lI4zlOjfDGocO6G3SoAp7krjxS1uQKe3fOynxK6G9F9cqp/jnPAIBzQ
PDIdOo7Yul11+uFl0/5+6O2no+tJsDNbAHY8vwvwzApckv3Lt9Kd4KpaEwjjs6/m2uTE3Tqthot+
WIaOow2NL/8Vk5Ct4agJOKRaT7cFQ6lwWK3mfVLpCDUOlN/H/C9EAbzDe/nGqhJcQlNcHDrAGHMN
IMSJtav7UyJ01lIQ4WMhFkcgR+GiOT5SgkKs4kfKOo8ePlN63NNER7YHZKIHpu7hJW0ThO4V4Igl
nVMaBFnlXFgOk6JT3PGB2hVPraaslhp1PUlTDGr6eGbaK0XazChWNRiibk0udpRLGFi8gY+t0gcK
2oe0Kav7dmINp+HWudXKRP/uwELglgr4WYJSBpt3GnrzLefW5/JQZZB6NlozVX2O0ZVEkq0fgPpJ
Q6rJB1/JfpIluoOQena3wWcMyyMX9vk9ZRf8o4T8BKwo7DoLi5j6zwPmDP52KQ56EFulKVvTar8O
A6KE8mYDPPXZaY98HYcd6hBMIAzq9nqL4aDkU0qWNgskdQiMso2inIJfGp0th5NR7I9f8csVQqLk
szMJPXv8LwDVOIx8OjteX5SJecJO6GvfQo4HQFUEqnDalKnJnxahJV+G8SUiq9UEKinwfm/GVRvA
3juUOHNwrnZm+6oD4ZDNCkT13+Ffs2s+kVmkuB/SE09wOsDuuGXXzuDgUj8oGa4ZXFQRnqU9osiv
d1yE/lcnAghqZ2A4xg34Ep1uKnSLuNeS9grbb5GzY9mhu8o70IuiQ1kQV886w0DOqV8xmbm6NznM
Uo0OJQ7uztTlmewq9TPsvOUMW86ujQbhxZ356u2u1QAW4gl2cb6N3IRqNhCrblLYGzE/K3MH1/IX
Kg4GU8eSx9ZePgcHYPOYMVmob+BY0CGrJ8AcvrZh+QMIB9nOUW3yqR+z3srOoay8duXw2N/+K6eR
7ZDrcajFk0WXY5OR5a7OaDHILhS6MpQQpuCoca7nuoxC/Qbn0Q3jG8a8Vb8x8y954gHjSSlzXQ0H
OB6eD9JjsuRsNcdG0/6IDJe+ezRrXT4L5Irim+/SaoFx0AyN2Rngsi4Ie1omz62TYp4z9WIBEU6v
xTyBYi6x74hX3jAByhIimqx+EmYjQ5Eeux5E2nMdzLYgM6gyB3irfdvrZL5SF2YwIAZU+hDUdh6w
5ffbSZb3JyUyTuxxcQf2Tww2IjkpenL5J1kot58OoJlLkIYN7Ttdsle6+RyV8ICm1OnF6PWA+s++
px3vPp/pvcoLcdwv2HO/Wox2KcXEFPvAT8PRrzw0oejTCK6fOojH+AtXEj1byEH9wCW3+6GBxlD7
NS1xTjTgLEh2QylSc61t1IRus3jmpkUEyPX8/6fDMk8iiHmSC7pq/m0cy4vWneO+3mL97DUWgmdp
yxZ/UmNYcLI0AeulHEIAUVr9iBESchXdKt4lLn5lOGdNIXJAAmL9Tcdpl/Uwgydi+VYP2HPxJpok
DfQKE1qQq70s8KmTU3GlPEaqKDcgI5quGipG/A94+JCgB8NQwMSDprD2yqJPx8xGxmb/UYp2KpqQ
7/LIP3FjCdfRJ4kauONmrnBCLjYizTeMJtZkb2Xh0IVuB1wUAKpaapeac/X5O+XQTahYaMdiikdK
IrzNN9713y6D207onuaJJezHwzW0TMNSm1ft5XH9t7W6b/wqROe4c0DTrhcKgWokuYQGcXmA0GbZ
hG5z7mDL3bX1HcMIiD1lgILEpiKqxRXD/srGfbMuV3DduiqElk2FF6+CAGwVAcJl7OK+85ZxL4Tm
txjrQ4dAtuUy4ST1wvFiPoE3cb4gITv56ofKYTnurvuIwezjYBqe/kXtHl90PEAn4A3dcqQSUl5t
h26T5VyoOkAZjFPPqPXIroz4wwLhV7WLvM3E5AAoz+R6ezBrILN6j/HazEsG/bnWBEaP948wywyo
05fKF+BJEEXld3OvkT9loTPhS5/UgVvx7IFzFmQYPOn9smJa6IHtPPo3knoYXsXUaMb4G5QMQGAy
4WmPHKWIKspUHKUK1SZvADsfrUIqSkthOSi093fQ6pylBxR6p8HyO33J1hmaBUm/t46JG0eIzyBa
nXFo/nzturdFrcsbURrVW0EfuNC5oUeB4oirU1dKGuqLMdlOPHNS+XwhBMSS98vq7YRepgWkAFEV
51g5nq0OEuxgXRCBQmfJWoKpgtEePPvTOPRZoGKrhrBx/FGTVQvd2nknHqX/VQ0JZ8ZPMdU5Vkod
bU1Eaywmyv1GS5tWGq4kLHIjsG3CyXi4/+kT3yAjKXo0B0dXCboOXKJ2TE8NEcM/AmzFVCQldQBE
41OL+oHaZ4wh/91X+LSOP5YZU8he8xZXqJmfCWz/i8YTMCmmpCnmTA7ZayV9T0GgYgoDM7GxSc0N
aqwVkH6LR9VvhHo5Nc73Mzl1LLvLYb7LNj4SKHWAPL93Ye8EPLZeQKWs9whZ1om4bA7A9jIUmqk8
p6QRmOlpagphMwdTbFHwrCQD/kFPri8e+W6DYDHXG8E/a3cpL9RYpVXJgzTluzuFs4mnU9XFCueI
mb1RuO/8E4ksdRM2+v3dYweVZIxpbrN8L0WlFWIEBNNcwYg6uV2fN9yqQqK1jBVoTGWPNyVg/nXh
ASj6iDR7dmKDKPUNUJzHeRtflHQYSRHTvrRM5gidC246eEIZP3QZVbuBq6iPa9Dgdk5guopFgiZX
WdtfaEf2VPhKsPvhp4Lbq5GL/TS+x8qVViSn4kQNwfHuHCVkP+GvLxuYiDnYVtAFbtFQzFJ2t6m8
dYGJzqvAsjpYX4PVTbd3U4HOvo2OF8rnJC4i0nNJ/NDTmjk9KmzeBImXwtsRcgzCchtm1QBxDLpB
tO5sJNjTAtTYcnrz2OIzVkOg40PSMY64yUIZHZuzZFO5pA6OK32iwRA46zmC68J5X1w2CpmiqR4u
faqULmoSUSGiP7TmS9ESK3pL6DBnqbo+snrkVTQJepCgeUunKryYKkhqDfwbtSUJHCETsMmN5BOk
uyfCm3EzppQeoWOwEUbvqYAyGOC2j2RUQe/vl9LELRRMrE2zSwQGH5O2n/wYvIHDamQhY5l8MV7/
NDwUjQiN1iiaiBG4TZkDSzON+K+8TFdGeCtnUWFUFJkBFJt/swa+nyvHWowC1nThGH6Gn1uJkjTJ
5k866YDZaN/1kemXZ3jIs8FSeLmCsh16ptVlWKUBkHEZKv+VuNKR/bPPIKVaFZOP/LVbbnMXDT6Y
p9oRyNY4t7Y9xs755xOkF8E+Sla2JwX6NvWogQ/5x8E09e7hSBnBIhgo0p6TF68kbUUL0A/VtKDz
mDGXirTKIrwO2UTmO1CTyi0qB/oC4j8yRHOfWV5hplvJ+7pmtqNnKEGsmhwuk202HnuoYJDwsEdV
b2nsHpgPv83vnkYLBAkH1CrLaJ09XmwVGD9sj5aZaUd0DtDy4bM0kXOgmr8gWYS/ixW/y0Z021k6
cDAXPqfeFQsa6Vn+FWaTQWJ298R96pmhnbFxPX5jAMVn8XGTpMPB59mzEqR/wpvZfBEoguHp6ICY
EYXHu5UJH9m6eKYyehDdYDiIZLUGG2B62dKIHEFz/pKqeHWrkDn0mqzk/5EvhI3WOSV18NQknzlM
IouiyQfKlEnSCZqhikH0R3+VapuokAlcXx853q3RVkQ6p18tcVtaxbtXj/RPqOq9mFrcMPCN8Ahy
Nf1hVHJAs/jItv1rLaLzeoRovLqqJnFLczbSxSxM5zgmq+w+xWGjWAyXEfRf3rtaGqllELtClP2x
IrbLz7fUreXaYJdxRwruPp7t0QS+7ZBLvcDTXIndNrhL7KqT3IO3yxAfT2zwmx18koW3QjpP4v9X
z9Evwbm23WwSSc8sa5I3I0U+tG8l68laIJJ1762+PWaOYECobiadj8577njKt+9MgYPAjxuOFejS
YIm/fHNI2facxgXR9KPbtZuRmBx0TmO6g5ZFGCIt9m1AnGXFMvDO4FLYoL8OJ4V402qcSIr86DJu
Hz9wBpwHPTyYf9cvHImdRzrdbytylsuttxgMmFql0s8aZo9CHunTGJNaUSj5hW/FCETR2vtUcml2
QOTYkc2eF+C7R911RNGN074KXZHKbsEohyPIf3PJyHWNb8KuMJ++/IsVDPB424+Egwo9pwNNr+Nl
bGD5Bjc+yuI1UDl+IhJ0lez1cU4l1JdvBJMKSU5Y+5zByEsQ9CYuOjs5agTXsnfo6klkpKAuXeMl
P9Xt9VFSWO82/piKKPJ50YK5i2lzDnWcODRddIEi5XzbdgNh+XsgLkXNRve6qMO2yZdpLJMeuucC
TVHHU05XoObnNz/XnXRKK2ouYj9X82IcWVMp9AdaMEb3cJ0L12MdrYTez20UE+xo7gdoyXcAqtPa
YCkCu4sz903g+MLIB4VGvTr16vmLvqjJhNpiis7lVeAJELx/AqNyuyYrksjZY/jkNrlWmYuvS+dF
XHmCr0txxJW972cS2DJPahRWS3B7NOeKFGY3xCSBMgk79sWudNxTvFKrJCO2h0T4vVgwhzfMlxPE
XfQ91rlQps46rU+aVB/rF+DW3vZZIepwXPCMVMZ96348Xij6wCfZPJ//b/B1fA1gohDIOWjHdFZA
y5p643555Ny+iNpmRJw4oAB4Mm26wXX94IqRiMk9dIaNdlhcqkufPA7TjjUNMH3IR5IgICrZ5rNS
eXLzUzUaCWVZUqdZupuEG5DUhQ/UdYxdgH2hFLvqq1yWdnko9DDS44Vp5W6IetnO6PxY95ZGUHrX
ASMlZhwI2s29zpsfBWVtNqr+yaV2HxgHNX2W6+v2wEgJIdpk5yw9do/p0Ghib3OQxy+rS+NC3pcb
7rGO+ktXAAyrgUYb6nO+ux/BpW6cfaqt8WCEq9frm8AWfur+w8T6btT8IDK11AiM3xPvb2HOlgax
hBHl17m60gPV89KXU8MYRxbyWTu2G1HFz9J1JL77S2Ljq8AZPxEaMNQGFKOrvKf5JXHfpxvYjXdH
E1OiUYvEu2l5m6DUKkl22KzdksOW7XLn+55ETT5Vq4AIjYBpUkxWRn7l/AkbwZVjlId/iSjkEwfI
Z7FdkagR3I2GcuH0epHnZJPcqOXDWABF5ZW52kIeiOlaJDs4Dfkxaqk6DlTIdD0DkUlFNVTeDV6o
djjZvoaCROg3MpRlWLIZoWJkpbJiYORWfE7FH4bw8qdQAHi49tWQtvrPTujuvRPz22rgdzuT4gS6
+v2FlbiQjU/hA6bpUIKAH8J8IsLjKOqOhMa6Q6V6Zmes9kf4hK+7EiFyFkq/DTshYjzIQ+HBLxOx
pZEnYvNUZOq0//DjLFy0DUz75NZpwgNUvpTu9CTa5/vVDWLmfDko8EIoLpg32+JLjy6UTgQvTPTS
XYrYS+Dfmd8G5nYQ5tK9e87XH4EBlkR21tpvAAwKus1VDo21Onsb0PTy1k2sPhi1ReeX+YO1AyB1
WBvvwR4VvWjN6i9sRd3hElSpaLa+TfoiaTAAp38AXwBCPE30dXoi+LZleBXDAYXPLAJEdu63vWmM
U/OXDklyzFJo/UpPZkW4XzkzBqbt5ZmwTh86XDHiJAzmGQcHrDXDWszpI2atma5tQlA7xtL2IUT9
vfCkodthe8InpZMidTEQezsnSqAWLHQ6IoeBx3rbSju0ELWegJp+jMbjh8E7LCtk8trHo5VNe0m+
AbyAW9TluIMZgJ+PkHH8ws/YGB5F/dMey6bsw9QWu1p9xFWwpU+/9+Hb3T3HJZltlNmdR9oO4E2f
v+71hNbJx0o+2DgW25VD54mFOpbjCVrebx/XmGCefL+xXtDQLgELxeOrLvAfNC8bf9eLkEVsSLKt
zovBe7R2NMPVRbwaZK8ft8b3dA1KjoGfszCkeJO5gaQ6+0+GAzu5Xlp8HayhaK8jM+N71EwUPoSB
NRsz1lGoxg+YhVIZZOtuI4UqZ4nrns9XHGW+2zD1uIKlhxiezxmYta8ADFu6ATbedYO2qdSG68cC
eCwRxb69eL+c36aQj37kRTATNSPSuLqtjFiAJVpNGa5QeOWcTc2+oSN5aM3/NRYY1PouHmZXqczm
YUpNgV943ItTzWN0jJlvuLdQjIqxykvWPzfGT2mSks9QWo337rrubtMW71iR2QAdxPwkfUKZN4sr
6tp0Ryb1/f2MArlEJvjIfS+p6pCg4JVQp9x4B1MrsSZ4iJWgakaqyVsfbzxgQPTGT86PMRQpz46K
vv5BZMDdlISCjt9acrGiGyAiPXB1yXoOycLi2/fqs02s31RBop+zeoH97+9EzearsfxcG6fOKmAx
9eK81m82Cgk5KdR0/uurjVOvuZO0epiWMnKTJHx2W0vcI/xXcK2ADHl21Ncfe0bE7aBLTFo+b8hn
5VGHr0RXGhWXZoJRgm+BNPHlXbOJ7Nvxl0y587cft/9smT86fIMzlCyTEeDSZJJMDzaPkPmrTgjD
Ak4ha1nhA3b1ac1BH3eyZQiRbd0JRME9ebNhtSckg2+XPx3GStldtCwEBYlmM8p6kS3ePMd4jPTR
ik8YsxmoOMQvqtfIB+1o+iGUj0DtbWisSZTw4Un/HjvDg3uR5qOVSbfrJ9qAE+QhJSY+epfLAbqz
tY26/upcLoKsPkbsmrGZknzcBDeQHRU6aVa/lbCTx4DUPBO77LMnKKNEmJNPIaRv2djv2uniRh01
XQIUip9lIKnnUlnkrXhnE41cq6da3iOt5mhOiHuUiTjO7Pa9WuTkVtILlHQzl1tXHBc5luxyZn7D
g1mhYU6l13aHPsDPBg7ww8SAIUQc3Rv4jGTXGgTTIvLidDO9a17eKMhvZUnt1nyU6lubpeakIOyx
ArvjeZae+T7f7PkyzIewyxrXYbHko5E/JR1wvHGaal3BxyhnpT+cNs3nKHKQlHto4sOPs6+j9wLM
rsCvsg9uxzJWRmgv74sEBGsjp/c1rXwdy3jX5rHn0rYWnQvzhrBEWlGMuEFr+tJU1OrK9MwzLtVK
EaMqQ8MUzVTsPRaWTM83DA0E932LsNlW3RzYCTSftm06dbSNTL1Mt+4ZI+5ZkoQ2RlHNkq02CZTR
l0nSUBOj2O9rPDlYfl482EBATAk72WpkuUgo3ikc8Oc/IPEvQcAO0R9J7vHCBwsROhlVbJR+o075
zyCAeuy9LnyBBStEwrbGbWvSqv/s8OvZrVb8uUSWhSKS3SY3ohghNhYY2JlkermkZnBl73D+1/nw
lzT0R7t9R/M7+zQ4phks6SvgrmOu4OugQk+PU2lxjQcqmgztO7fHrk7wLbirF/0bSEo8P5FvUzIo
LSuhHVThGV2x2ExhFtTrMag28cB1UF/JSA2nqcgueOFamGsJiOdcxgLw22oQARkyFDqch0HA4hO4
jfyeCCjvR/WgAlpsM6CwO4Mbw+408V4hxPXjrg20eEQhFuYkR3+OSP2SOUvA5wvVZp+CCRC0osav
nwf9bWYbQN1pKwf5A2XMrPIWIadubiOW4WQT6u383h7xSdQ+LDVgolOKMwv5ut4CkvkvvR4UB5VK
R/pjTY2CKn8PJ+/p7GWmm9wLZ0kE8iCLDj8WtN+Jnp3OIyndb0BtiB0zv9FSyKU9aNR+pn1E8bOf
ZlOTjU7qBxC/DKOQiXnF1uOrNV3YcdkAVHMPCKwwHVBEDjMnR4qI69p3N96DYgU4irdyapif5IUG
QGtj/UGSPawuhD2errJsmPisNGeNJ4Kw5Pxf1JgaycpP89ctuS77nh4ZDtAhXbFk2drN4AOiBy/N
oF59GOLLpch9gUWxxDSu6gcQTUS4uMdSOU0s5Q3U77IHGJ24HOlR9ZWH5NkR52knumM+SUZ/vdLw
EAllCYAf2wdIYiHrAQeJlmCwMdcw2Mvl70yJtNIOe4A2cx0evvYXBOi687rOprkMpfbArpfBICiI
pggyt8WhbqivNu0X4gyKejQbBbwTIj3kWUGtkql+LChESxGqxU26iZTA32jnGv6FLtStH6QM0uxF
EZueTD1nnZwiLrRhsVh8+XBwm/dTY4HS+NXz7gXFbq2CAbyhCuG6ZSMcrMDLZixnGj/P+1mlizf8
82nFy6rvGRUX9U1PjwQqiZaI3oUO+gfZ7iuZMwiU3aKKWSnoSJ/2h0hf1CTxHeFlT8euHaXpf/C/
xtVZbvMgj85TFUr9IpMvEfzi5u/yKLND+S35w+n3xpCLklBNvhmc4CQ5hnpunOa6N29EmilPrdTP
OFQ65j1QPP3x18IA+LpzguJL/8Y5cbt09ZjZ6RvOO77ciGiSlWFnNt1BGHOZYqoTWLwHjNEcZHdB
DQNkvXwnR8oF3SfMSvuigc/4h44+O/M7dn1volwUAMJfA2uSWKgNlhoz9foqCR6cM4xxejGMLiFh
Jl5Y3DA11ZylqEIxc1xGo6aRmjaABIA1IDw68aYAh8i4ms8WOzptPwPRf98pL6zk7t//ypDMt21k
s2lImObfDDiPA0ePAAK0D3u1Nu8u6AihHpdZMkK7CHPJc0+IwexpGE9pfcO3qqO5NI8cdNiTTC8X
rJ3TXT1Gj9hdxqrmPtL7CzNATWicRZ1vKAjQS0WF+gOJ2Uj0ccTIhFiU0HRJulv25IMx2/TAfga0
UOeyiQO2ovSG7DhfBtcvb+eFEGJ/WQFQL53k8ZrYK3/doGtZ0bwjHmhs2Kp/vdmPpbzFzzVetcq/
rctaLiRblMA01sXlYE7CkKhmQjzJidbmUd4rSLrn1/cAmhWVU8d7Aj+IEFirvARTCZtrINB+U7H2
CFaxJNL3IjRCKETyIMqgrnQr6zhWNfCxhyUYjwtkZcyCLUQvp2ewoY0nNR1GwFvIL9oVqcqt7Xqz
MlWBJrYOfrdW3R6ory/tKEKjzRJa642I3ugLi9wvVUYbEs5sQ+gNjtHTpgRoA7QduLsr3kI8k9AQ
UlPhBSvhA2a3sPqhDEbDTih1FFDIxqrAYugblB334pJs28GyF0RCm/j41yyIrN9gk4yZLlL8tZsA
ZIZLQuMFvi/qeujzcCGxT43Hmf38M7Ev9LY1IMF/r/GxDIL5vFuCLplT6M3RHIGUJEpQ6FKOZs7E
c8c0QIGe6iIvrHMh353B/YiWXbPdv/GtE9KvHeGSWoa3nnCa9aaA/1JxPy0LLOqRD8Pw/3Xfbku/
wb1Kte/z+8O3TpBd7yER8lO32wfLs0xQXfErjFQq0QJ0h+ETRMhBTexCU1YVaoneX54WbRcVQdGm
P0R/rpEuWfax39re66MQMUsLaXJXFz60SLOBnAyhzMosiXxRhTfAouKd6br1+theg3csy79m4Wch
jNTxtGZiOedAlzzzvBvQpXzPVwL3zBA8ooVKu2NmPi3BSFAYc4xFaTNgZ3pxUZNWJGmsinzL/kPo
tBofq58pUwTAXhVxal6ITr1nTZyNEK5Y2SENLNeyQPxrEcQLOLIFTfSpdg9Y+WVkn2KP0s+D1TAz
PIbZKMVjwdJw25DADeyZSA3kbZJM8ub7T0txyrJYvwcz4Ik2KJCUpf7vHrpXFuwYpKwlYG9r0rEt
N/txfuRzMklNjb6vgGiozIULzy62zyCrwwnlmNEzSVhUAo/yXNjn9moC5tDzLbul4TIuLsM6vT4r
spcxqqGyeqiQF54Ep1L/dz3xW0JoFAbWYUvZIofTLp2Pq2yKJp86lkTYMA1xV5bhdwUKNejN3gqS
q0kABvO5Jrt/qd19wDWFRB24SHA3LPGKz0zUo5imCm0wLeSBy+yyHZJ1FDLvO50FwzM2OUQojCB4
PRW69M4XPeyu8HMaQbAt5AoSxDLJshwS2sokdp9HQ6GzxLw36SapSlABFdjXSsw2nSyfLpoNPgD4
z1gr0pRks4xVPUnz9OlEU9vwVRCgC/tkyLm6Gqjoc2v1r3XAc48n9hXAkaFEa+C/Mb1RzkTlX9d9
RNN+yKhvjuYHXmA7qO3tomVVDh3J/dyfaDt6/iNf9pzfmjAOmpxEpeh2mCvLAo3g9VbjQRiZKKIF
0M+0kV29jaLKS//2gJgbDU3hKPUKDA9vgaZ9CEjAX6S6T05/LWeXV8liOvmGfWJBgR7zK6/7pCAl
ug4WHXlrIUfV21IyVObcUvx35qpiTTTEYFahiGMiZFbMC4aUJMaEmayRLvbulUtQAiXKia7NXxVb
CV7Wzrzhode4+6rmk3A2g5GuV3fE+Bs68C2qopSj0MBSogqaTmmt8uwPX0gQLg55U4IvrLtLrlL7
V0T61RaMMz7XD50y4SBk91K4Woq7GQcUH71uWfSk0wNXAUDIw0TN1jcByxydcSeni0olCyXZLs45
cC9MOIii1V6pelaZeJRnFxja+xHakA5eeEYAi3G2cCxDP3VUIIH/V3ZkSy/H1bhzAX/y4RCPiL5Q
zS330QluKWVhd3ffOw9CkHqlw4TJFswzMnGjVVYB5GV3mxfFxGUUj5JPdPuxrch/aQmnnkBOb8Vf
tg50xZKoTUNqESz5/Doso36ttsGAr6GyyYPLjcq4mRwLqy89cDIyBK8uE9zFycSIswc3DSbIkJpC
WYIwn1rNeGlnY3AoqtfrPcJbZ/Ti21jniSnrDEjPoy64logaTNXniqB6HJ7fmAv5JM9n+GllGHMT
3kOL7245wpssnkUcdCP4JzJCsebR40umK1zkltVGvVNtpXpTu9Uom+CDkS+hmNvDJui5eqUwxV8M
wVfIo5EqKyo9I9g3KeV/L3Ns9j7QNeS9iaGT1gHJhGj+bzjetsoT87xjIVVD3PiIUM8qV0vl69t4
ieuLtzjrOJZAB2lMs5ffD8tCyHErBpOimPwT2lrNAqjrhS+Unc4WvlbeSXlA1cX5ZvXHAS05fTMH
BETTMCvHUkf3MlcpU3DHDFJtA9I17Y7Mv3N/WCNexRmM0qwLo/6T27WJoXNHKHus/TfY+nlBDTOs
8CfthezjOIUvq/+Ri5SeFRxh9j5KKYjmvkhtqx44rGrIHD7SBfn84oGjLis4mc4XXDMR37M6pdtf
qZANnTWNRqq0wieLlgN48/4OcGlcja1qizIZkHjaR+M+e5EIesgRvJw/Wggyzkm6zZWiZScjdQDF
5LCPYyLOENISXNun6KHsxtMeq+BtpgfE1foArxIda0wXd1bW0LM/JAMtspiqdGT9m/TabCVaNMnx
D25v8HwdLO+2yH+ojN5RzE7Qcx5RaLrfGeW2sIchU4+a8pOttoPNnxp6PqVhN25gEVgSUkTOLSMK
c/vhy7P4s7Krt+VlZBgLVWaRyXwYOum9XK2LHiBaI7W82TKeFQ9IM5+n003tx3XUSWPU7zXa8/H5
2QlBkTv6Ie7DwmmlKPwZI2CR3Ij936IBmpxn9TK3jarJlRrzXVJvrl5IpvVqT13rjx5sl/KbIUMZ
nUaSCywAx8FQUorIwgcKzoc05zMYRgYynd5JU/E1NHyow+qJugg3CMTZzq1r2KQZyD+6VCljPNV7
aavWcxUmb1mZXSMTN3jgfjcCIBSVuKt1pHkxhgJf2BkQ2u4j0fkaTNGdEfoUmi7wrBQR6VxKBT/s
CZSk6fXpvHQkK87K4JVyP+B0vW/o9XUfifOqshg/7lXYkDBNkJ4M+ByjlKoPTQRURiN2c12Kezdp
ZLLR+0Om7qJ2OFB9oW4KqcRbIOIb4Akmtf6+6y8+dcgKktmei1mXgEhpcWQUmLzpjtCiNp8mkOpa
2xWYso1bw851xRdgM8UG+MD2K2/23kngx/ww9Zw2N9RvtARCao0LkR+a8TT08kSabtS0QrLS17Ds
RPs3esArn4WtMqRGJOOib5uHypA4++qADjN565CvlBVNtC2A2s4GBKsgus1Ok5yvZAepJgoYvwGB
pn6+9HYtZkTNm89tjqL5Nf+UWyo0wIZnAgi9NgscMqckoKrNWQ/Yz40PfkF2u4nigipLArj2DReX
dQ8Y37J0YD0hOu5pX6R4PMNNuqCaLunNzxUq1CovQumapjeXqcWOz8GpUaamBITP3gMyF5WP4PAu
j024eVx+I8SX3lXhd3JmFH0JMVKSAE0kNfdlQU6ROgEtuXbRHL9iAkAgosZHFmxZQWYIADSMs8dP
kkEGuQksmRr/z5kNVCWxrBwoAOxr/xmcQn2kXEJZJzC/CKz6YsQ0kFq7B3AKBjsW+oJc7fJAqC/R
ZzgHZI0QdHw/Gr+oZTchSuFdDTka9qBM/BXET0LzdZqtY1ovrRwQC4FvkUGQNG61MfZl4jFoNaTt
eXErL692Egxbcm2nAOygHUqyA8Z/l/VhW2rnjEAisV/+Kc0CWzDMc9I0DdH5b34TPDUVOn1le1W1
AcFUFg7AeulOLlwppJudAaVVB//QrlG4n3VHn5Pz7hUEp9oDo+nSwgyVB8MUHZNvInwRtRKXUu0y
O69msGWHcCvYTJO3apmxdcajY1nb1PH10uw0SQh9aI7PrHkzCHINpF9h35AoemWTDtcEhXufDF4k
IivrncLYa4xR7CaEk9mM6zG5qiJ5GrsAoRDDs6MvB31xU/ukHe/XGBsTQVLLZ/vH4LXgV7s9myGr
QvSEk5B5DQ4CX3T54oeE62kn9FoPxsCxa7whv+FNaGQl64I40FuYrUPIYEpLNBwAY+dpS1kE7ESl
WnffcR7ZKq9cJE2Z7/la1+LvVxB9HsuqSoHQAq6QV0I3sZUsefeaBi2v770W9Su52tRzgkhphBNW
DEdmr09bhjQvGMUDsHSuQCfypIDhcBEPXG350hyoGhhKfj5p97C8MTSUXVK6jx0LRACkCccODO4b
ea/kbpQ4h51GGeriGPTsflF0aYBbprFSx/EZIMW7FgRtlCz4g006OLepLfjMk5OvBSF8vfGeKzGo
32kFe7VdutsrENYgR+w3MwuTH9qItB4z2QHSzTAbyc4UszUMOmJrNFoKnSm3Z1bqyFZyprD4Lu+9
O1QdX9BGEWvlTrkmSZHvgeD2cmBOnEDF1EF9WYljr97flLKh8K1SELzIb0nuegA/pe1MoDxTwv/o
km7U+CNTkzb+kcbtBmLS6xHl9A7wvDodHtfZ3nz92sZcbFl4EgAF/dfy26iAdP7IjWXpFiwNJLTQ
jGTIGnIJEWeNIBa88UiQlhhhS3CQkGXONTlClzZ1L2Lku9gQKrg9BcPTZNpxTu9PvcGeWevwpZZO
OHlvHPEjUK8K5kl9c4GusMAspcHvOh2qhOXdG1W/RMgY2g4JmWxWnrVHIIgyxDboHIq05FkAY9m8
edzVNEs2Bii++lD1B4ZjArN44RcI6FfSikCNATlTCBUfc2MgVPFqPFTo+Z6otmNu5Qf2l+RPlikO
9HIupk9LSmgYzzC1AVLeRwocHDQAUdaortex+Uw/k6naHZwr01H/2WKaCOoIWwYWqNcOZSw89qji
UPqBV4xnFAXkDC9ZIg2fxjOxysPnWdFsjMadPTkdgSKSkj6mFAgYcukrfxu6mIDaTwG/xhHARA2o
8Ymss1fsyh5DDHrHkPqpnD8pYVTYbE1M/rwBAUPPcS/hXgsq9Mz9ONVhwZMcHQrFrx7z/xGidkPK
U4wEANtyDdnfnjJ+8OqsEufEgLGsepycdUUWHCudsbyCupFUzzEwvyVpb7biDTlRhnZieMzYle3w
G7V+DSWrTYP5wWwkx4NRs9d1jJu3pL5es8trF/0Pa3jhl4awt8OKXvEz/eNVWNKjndf4FF9WaVXm
jUf08r3mAFiAOCcDfepQXZS3pB0aKCkBK1T9piNWcHcyRynoHT5v7I16cySckN+QLAKmAbAbO93Y
B7gAE0O5s+6q9m/ag6EMgi8x8zPYeAC39QomF312UvstGUjgTQ56cv3FbKHz301Gv8bIMvYUs5td
yipAKdYOFg7kHCgvYPVGIfJgZK4o2WynsvAa9LZPuv9L4+U5tPJBcRkx6863jLvzTxFPPKONA/eo
s06ymXbiTe1CX+fxT6LXg2iJ0LnRX51xhICjGfZgs4mZSL0nJF0Ar9zBJB+Bqw4ps6l45+XdYFyH
A+PAq+++m6KnycyIYicHLpBepf4Y0UdFEWzty2xBIr3y6frx+joDFdAzKMEswCilmsaVihAUEOmd
CWAq1FThOsTYHKfr2x8u/9XpXQylJKLxBOZjVymvtBCHTbm0oPojWqkVsGtt1l+HxVIo0v0WVoPP
RshG/Sx08TqpbIZ9A2OLKuWPqAeFuj9qcZKAU58EKoAtDsIr53PNC4rbu3BOJSQxz8eRih2DSr5E
AQdUpfTXnLvXYzqBAVnQIBEZHFVz5/edUKwgR3PsYwU77tlfLAp7rNWfiZq6E0BNphADndVRRIF+
qCifu+2zMUKAK8Rz+UyPSgDzP785OJy11B3ZC8Hir0dgD0rDZAUTnEvqOmY6pkk4eB7y1v264Kq4
KdWph7D62YZfAhXhs6mBsEN+wbAn2ekV2Q7s0l4xyurkhQYaxJRZHghTTsocncvqq8jEz6ge4+bt
zt29t0Dj3zqZGKDaxJK8EtatQzLX5VgntADLFpLEbe7pwSbmgQRkJiS152V4Kg9/zFa4Qt5EuN4g
WGHdDy3S19qn2Kc4CJNteh+PkHIbmALYVnQXTlfVKH9Z/WKKAE7qZHz6GW8loD7hz4jxFZeWNT+U
rq2n/PQNoeMmntSOuJ/0WrYaSMyDM9sQTaJjBah7i18A2FU/jwMZv56/quGXgg3XTTueWvNf++bV
637KZIpLmA875WflMj4PxCfc5Kz/gcezrDxBL2CKRsnw4uE8TG1sPPk2WHK5+wtKtELTpFPRo9Po
ICNdGNY9N+D+YSi5SN7l5YKTLzTUPUVTS9X7F+pRRGXgqXl2ynuhAKdXYO4xFU+CSxDZ3HQnRKPC
88VDI+oFlM/bCdkCpX3mRq6wmg+98p0TCvn1emu5IQ1Zz5bAEHV4xpqEq6zhycBM5E7wBNdO/9DO
+tHgDKKpwY4/INf7jk81kgS3zbE92ZgG58AmA4B6A+NOmXiYwZGEhmjDoXtJNCI2FRlYv7/WQ55J
kNVzuX87RTE9iqlGF9iZRqw7/Zr2+g1lJ1XwISDrresKs9uWqrRiVLuAqPuPXtcEtD54uF8LxqHF
Kow5joDRMWJ3XFNh6ITyYqQZYifAxhIw06MHLDX+JLbsJ3QOqmb3/l4P/dfUyzhK9XURUf3aZzWI
C0DHz6BoidZSZ1ilTSdSLBqJMsZqKbehmN1UMKC9ln1L8souX1cS1DWaWwzrEIBQo8ssYwZcdiir
pD5r8E0W7YHYJ8XV67M6FN4ijVJ6dWaYVQRA2LT48GlRpOfE5glH1cg3mNz2OON8Ov9WcuDKw08Z
bNnGPp7avzivJAR5tXlk+fKU6RmIAZZjcF5L6jC6djKtV28JctpWeZT9TTJt0MG6IjpAfyC6bZwm
RA5IQq43v5/iG9IBdRaKiqne7DTC4c2P4rtKvRqP9BcbyzBXDW0n3EsTzrtLWVWo2WcpkvaIDYxS
vEBLnN0+sYacWzwT/cBJ/10LvzaOD6huCduDZP0zZy2hgDULGVAvkHU2UreO44VKYK8WjEUMWxPg
a6C0nL5FIQaSk6Wl4GgzIQpaTef29xsW7LVQneXvS7ooayyuMCii/knMn+mJ/CsPdrRHD6D5RKM4
l23FoCkmDFi6UKQdMt0FpbXyNrxxwejjvZC9aVDb6kCcD/2/+ajJywWOkNrmp509ewl7L74w3+N5
xrB0SkaoJc6sJKbZt0p8skImo2h/cZ7/Ut3vGYAQXnkHL8vJwe4wOtW0FXqDD1h6R9gEdElqhSON
55+J8pOWlMKECMBcXxm8cAluVmbn3Jo4MzhB6HR8oDedl9eUbYBRnByg3iATCR2yU+FbHiXOHNQf
GoIWtqRsBdFjHbtmuLhlrBkKZANvv8J1Olx5MfgDgLvofiUd9HrvQgjckwgml0dj8yVFkFP/DpHw
36vzcwiAaA0mae/w2lAbQ7UAf2df5CBVFplqS1T4DSXDLIznqMx1m2FkLtDtTZkOT7asOttqXK5z
xxgqYaEzcpCecRYsF2PgFaj0UC4yzqCH/nvCsHw/8cG5e7yvJhGJ6mN+y1bA9kv/YFnKIuYuz9my
WO9ZR5eSQurRVWuSA5VatXp2Ncbm+eFgsSIEHidNYZigubLIrkBSj+vICX5ei9k95chDjeDI+IIr
u+18SEs+ky5Kq1ZwVzXKRkNa4b5Z78YdwG2/jmNAXGZmtFXf8Y0GDCXw6wqGDqc/gG7tdqk8rnK9
PiVRkJb8HVH2zdwkc5M1yvwTMBe5j0J+UuW4upwjzH+LLl5O3X2WzlGBQov+fQ/sjZOLDUGKoxgB
JJOFIRhhboMEZZzmynJrwOFa/9rSJUH2ApMIV7gsk3UfPtSz20EQIjW3/Y6xDpZv+r110750YIDx
QCbq3tZRnzT3tDpRGS2fugiI0xjVTgDWQjGUxIjdknDRpSY37NNdotWeelAdDjSKxq+vqoW6muiD
tvw3QsgXYa+zIetbHOUtHSY780isDMn20jQ3rHz7KeerglFLngEnAst6wgdoEta8/WJxkVqVDSLn
Befg7yF78ufAfFIKpHT2FVe1zu9D6kc08bvcUuuskzbV8XB2C4ZR+fZxUOA23LD0wMkAbYanB5qI
jwKfNyNVxKnfrQOx6F/HmN3Uo6mKnot0MP9xwA5DrKtlAn5co35uUER1gJWL6+HAbR6hrXQoDKzr
7czh7GO1mJWXkAbzTojmo06bVljlNMAhGu2UGMdjswIPcIonuEpz+35p8wJqvQpKYrrH2yFmTAAL
is/LS1bx8YTuZq4v7E0+dNoo+RFgOM10zORXUBQZAYKgvi087xAyYtYOGadGo2livgbh1fCRupbt
2AYxbMJ2SabXgkch1uWnaJow4wDT+NcCjYH5ODr9X9jEiOJJm/enA1PWTrxQqVOm9RURlqwukAsi
MgtMMfzoPwsZ5zFy64IEBlPq29ExTcEolElsnwshB7Kka/KAsiQ20yH7KxuSLJdTvssRuRoptotI
qxC9Jo9WVbIimllXNybh1hXsWdyIjAqyM4u1ePd9U5bDq6lXVLiAenmqbPFBjALLpxTDll1xGR7b
b6J2rkMHISNWsTzD4518D6vigkVFYS6S3m4Y5jXVYbzvw/VLwOYLK0NJ3lkciXKFmph07qL356cg
qMPVug0uLfSgkjWGLFbNBHG8t0US4J+oSIx7uRdvfzsLepmfXeja2wl6fsyuuCLH+IHS5tufIz9w
rRwUs7YWBrj7Aem5d8EZQWO/OwPj3iSfOYBaEmyGIOMtXu5kMRZsEr38vp1x5Kaml8QWTg+/SaQG
XSYAOSIfm3o/UGZcfhhuna4jPgLglKZjcKir3k3hWRmI4x26i+bvGHyGHV/Fia9sOV5MqjaeeqDy
axrley5KZ5+OZhwUP4RedYsK06wl8uqjujwtBwkpbECc1r04yZ6MkxnXemCqdt9YO1/qxllkwaJy
3IhUoBLBWUzgFU1gX5+1qOJXziNJFDkFwQ0LA7lCXySd9LCMMG3d5+4wmR3h2Hze750NBfSf35eH
74tpHd0hLqnRtCpi4UL9SuVgfe5FY/Fc3rf1BHWghxWICKQ4dHiBnRZhVTFC4LGkowds4xofOUTO
YGz2Hab3OviUNQhlrxp6FDf9obXUr8Y8CnNf6W6EwHEbbEn7t6NSddbjNKYLqeLKIZkPQ7U1SBej
0gXOyTeGImhg1H9ZPQZrDOepqvGvitnFAeIkuXQu7JsN2ix5B/f00o8F6tykFeWNydnjoenigoSs
nn+HjoIb1BMnNQkhk6ljV1Wzx7BYek/M50dvL6gTDsJFdPBV7Yscll3AtEqQGQx0iEpPM91u1rjS
Pz5eZAO3tpYkkbS7Rjo4pZidIWvFby2OZnnwwU1MHx6+Dynzo7E3VD/4lfe2MaYQUAPqcpy/8W+e
FxMiq6t+htqD0/TQNvA0lIAxqUOeTc7DdZdb7AjwaYM3hpLF6e0rxSasElwWAB5KYixl6dAKK0RN
innJVM49s9Rf808TjwY+fqIQkMPsOaAEzQKKl7FSvl1QuS2t3/19UFzuQtqRCn4WmA4s4CLsc5lU
mUjxGHLBfWGKCNJCIIFolcxUAGniJ4vmdShCXBpDeL4PfNFFAwvZdegAzhlxaEnieRmiph826xhy
OT/JVt6+y1iShXCRiQFhZq+C2I18uIZ0IV43g9Otifo9kGANPk1EzNjEQM9NG8zK/S7eKYCOAWMn
84iZvfqakLb2FxNJD/ouzuBvaZvM3tYNIigKs3Nsd4jKsktERtc8VuQx+ztVHVt3TJfn2WTCQHxS
WLJxtJbCbyGxFii+GpY+wrZMqV1yRfWXUZGkQbL50MW3xpCki2iTObvKkX8zeFR3ctb9KoqqRyZR
ZQAFmCDBxi6O/VkbTqgDOewLAZw3tyUpyKWsbDtJkfurKuWXaQku164ughCTX2fy4lKqJxPZEsI2
GWqovNL2rNOJmhsbY6iWWl1f/eKsL8xdxnUf4HGhbOqwuJdurwyxxNkr8TRWREoGKn9gZn28KYCC
2ay+vU1SZcq/Q741pt0JxNqz4B8qJ4D8cEfRtquFYg+W3SncCpgKzmrM0gGfABuy/09gOIh954DR
hJ2IufgRYgmDAEd9w+7RfJOFV+DzDQBiauY1irZ1hZYc5HDKpZEUC27Kk2TtxRwW6+H6+rGC+8V9
fJzbRxjmh3CYwB9MDiXpL4Pt70GTzRRjTSXxLYT/+kIAgOikLfahkOzXfAPEvERy1CogVMlMWrJK
ltVWKlA7oPmHe+JZjlPPzhRowqtXNkwabFFsXZCcadrGbgLSvJcZ+/NQ4ElyaQ/cfFK4S6SGnvdr
ec5ilJvMop9ZAxxS43oVMBDORPvESFPRqWNjxfdf2j1Y4lbo9d2XAV4z1G6WomodTMqhSvFIxDX7
oo+e8IWnmlTmpK9cHo7hbmC86v2c9uQTL+6Z4qEE4gIZMIxugy8i8VY+U4KPEliLgmgjsQkdZnV/
I/7ZHhVDwyqpLL5+QM/GtEU+HOUV+jaDNeUzg/YGsEBFx21NaGOCOP523I8hMqlzhiFTBLs2sD+R
JNIUQgQYBuuYG0yPGuDyNldWKwrhcByrm3peVZIrmKYOks6dS8mAzKO/w/eP4GCDDCLallov1q4O
9XIBfFTfN4rc0uoJTFW4z9LryIXxO5BLbA4qSQ05EMYCqSXvO1XnO6fgAZvvd5Bj4xU5AOH6gHBq
J92Uxfv5pchO7VfSD3Wq6ALOGsgBcHfuGbFZn1cefl/5BYf8xYynwpyarSjH7mzl4i+W5Xs2dQEN
cIOkVp9PtFedM1ZGetg+xGuwEt48Yg/uuf/CRWYD6UgtIMNVtmjtFU+l+Zam1/E3FhV0Sr6lQdBZ
PVv1VuJXnxHTYkHCucA2r0QREs/RADM6cxYzYIhSpq9KhFzxkh3ztHj1hb01SyqZ+4v14KfS79Gw
7YIStNWTHYSE7Qm+QzT8KdYj8KygVAZPth0r8JfJNjjH77ajQuS0DTpyUszWIUlMSZ8IGcd32co0
9vtzkkR0EeEjqVWX9MaEBsqDacH+n9uqyhrzE/Utja7skbZIXUkeQkPz1MgeAoFbt8YmrgVDh1XD
mffrb97eVOgQmjh77e77tQZr8IbA4erms5Lf0gyJrE25V3YMyozyNdCwivV6TXLJ3YmjxkwCWuYZ
EX2YjXP6TC+KEbBwLX5A10d/8ayKFsbuqLm92eFJBaOBfOaCWRrJNMUg9D9posqQUIviPdq7WcBH
ylXdvHK7iTxhy8tXgbcDd5avZN720FIGEPrkl7k+DF51AfVJnLSk0/eORiIwh/EVm1IEJxS3xnYN
Xf/I7f+NMDmKdfnrBk+cgSbOAVwKSusQ9w3yabwBJ9XfbppSWhhT1iwxqi9p3PCN3Vl+h046e6Ix
b+oKH21qNRXbo2A39r1CUtJboJHE57sucSnAF17lnGsmz2SfY5JBP36LHSdxit0HEorU9oFl1Sep
UcLsBO908drL0ZnYg4ekVuvt98XR2XRnfl+MwOUpN0W1qHb5KqdW3C21dyljt40j37eO4Ov9ES1x
y37VXF/jTJ9R9rsmWrVPEcm8BKE0dZVQWiaUzZsWHO6RCnKnCjxPQEGOSV8+e6OnXLZmy8EZFJD4
/GLcnPbl9AoMSoFfzya60YbSw7n/lJJcx7++cl73XHJy8+cfMZBf5E7kisLIJVHarz6arRXBESj4
aEzpFg02QwpWUEC2Ih9eYZtwU/iPuB3ooFXjv0IvG1KOn6uzvomLWVoO3lgNbu7mlDw4UeHWSE2y
aFjZNDnYidXGh4cYOvolJV3ycDBYNU35CV1eTCj9dMQAG1QIdlKhL3nxRThxHcoiEEMJIycKITwg
o2zTRTYAynhTDVMZBNB1GY3cXoEAvL/8840xV4iv3B3xEIpwjANYtVmOrNt1ncoWjPzpBQRT1AJy
Cme4e4p9MixcVIXfIB2PQf7FLB5WWSKpU6U2+GfhC0VD2NOsjHOkcUQHbL8nQzQ905OTbSszdE/+
+A8YI8B8RIGgagnzxWJbPa3MtgLgSoG2vrGQaRW8F/hNZKqZnKB+/BY4DtHtMb7BKMTerg51T4GM
CyRJYQx8p3A2dl74URrlSmzGlNw0demHzvHYePCX1AVzviPHaGNfy5HKVu7KOFi12MB6a8GPvTPS
Des4UoOaAvFwowtrCLkOWmfMZYcjAcahpTyZOtM50DzmAvQ6ok24+HHcgrmdnsVQl8osnbCz9YgB
e89m5t7ghIVAnaqKdoDUXy3m6zmegyqHvfWQTNP2YALFDFXiuxCRg3XSpu00CpdWGEzrtRXVxli9
fdbESPHJJ90b8aCuPXLf+uJRjjBZ4MWxSKDXHqSLJjU21VKQeTimw/X+Op4Oh4IJGgsfHmKVz4Rz
aeDMey+o2NK+Tbq3IPCR/Y6asaDdmwUSolIpbizZ2wB70UNiAUZvMStiy+c2XX/vb608yuQtjbIh
020eBsrQUuCgMbK8QiwFlCKUl6Kz0nQLJ077wqtcHDNIQ2ek5U22opcwa1ng3lrtmA8nje1NxPQp
a+44pr+RcjrT54Fv5b6DocvWNNX6F8aKZIoBYA2+xrjvhB4LRNk1XKLlFyKeXQaelVtPA8hfU5ml
qu5o0wuI7n32gzbP6nKU+x0d4gLfjcVyxp75gweHysEgOytKTAq3wAsO4KRUPzZj4pC6msbKASJP
G4Pf6ZM5+n78jyTIWBCmoKnvINMAj8IV3VUg1Yp4imwNXKOKEz8bJgB2lRyf9JC0d2Kilnvc3tdz
csUrOk+Qo6I+A1FMAhazUfASNYfff2LJdX6RXgJvRJtoqD+KtLGEM3e6MbW0rYrlut+08WPrflTX
FJ6x10GOdtZX5/ncWVTMRDYJSMnyB6xK7961wtNnhDa7iZajB+Wzi1c6I8k6dFOFBewuqW1veAK/
kSRtNcXruZWvfPMlNmmDyXeuarZ3+0suu3mKsvoCOq2vHP30IgG6kUJunF9408yuf8PN6EgdlbUx
HVhSesHpvtAwd7Sp6EINlOVv5F/BYwfwt8nmQ/N49ljBR6TNVMyW9OOgzk78rsTDW5z/T1Wj16mq
cI0hZV0Sl5sonR1kS7NjD+G6SHWwkFdqfvQIr2/jjbE3K+eEs8l5b6v62IbtZjcdy9MCYY1DAwvI
8lQhmifovqTokOGyFWSZBU71W3AVhi5GzmcK+jzoD0PuQdtNL49n0YdW/vEu0nQwVvupf+CjqmHs
50HlMM0PxCH9w4Sh8mtkGpKnnlrSXTTVZ/R3yt9epmM3y5GxJAeVIY4n9hZFrqR6QwbHWiJdBiUW
d+ROtg1gnZgbDqJzmJZ+gPHmKy9dWA7lqaHRqYv6hCrRX/Xb09oTakc6gdYFMedY6r+tg5S8AWQN
3IsLhw1a+1Ci74jgkYvpdzvfdQeQK+5xTLS/t8HRzECdH8zriQTRjyP53gcLshKvRHtL7CqxXRRK
Td+Kst2RTRJ2YpZkcq/fifvinfs+p4jhgp8npww5Wendjz/+XY2ryKmWlN13z0oOz6kauIaMv8Jw
if0pVFMy/DZ9j0JJUQrFemzzZ4ssCLELThA82VkFfjqPpq4+DbHGdE/fQpyENLL1FGN5jg0M9W9k
VKWfThgbwoB7yi7kUQorWEvHsM1K/U9kGfbmCyNzYKfA1x5jTTPtPOuRoRBvgAjlmq9cYhD8A20G
W9wr01bKSPcdMfaCCC92N972p2NiaF9NCqTjLGtKl57jhVpGJLFBFdGpa6NMT0+vYAXvTneeFlj3
mMfDB6OZxkGQYZj13onTcnpC8E7DXoJzKAzqgFxOzvyi9SDILXjD7lkWbUu4w1O4loucaShocgmI
pgra4L1XTkp6tXpcNp/OxE9Zc919lgBYHXjTI1tZLG//Wkn9KtKB27yIsGg6X6N1KEFwd+ZfvvSg
H9iSNWmew5gIVSZdduq102Bd08hG55JPs9aN3E15Qw4XggPgQAr86n+yWMuMATWa/wjj3Yl9fQxW
MYUl/bFNGsKcBcRaxwXQNR1kZjpVfiDH0Cvzojhw8lIcY3Pe61GjH0zL5J3ZH+S6Ku9ipbd76ATx
geTVR+GySo1J8VIcEWXjfupaNsc/T5PUO+MQRyZkUc8LAs1g/NF/pcqzvZ+cu/usTl96i2bygBFO
NhqDdbo2glB1NH/6c57/y3tjt1Sp58rUkHeAxkw7qpH7Hy0ORCBsrs3YZ+q0dKquEfqyPOIX3GcP
rO/oafrtKe4ERgyWO8D1T+RFdqrxD06scXkvwJaLC0dnSeDGdoGQY4hgvpKnC6qM3cuUr6uzfEGl
6QQ5oT6AGnUE0HdokMnDU4wYzV1khAgVz8vdU7vYwurg8K2AYZI0yg5b1yX8Dbyo3PW/XxqJONX6
7XmoxpXVfAUucCf+O4Um9QYpaDYqVXr1Thac9Y9PM2Mz3wckXF1RG9OGtm05M3TTcCc8eiH3NXKG
19tsnfQXTwzIMzhbMx15sfoE9ToBcRGHJUatOpdLo8e6/0rKSWXyiachCX0mCivXn1KjjHGrUDcG
INYsFSrPSwZtN43AhhkhIqZgiV3+nC0W6VfQoSNP+I99Xp0VVd5yIqSirnVf5ZIN0o0tlGNIg/7j
A/tpD0GOazFfm1Hj6CFJ7WFw28Aop2BCzK0PyObWBP4LsywohKF9fFVlxR6h5/EF0ZeEKYmQM8Gm
zc0VnLRj/hlYWA9s00YVkvWyznIHfuZas8ktzIZPfopuRvNXLdmSkrshRTFay0AkXBQbA+RqU7YW
gJfdeSqMqh5aL1/GQC3QED3ScurDpigCK5vPvUUnhOI/hfLn9WRzT0eKxg2bJ0CeBx1t33PautW7
c+ecIsRVVpu86SeOevgrQX8ikJ7Uxw3e2dtYOqnHKqg5V5lwzpQiVYvsaJb/+Tzq1s7Vs/cQiKWj
cJ5YComu5dVgDD2D7CAeQFbjiLOmVCJlAPJmnstehyi/IlBud1JyePZ1iyY9ibZzyEeQiIGg+Dqq
JmoX7gh16GKAzGPBEaZayJT1FmS7mr6UpAbSNlV9BgMsY0uHzOtD3HVJ/XgvZY+PHxXj4IZ8eTIh
NUcF66rJu3Q6NDgn27GHCtpqLVCNH1hupIcMuc3Q9T3VbC5iROdWfF7nEFHxjKUpU4X4L0UweZY+
zzizbjALl2Hu0djXvrmFE87nXJqoJgPPhvrRVAUHaY7QZEdPfi/uoT2YsLOv1ifoalGZVnOuTWB9
w6QbyFle4T12S9VR1xUbVnO3nYPyhfV1GGh9B3QGSH88wKf1fQt8AaS1LRmok6B9FjUd6R2hVMKz
LC4dxjRLfOI/S3C/l6LJyCOvTs8lMBnIgNB8yGQaKhx5KC9IFPfId4D7W+T6rEePsYxDhgrkFW2u
ZrBrHgNBvw9WNzKszG7GFZXOYqU/LvmToZRezJiyR0j0B2XNEfYTXwL27rJrjDaFJ2GWo9ApplQU
IBFZw5nkJ5bCU0QjhNVhCpYeDJIiEbPu2uB6u8kOk5vCBQ0KD0wMBhcJmpFpMxYMZ9yN4l65Mc3O
hiMEL60JsljZSh1hrIYzboh4LWfJ4blu92YTxToxA8o1FwQh+ZerPhHADOV62nCj4Rl9lRClQDFb
iFZk1Wf95JFxf9tvf0qKz1hRJFYAY/l40m5j3bt4N7TqT9OpqsTJJGr8VLEZ+zxR9WenW7FhQTH4
F+qT652avMRPSPYW5pXbB1ZD40OUMgcKPCbIfaRzn9j0FomVW6vP7Z9RhsiuwRBBdD4MJcW95wQq
0mLLK1bfckPcxGdvyngctuKthBGqC2vnDogt+Nat9RfrS/snMgriwpjH1UFvLg62/tsaVZZCO5i0
HOtTBSIr9eLZxaxvHqSGbWu9Ghj8sCHA76p6gyum8BqG2exYTrd+UYjhA0ee3jxJaNpCBVBZSvB9
bF8+WRKZmGFaJSu+T5dv9WWPbKqr94+V0Yj1iRwBNszPXByb6d2ZXXejzGsVrR1yydQ7nkaVVgjc
/V0rWk7VJk7pd70alyu3wdwr+HmoV0uxvd3+JEqpTCfLePQo47CLbPpXQuAFm2L8c7L+xO5QRpjU
AF6bcWF9GZG+QeRsU7NAae5UXZx42uVe6Ef2ccuAdZrpvlJyaj6Z8ZT2BcRtO77+2aKyY1N2PcuT
u/RzWxyIlroamkKscHMu6R0KgEo7LxVsiYFOFAGHP0CDRZ5FjFcdGbpLUIBBx1OPN9uDhXil7SMP
M2fWkvpgYTzaC/cqnaRjrVnC+mC8rEnn9VG8xqo0UscuIcgYyphSVdfq4g2lj6DUITcPhHQyt4Ax
KexRlFg4DA9YETbTs99yxG3CsHKHFPnXW1T+YRLmy2haRbPpGXvs4ApuzUHryrcqBg3YfOEFY5bI
SfIch9MStZc74cwZG7KX4HzYQnmrtbaY+ydeMyd04oJLkvr91JsHZ7QK6HLEvFhnqk9Uqh4CNqgI
KrK/imrHs7JE5RctVll2mOY2mOYf1P1Z1TTW/2Dx4CuY2NlXp1w0RyQpeT2GHGRZ2Z71BqR5LAvr
MXyyqRQpOllGBqy5oDyMhm5+2XusdZb8UxfmG28JJbfiTa35K24vvvQ2AvY5+X0y+bjzluCdQNIb
xmj5au1TvXdFtGpTETsJEi3hh2Ns2VoEjizYH78AqUiZtCY/cB9DByP3mrzRqIsbSoKemVU8BflK
2oNFeS8anWpaMHKPpMHTuonaj3wHuTeSG9iXFz50xc83+BSc0avoztKLPspfMAqYngcs+VC92HU0
4r80DskxAMLeaTqLvBEqXTQQKaQF2RDntKZSB06PGb1BlKhAC8vwhF6NiqNKFogRnJcKbNOMV41F
9KbNe5YAeh6yBo75ZfZjOWvxoCY3nTal0AmWSwxiaLMQ1ZVZ07olidpW2jvxR2ypiRinEOLofdOY
mbjzSCc1x4ZggKKb//iOBhNdTEHNp1UpIiO5+ZdOLWKcB/fQxhhPbEyUkA94NqZ36Qe6ggIIhENK
R32TTkSbrcqk7OwQ+R6mgZV5uSwBKN358MO0fENFxiBlgx4mXrMLGqJiiGlm9eNdqLnGGrosIyZp
elXUZUZ1AbyevGH2O15hgABZA7eJ3qTTvGoXN91P7PDWUtIFOzcHSdrVJC02ZjYtBGIr5KD8nFGq
GnzxlEkgkrSy4vyfg+gXYo2lTXzW0uQ2qZ5YdAFcfnSU2ULdNwG0erBgQuFH5i653KZfYFwc2bSm
xzKfGWkWGXmcsY9M7NiMKPI8+y6H9n/XQSO8mdjFWz1uzvh2AhA8f8KPvuMVtAH5BuJ6BO/AH1XH
Yv0GPkk6M2qXtWQXBQu4RTKLq0dbD0mFAXAlrNZs7x0qiMIVHVCHk2mTdyPQm5b364OyvRB2rezO
T90Eo2gZziduTqfNAKcLf/FEZ536Jr00VT8RKU0CAfHrvawotbFuisowiRvLEZtGVgWR31Yl3TIL
d8N9LOPJr5KiAp5+KaJVEbO4pEJhoF5VbQnzPby5VJUI3rLaxnOeVSWlwEliI8TFjHbLghFBU4oE
g98deAin0aYWLHL65eBDt2hqb3NllvPi2d0IsL/zZtVmT8gFGOimpQUO8vBLRroEMCDIVsrfzpV7
iuD6kLeIvw5SvArZ177OkbGIjcQwwqN0mgu5alVAmb3hOuakqjUI+WiABOo4pbHMHbmNlrH6T2Ru
TONf0+t6O9hTKMg1y+u6tiETuo56oj3hmyCF3sUaOXj5RNnkIIE5X0kA4ljFhF62xiRZfLnA+sZP
+t8FmMTKfog61YQNaIMQC7mYFNGgR2DHPtUfKPgf1I6SHN0q9+lE/N0kvEX1m9vQICXuibVjr59X
z7pxt3kjv6tV9BQeJdSDgAdsI0c28R8roXVptgvJ7ztyLbMbZMdDQEA+nnax6msM0tx9igFDLf6q
nd58feNJCMpLvUt8qCQRVn1eDAZrj57nobluSdyZ7vZCMnKyP+1qwSXabZQokNjV12oYrol1RlIx
0fNBvtdBcHvU0UKb8U82KemOQTmslSIHSCInXC7jvQvtRoBlNu1ai3Fnb74TIcM2Kgqi3LB19hgF
bf5mTb1gqtQHZ+EUrbZDHjKrbFCn5emw3B6wA+D3H4R6AbDAFIRhb7ZCF9LCdI/9dDBxysGHisWc
zonUNf8O6VfQ5l31TBfbsjaaC7D/+OSgK4hMUB+MTO9M8AsHhRTlu32q6BpASDyt6idbRNA4lsal
uVKriA0lrvxKIUzlb5XPv3Z7qHhnm4WGSNMnsfa3qYd9Hy38wTZcHvUqf4Q60jb3aTV5DCSoR48M
JoEdON7x5yLsqkM1xi+6pzB2KLq0+4ikAyJqPLh6fjJrHlF0pvaSUiaUZOYxJRaFM8ezHqll66hX
nUYtVUzfvhe5Q0PTv9GvXFb429tfhVKtLS/f5AY7r+uIewKYsI7pJFyG1gQrNMnUrHUBrOF8dEof
p0lm2zIKC6Q+f7lOA/SXOB9taBF5oYDrwtYttHONdEwp54akkOoa1DzzMo89fm9GtNeXQPajUwKI
HFmZIeZlfvpDt28sRR2k1VN7/7qVfyKss4Qovk45rBdU3eMmujwcEX0hUs4HpjB6bz+g6j9XH5vA
NFFd782K3jGfIbSj/wt6astGzY9HnB1sQeocHb15jCATaXEGItLOO2vzlZgXBGXR8YrWeCDwT6ej
yhDxLd9xfW1Hg7IxUPREW8ZZ5n4/Oy1dHtRc5um/c9t1Kb3RI2RtegZC11q5dTDPB8EVLeGEIktH
SFLcf5Bkz1aOBiIhLXZcf5GYRdvAWocdU6YRJXdpVFfwnGZljJbCab//xgSlncgcl2HbcQ47E55m
yLTaLsD3whXmsVlA9anxyw7t3dT1ELOgk0QvmaRwK61gCTCijebtFZ80sJtHjfhXLqv/ori21Y8u
p3OpK7JP2rVZTzaQY1ykZRIK16mV51wycl6YtAzCizvES0FQImee4QNCt1N8sl7MRQZhn1960s6p
DVCwzULiqNuomFma8Gwr7oQMeV5tepUiZj9zAcNjFkJqaNbwObXOisEdpfg8WMoTPAGb6wkBXffk
jgHhj9WEdHMGj1JcFrHXj5JWE3+QnWQfFpHHxocapamxMobtImVI69suQ/u65c0k6s7u9zCBmetA
8pESJqmovnUBG1hkJF96U3s2cky9jrL63sdZFevcy1AsKbuyC9GS93MEiyaQAnrp6Z7Ea2B8N+gs
C4kEQM/cZEeC10bSQC7hq/Fn7zFbfde97osCzouZGq6F6iRSlrs2bDKiReH9miXVwITWaDahJ+BK
pNse3z0BlaiorJU9HOKH/hXleMy8DZvqsNVtJho/sz5StN26B8e1Hwz6bQp3ly4jqRlCCG1lnuRc
bjQGYgULAH+1wpxCIqeE+X4cPsLJwF/fpjkNCJwbGqSjms3avLLoxRIpPvIbSNICEMQeVDQRaxeu
kQVo2h/lM2dUBIOvXKHQvxxerSqdGzgjJAATaYoOdyWoBZOXY8jxi6qDOCgtEaUGFMFmgMWOvyqp
mQbQmBI9CdIKVVXdsYBxyEbWskRtUvCp0kPei/3OUdFGgFdvLB1DyeuHQiWklOkalkMarMzga/68
b0Z0FoN4d8WU3LC49rxQNUSBfNNzdb5rdyJQDEZn3iKGJGwvJQPlaey53tXbZYaW0BA+eZE3+mV0
2nTY0XMAf6UO/WOZ+ofRaqURQ9KpfFDjBrkaH87wq+L0H1IApl85dkU5YFT1h45QYhRsNbYR0L/u
uVsS/KHf9ciMj4otd02CaeruxoJARkqTJR00X9BUwzp/aWgILxnCaYrDerK1Ju2rMSVELosc6wKI
HmOoZayO3fk4KWq07iLjK0sfhYsVsrsUw/6KLAP9Z2vgbJ0mqzbshcBCCc03J1gGJvEtJXRDkO/M
s515N3xbu9JNK0MflwMZPWIVNEqZp898IgYDknhq3GV73ddwhWvVd3lMmFl8dy5RtUd0b3Gn15Nc
jb7wZOT4CLKPtyBhF3+9wXqjo8yYI5iEK2Fu51tz+y5KmBSDmNMLFhsuLqLmx2sTb8zW7TyMGvlK
rIcE4v8k+I5ZEksV7t8Obfmgl7jaH8qLxfsnxjSGLgIxG0zqNKFPVD96eHqbmwMy5ZlOjqREov9T
lStSerfZ8yt+OWlhN7QRZVTVeG5x+OrGmrUCjT6WRITtgWanBkeWieBl2MVmiQjxNpB9LOppnG0X
pFh+AxZTK0ACHe84CGe+ZQpQKZnrB1eaZs1W7yoT5Hf1BG6/Yx1/aAjX0EiJYLlPef20cHVqLrY5
OZj2iCNYeVBU8Tn19udAu0VuUjtshOWR4Uz2NqMwDCUU/nrQhvGpbniqiXJa166eXXx5sHbXkO5A
OjShnu0bW/wRBVLU+U+lE9Agty5ff5Mx/2JoxxhMfhiR0uoaXtmnhpwcv+XlgNqcI/BviImasZQq
LLtrQVvtTMIorAt3T+NPXV0dgfW6AXG0n9vU8qaDVls61X5fkBBAx080VURplooiOrT68v/oOdDF
25bB6/38zviGcmw/QQfZLnvhHCUh2aIovDm3TR4TPxeLeMqRY+nCrjs+EmVXUXa/+MJtgf26s3mN
FL6raxcCr0Q7UC1pBnJDt2pP4iYKG93OCeYe3EEuPfqZy61eM1gbmm35FGGeKgN0hsplvB3fBEZU
tlf7tAPX/fZWGv5Szs/EW4xqVG+nq+fsfQ05APxEgw2xw64jOHGGl5MmqpQBuJHM0TebW5PUaU6x
k0o0FgzXQiW5u7Zjr9V5YrLzFQJjtmS0cwe5w+Bj0DVwAAwaAeq1cPKWKfNEnRdFMcUeoYVodmWq
qTvQ5gAGOVy5Tjgj+KYNnefuDjVFHjLHd4cUVlD+mjXk1gfs7JZ8W0B6gQkoRzbCyASuRjyaFFr6
cSSa3EvdOUx3mDsNNeoqI0iXm+UrurIQXZh9yjcnKHHbc8nEhCMNN01X58JdLw142I0HSxDyKsUX
8TQz8NBfKAMo9B1iLcuOqmbp6Ds2GfZ9YxoUfzuTJXvqjtiqVa6w+GOslrK5iBRaohtLAhXffQit
icIc17JKttK6CS4evp1aoY/wwfyQjSB69jp2ocwkxEuY5OUMCrGmUkf98agM8HRHdbk3qauFclzs
gc0EBKm9QTx24YtljKE9iP0wb1TjgQdc4tXzs7BAK9gO9fST/W3B15KhQjoM3+naDYix0Ihbw4Pd
+Qn/myWgGu43BjVDLVKQ/+cSrGmLVsa6siO9KiPHqETrV+v5Ymb2OsQ4L2G1AYrNRAvCMMCnRlma
EayrE5x/LBrKMWvUHZvCOmCAGF+9jqgTDnrmPfDgLpqLMynoShg0S1HiDNCEghqiCZV930ibxfYG
ufMQHrQ/zLYEKMR786MtBT4hECT+s0CK9l2P4YTDV/9OBhyZ2c3tRBczK0SQ/cKsrXmBA0wyB6Gu
CdidoWVg8zAOKuqsxn2ULqZgSSAW21+lbD0sCM79AN+8NObbLFS9d7qh6MQLBIHZWPSL5h5RhbWb
8qDB/RhTwQMteHBIiLgLlgOow23NpAYcdvka+0swBDevlcSHTc/QBr3in6nHv9XGVmGyGGIIgeme
pPLZxlKSA56N31KLGO3TrY3CFk7rXe1hD3xwGl5DTKnhEACiR/zKx/N5Vn22qTJB2KrwXWrqGmHN
+u/SB2IymwpiCvAc0yQ1EgmyLjaLxRUaugUzf19P920h1mWCpoluQo9/c2bFOMRHGEjvJomhq7DC
dGVRrpD1s4PvS9pIsa99yta2/ae7+RkF+DEsZf+nuiQbK+Xql1GSFY46HLjIlfuvNqT5fOcGzAAf
dzwgwP5t78Pf1c2HcbL5lNN7H2Nc3Feb/0TiAHIjLXezzbcg6qSus3u5ZEsCuR6MagLX7Zd+SYFH
HoX0Y+GQoBnrqKnNNcD1HgWSsJZVN2kZ9D8UJFHLXCFPVfsDgDwTJL+6kZyhHWUDMIOpwtCb/o7t
qNG7VBr4HoxX/lsYVIP2w7k4JDVUZBTDSy33umYk37vVVBOrzFMRBQd8+2aURv+OGL1BrNA36+nf
xsQui1qXnCkR6aCV0/OP+DItvHWJCDongWIJ+d7+IZKQM5bvcy+ghumL5YmvfRdF6zmLZRheSh0s
oZR6SesyGWoBv8roacFBOaZmbBca1CEhOzb9xjNf2cR2+/SS7qE0My7nCEmH5uyfqDIgByXIZqTQ
ePQqM2bksm9PJP/pbfgCf7G0mF0b/znGPM/shzkRf6LVBRK/13FkiD6JbGt2P2pfi/CHRtCu588o
IlN5GIdj9MPh4lsKhwbts3MOfZ+E7O+MphLXy9IlhfvBlMadmcY8Rv3QKR+IZzthJADefvOy75y3
MkJCtsS7XSYgBXh1CC436eKSybAsdFrMgPH/2cQ5FqTu/3DhjuecQQAS8KTt0CKoDu4kCjSAJi2K
KoCaKTZesEuz6CX+8ecG7fwOt+voWUPfYf52vIv0Yr0xXEFlC81qmKoLT9V90ju7Y8Kr5TOpf+PP
JLVuBbL2GKH4jQWY2I7vIJb45aSraWEP9U7Ly9KfLfW1HkDf1vXSV/L3AWWLhpqG5UUzpUZbWdF/
46w3PKidC0qXUm0omiEht/VO2x8YIjcxXI5wbNvW+QOIMNv3gD5YOrgBXr/3XM73RGcePub/DKwf
15Vn1wjU8aMCJ+ef4sxGB3AklMgDCqFc3mFuX6I5dp+cXsO5RZ5wvn4VAdOh/DbXbH8fTi0qLoss
Nd1lASsQj6rbR8XUNIJq5bA+NpddThKVdm3YgUggs0OTVwolk5AIgB9qIN9rBmI03dEYlVufRwFb
511VKFt8qRLHNrr62uZ+pRvDJL1DmrIS/Nuv0swipJQhSbIeAd2u3oI14ZfbfG+cf7KbvA3bKhE2
JhDBUzM/U2CkxsaQQqHMkfLWHvhkv/0xbx61Mmwi/3nyt2BXMtHFN8iqvscLAPY57dEf20nQ/dX1
kAPFEJ3w3RVxK7qnfW5/b6XHr06hTIFs/CslCsSF0EEzSXnuvF3wGVQq788GIJviY9s763iNGoHr
PZK03BDQku3CqngqDbrKpPlNJ00f9BzsoupW//hpmlVr5F4/09XTmoOH4a8ciIV6Lz7QxE7vOeOZ
MjAyE37IGuQ4pSqG2cxy2wotJvIcy4SgYtPOs93TffVeaur3b2FKJ01QPuJXrDXgNQS3y1TdDpnH
4sFBZSPYLpFo7hjw4xduWokw/2bpIfokxvE5pk8IHoVF/oVpWVUrXmnuDWAQrOi9Uj8epRU2jLSa
zyhKG3BHg9z/snMCGBAehzzbeQUxubHNAFz47Sf4idbs2L2Ru+EHjHDGMOnMQq9mYANvtL/SSsMI
x4CUnsXzWyo24Ds63dnqP4hNaJXWNUj6LGnBeWmB2Y1t/frxwXCfO6/VykoFeF9P1nYE03WW1Ofi
YsbHw9neh3tTnOd2UDQBDA0Hoz40ihC8gfamhwWlxB3UpKbyoYA0jzFri5TYu39iYL/0Vngrq+vx
oFq8/XKTvkexoBqmt9XILezMLUHb9u4oHlwO83Go49voIxFei+ge19HBuD0rEjk4ucofNQYEmsMW
ZAIWRXldXPumRV+HKM5xQ96CY0NynLKY6uP4gQ6nXrHEFvfDpqGU8h29KHB/Z+bYlDgqKMjtku41
viZxoyUQ6Gr2S2WjHMIBNcnoWFB5SelL95RZKvTLgShemEntJHuVHzdhlV1azwNKJ4CmfYQQeTAs
qYkinITnqJpJIQkje2ztVqi/z98qZjIVcLDcu+rDPazBo5BBaz45KXw4lXzC+MOmzRjizbtB+7o3
1a55NQCu+b6dRTLXH+mReZBNRNNC5UHVUCsKTWo+pDAr6jdma9zRjqSxCAUxx7V4VvH6R39Ome80
si7Xuq6AMuErWDv8y0h1YIMMS2rEWY3kw/D80o1w/lqOseHvpUZDfHs6njv2f1FqAxKdUTVeu5R1
Ms3pIMioBHpcqGrcqRFuTwNWCrJLa9Y2q36W9BuhbybdZn930owipV9lPsp7N2DxNIAmNy+5gadM
R7sEWZmnHnZR/NssyU1y5JSlue4uCrSz7MZX8LUeOW9cre6rXlWAn1pkUkhTZwmJW9cUpAdGGHsY
vyfcaTNPQHd8bkZeXv2l4yCfY0UeTE0lMw7nLKTZ3Cx75cX3K4qFjU/giw4SKj2pVLK1GyqFXyZI
1rkXBY9Lcyoto7Y6+SSINLbGUc52/Cw/LkyiAhTPQeDJaFNlPcO3wtwVGcjt0SautvTvuZa8keJS
RtRnIt2l8T0I5fdQ/n44vNoY1ADmTZzi+QiBKEqflSUduIuUfRINfJUTvCpW0fy6UPaUiBHzi3BW
ILoL+yTnifhsDtAOkAC+ASkEJy1BV3Id7uOX4M7T2eYngnKTnk3gh6K0ACSHOJ83L3p65Ryt4S1E
1XhXZlmUWrz6APEwvYJoyxYkVb5bwxT1nif2FxUa99kzFu60Zuq+l8E/M0cOfv+duQYpjjYDdQ/K
lQJIM2zPT0S6gApwk66sJ5kPEJITEiDYkwvMWJiU5pw24zUmHPavx8kJsu5sMoz831xnls7hbjL3
Nw3P0G+L8VDbfG4W8pf6IutlHIVd6lxY6F3a24E1ECFaZv/V0AsQdbBFeIYW068DrpWSm7zqN2qQ
ABw1hslJBIpPmbqY44NDrRVr4P0hrIP7OTfkXPhk54mCoHdvWb2YUJdZy8AHy4R1QV7nNOMa820j
nQ2BKVrcYzGo5mZ5yWe4POoTaQ2xuAc7aTWy3egHV9bjZ+fHGti5+pCGPC9LL0H8tta2k0vznxjd
AsaW+8XiCv47HMLzi7e/zk3oHC20cBbTPbbKKtZS9dMeQ9tfJlE0GGF+5zmsVD6ktZplOi69BD4L
mJK8c21o8Bjc8GxBxHR3+hrz8Q0GE6TwIjKzhfAaKV4P1n/QY8+RtRywO8Mndu4OBeVu0MISAwtp
Recl9CWetS/cceVGN1sM12Akh7IDgDYyNbt7PYJficGbM/tPDc1wtMQU5KFpreV7vuaMiRXnj3bu
O+8JxE5Pdxdij+VP8Kj9JZK6tzKpylww1BdhLZMs6i/Peo2D33RAWT/tg50wfN/FkdYFndufrQKn
jSeKq39p2g8zdZkgUxBQ94fLkyZTxLiUrkJpnfDwI/7UZ8RPDd5MYfqZS6iPdu81PBJU4+hzzhXU
8NAJh3jTIb3lbAwdklMEXwsE2zT7G8Mq4TC7leaFyZC9EXHKSbaCylgwJ87U62Ql16f+fMoxdHol
sxSt9E4WmlzbL89hUNO41CKlddLfXp1+4zSi/AOxxx65ZxVu9M8PKiYNNbaMJFrZzqJ9CCImLnUk
M6GolsaozyHgVu1lI6GL5xYfopmwq3WAkWcWa8MOw02h0aljzedDjQP4auk5vUaWiwCy6MY3rpyB
7RcQbfiCUH7sU77fS9h9GrxiwbyjNT3sfdSdp/RxbbHYd/muW1iTV3yLelPwryE7FliKACmYKUQl
ZtBAh9CI2DfsYnnAetQtYFHaJEd5ptj6iAT8eP5wpgCZ+HU8G5Xu6dPTOC4Iis3YXV8fe9e3LRTR
25tU+8c+qu/U33Y/68e3PhbhFCroWM7ZCA9E5QSTM9uEn5NrAzKUumnYTmAEmtUAmDVrhKJQSP5M
zS3AVPyCPFyjiHoem1h3IPm0W2PGW/Ncd0ptZBDwKmDDg7w3nJUvTLcJrtKYfTuMPa0y4ICevNNw
G38iWMir83VBxEQ2IDw0K9bH4QGTu+r7mWnZvx14hPdjIF2mcHvf1hIiYsPW3UjmJ0QTXcWGvSoR
2v5T6ZAC6P+zKVgQpv1ii8TA+BJvG6iykRJHihipRuudPkqrIb63o/uEH1V0oaEMXOd33fNUGFKs
LEdzCDJwPY0GyJ8/7A+TpEuGPf6pgT440GoySBS0XWkkj8yzEaxNKpjh2dFSZBzBidDEyRqQpMzi
2ZAG+IYP4KRnrceM2uB/VY5VkF4xYfbJZDRGHLLGZwskCp1B1GiiR+v01P5lEoNmhyHrg8ELxa0J
eH6hxeieiUU3ov2NO8h7sgHtbtn2NSHvgfTZXxEfSltssM9wV+b8hYc+BYndY3wJg+WhyLvyN2Ty
SCG4hU/JArg1DxxCsty9maJa3GrvCC6lWA7a6trrDfhA9+r7mhppukCf0wH+vhaSfamYCEwDOFT1
5pAU0zKNoRBJaBGDDDjJKS4E5bVJ0dPc/o3NHzJA2cSzCL6o5c8qH9ljn+49/FWxf1jOBXcbbB1V
PZ2lt5tzzFP6I0rj2gONHuACVuXAuncjyRKrW++97tJvDnjx63izG5pO81uRR00uaIXsmhOf+62t
dpN8veSvSuQ+5pwNaBuYoVYOEWoO0HD8/6j1W5V3F9NV46lnS4+PZGAUY/ye8XdIu1mzrtEf/2Pb
Dr0evppKvb9x69dgqsyXkmTcSk8E5PoxpbLdwcRO1I6n6WpeaXTZQ9U4EfiG4ThALHOggFWLTXuY
wAmcLeGXFL6Aqa6xweBVmRf8uunZvjAMvbvc0yrkfz7R/PTF221zqs+na5gciEAd5oy0wrKaSiYX
FOfehOoJO+ObdYIDC0U2wU7XPhcVX/KBM7kjPXJ4BBMYdZu5QHDUtKJDF6n/bBs3dRjKYAmPeOLa
q+neFhLhU1nfiikYzMxZuo5hbWvsd3aFrjRWZTMHEy16PWNBGeejQNSZ3xwf9E1EOVQTok1BEKdW
yvveVTkZ0yBgPP64SMds2ZmG3RiLFgKu4DKOjd9wk86yKfuVKreKST4cSmN+N9/i/E8mx7JzngGQ
vrEU7uugx9XFKg/sWAYMJ/XMY2dRTulEKh384cQVPjHaZnXhe61J9m7tYvvb9o4Ho5tyjpCk6c6J
M2XdH3VtqixXMwq/4eNdXcX9JBCAJAmfbJ3+jeXrjPqaKy3+9bHbGWwoQTq6Z8AYN7Fe5LtQJuqs
SvkhFGshxulBZk6q4aTlkhtD+FwV8r6LIOIn/8+jFWhJbnArBwPVDDbCIadcEPazgZDzRxqpr8jy
xVrcUwXBWoy6J/HynjdH0wIBO7HbS5Jtx/HQYELlkuLRu2OxPvPWTBV8pUi6snq09DmN5WpL6Rwo
pfpKznYKkFFM8FuK3iSJEE9zzHTHZI2aGIFj2CPYbM4AOd6rwsJW3AGZWzMzo5CmEaAGPVT2Sdwf
iMaAg448IIf3pQc1GOQ6KLmwa7iw6omlWLFd2F43ZeeJ78L05abtxPo5aa6ts8hD8eAWyQd2MEjH
H1OuVm3eZXCgDT2kQ7UvcJHlWGJoXIzYKCLIh0N7LSLtHcZcjZ+nzdOpefD8+VOAiU6wnUogGVDe
FSg+IVtwpdjMQBzKJt4CzniuIJJ7PWbRn6se6a2ZjvpJdpSZEX7z4nxfhpI5G11cumRrCHN3A77f
0sRMSewO++FMicfqmfxJIjmK8ztP++9zx/0hZpMQcnV3evIeILqgKyN+aW8nS2KuIOP0RvsPDqWa
+8RPxNzq3NW5Mc4Fa72nMJe9ddg78FD2TvU0LCS4goFjMc5VRyLQ7K356i4x0oLvPFblbNYKtNKM
RmmDcVMjjCEeFJIaDegWEnJBAzM77qpIAGIUqQ7K/yq930aitVWH1h0BRQOEF/BhAeb8jsnacXjg
w0qDW2+Vzwzmo0YVLa150icZNq7kBnOJ/N91zAQyYsYJkw8Y/lBsZ0uH0O6+pToxulsk+9BztFY1
+XKmVYbipLNVWHTZRJtx0J07HCsGPS28vKd+W6Wvs4qHmn0f8QgBjXdT9QT8wUrcFr6j5ELS4B/l
kiqilXTRC4xYdGSz0eSpUc5sfKDmOImehXL3viYrgnfrNyCYX2pvaliPa504W4D7nGrE8NLTrfI7
7lGEYKKStxvUZ+muIZj9uoseCp43XHVuOAK30Q7TAYKxW0AXphakwUNQGKM2ypuXwJDXx6anmwwy
MjVsye9HUevtWRrKDqOGxWVEQakpJi+RgQ2aM5ywB7K7syu24oWMGBgqU7SKuNp8fzcA16UfZLrE
+hv0OwXOacLmRyTrRZJEQqC0Oi/Gc3bYWbw+piItqhjA/az7250GjS2BJ/UszvcFOJHcdAYZVwbG
+X7TYOE1l4oq7jdv1PEwAKKcEUY6vBvXuWmYWXYpwJn+TvFUjMoGvjIxRaE2g/uOhVMjme4fwvYF
YBCyIRAPqnc2zt+QoN5qy19DCQ4ekxkDDwdpznXeZceti1g65xzVd8Fz7iRb/N09/3IymZNXLf7u
LWF4Zs9IsNWRkfHYNw+uAGATTZKEa1aoyfsKkGYgw4pmsJWmfuw25Ru6o+dH4mPAMS0jJAjZih4n
Azft0LiMTjqM5hUVlIkS+zNe6bOmVgiojKoELMXRZcxolV4jqVJosrJDmRvT+bztugfpqBN1EXHq
djk3kUknI+JQiYWYojhb4fl4XDETrkUGPPtt4ysOnWUlGUcS2yazd9Ejk6HpY0JvnO889dtNN2Vn
EyX2XMzT/dUjecaMWQDlRhJBa6epLQG9bUxvjrDChCN1UIo1D57+P1DG5fZrhbEs9LhqXrilDijj
LhIKwfC3rElx8CmquUXzbZgNBd7oCHFYmdF5kk0laYTcYfuw3ss6I1+sNasWlNvRX14B3xl5T2lI
N3WCdC3+cDfzzJRXMvOlGT5wm0Oxa4EVjhaseZ/bGRrit9xZoD6y6rtUE3hcqI+PFq5AtoHmO0W3
EXxG6O2/1hB6+f+IXj1na8as94zLpLMlW49f3ZZbNXJImU0qOl84QObs2fYX4Ha4buF/nryePCnO
6aDWYF6+0GuOqWQhIpARi+wrUzyi4+VRu9i38nIrB+vwRy/Ewr8DVWnsUgsikHyKQW38ou1N8WAp
sI8xWm4upYqU1xKZCI+UTM4Ord/HnlnKAV9Y3oDeWPojBa2JHJH/u0tNLFz/vJCsREwXG3UD700/
MSMyQGB0yv1p9pHxIafvzNKjFwSD8kC3Ata2PXDQh8oJJU5fpNJRI05OAQOVQfPrqO3sA9z91d5O
Ld0h6Ssv/T6caSruSN3TL+TG8B93MAVAfuyrEjq942W98vOXIcFyoi7PE9EnClVWkinzIIvrvqhO
CDpxhuBqG+2BiJs5y6tNkOR/qTTxPbV+MN207yquEXhNbHBwMNRmFksGA0GxZeZBnr8aW0+HFLDF
aEty+mcsyJi36nNYvIckya44ZDul8m6swjJ6MLRCaGvcLp1Z8vdko8tLo5443hcVlapFBcjnzRCX
UaMV5RCTfn2pl6n6zm49zDnNGWLXDF2JGRw7HLSsRQqr51Tm2dLI6jDUS8q58PTkYOt8PV3LJwGa
rivMOZCGWrHvc6kBLMaerPzazoFEh8MaZK0D0gFgMpluv4izYECv3O5YF5dr5ZPE8qPnG//uE84u
IMLVBGBebTXJ1i/VXDqIBjXbOfJ5usGi16D92fF8gpy/jriqVUJk7+3c6BwdcApsFRL0l+jBFG2x
ElK8/EfVmCUwkd6TfpB0LWiKVVea71Dv1gsNGHYUXQwc1TEPlqnIG22MwEvRxaXxL+G6xTWp6wEU
QPY9Y/t/xUY4gf2yLSVkhZg2vkvQnfSC+/zY5wKBUdFZ3VjLBv2X6KcB9ojm3BfbaWe0D7/hOxg1
JEDZLcOamemjLoR4E8c23qkuYR8okpogS7LefosFexiMZq5ujEaDuoC2aw7Irnb/86g+Hgs6lSdi
drfujwTNBb07vJIbIY2urxN7gQFaUifk8YzVDQWd6NMKfGwneWcYxMofJEDsHrf5PTxmwXYvpFdK
sTEsrFmokuweBD5ebprgM//LMyaxcjMgtT+/zt+9J8I481rDuOeGfu+3TKOEY2Q3D96J7CnL/tM1
uFAcvgJ4mEW+ZJ8jQA4+PuGP7vgtwKGqaY3CBatC1U5czUbnDTY3s38kwx8RJ2g6ldRpYInAXBm0
FfL2avwHkGH9rJsPcwGGs8iF4lOEWELtUuJQ51Z3pdaC7Hg3zMdhmNptUi9EfEFnHcVOrDCJ/rhG
P+DNhCRzYQ8UfEbHUAQQe+1zW+CBmdXiztxw8KfOZXIjt/JMg8goJ4Dn1nZYzd+Xuo3+dl92kGCG
Y0Xn+p2qiIt7NPQ9NjMc2frXXT+XdPixkL+0n+q2LojadB121y4b3nURH+/SrYpbrEebjgk4tTsI
7iMsuM4qrUEiqBTLBfz6CYpzY/OI6mBZiHyIrKRAEZuULxqP757HEKDKcUw6TxH8IOP7OkeQMF+F
n4P7PpY8DE7UJTlA64g7YKPka9fOfOai4oDfeSAW1TXkJwbhoXWAXrjUr0RCXiKSc3qzl+ogPvvX
IIOV15wQPSMYLHuSTLvm7eCXZZ6KwycbqFEyBmMnWZKAo01YrZTEa8dsxNqMwJ3QSAZ5PKenRMDf
cNIJUy3zCwphgNTa/dSmUtI4orXs5batEt4Uq25r/V8k4HL+Jw/U9dURzOHgFhhSELmjevwHBJRO
FqtVHQhQTcbbTrm29ohgFJB2kWyrubKvmizqP4eYcd6D6FYCQh6SCkErh07oIjBKdyKb4IT06wnV
xMDeRUDesXqzfjwbja8eKM/kE3WzTUrPMUIpfaue1/NCwjZ1sf3C5fW4CY2EAsLrk4upkNrkpNGG
2q9NrfyjC8iZn6L3CrNkNJRkq9T8Nag49jcR6aue467EbSqhvXnSXGVkV/JgW0EOVg6nh5vLaJvn
yKz/pWiLlCHc9wHRUQAzn6vBptgVojxCXs43d6gDLcILHhsPG3Gj/qZtPRZg+9iZYusPDbaRPphC
4VfAVUUDUEHjQchfqUCb4t2A53rCdquL3iza9JieS+xOpIg3lIomQVPD5zBEovn4olHERGd8ORK3
CIFXPpOb+x12fe7YgdZYk7Q6FgUZDjHp05HfrzdViMSWabzN7WdghNxjX14DhRb/0L1oG667ys7G
gfs4hVQvc5nBNQv+I47/jDquaJtECN5mbhRvLkK7Ntl8fbr6dI8oOQEHep0CBPsNuIpcFi9athw4
VrMdT+PItMtXSoPeXyIF+ftj7+JqMSR2j8aytAxsmYjVoebdpLJ8lQHo9nUVWiYNhwon32HP2Rfb
CKrgY9J4wxcspx/QAIhAngRGrouNM/jh43ilAUEhinzBCX73CAa6iktbNjywBLr0loAtpKYU+5Oc
gIFlXnukes6R6jgBnBc7gbLoQLFJwmq7i9KK+Vo6+u0CkF5ql4U18tPUpOfzgChFp0yRAAwbjlwS
S9DMXPM8jFxY2Vig7Te3lb+dY9l22IqabzamKUsA+XZ8E0w0VXbL2SGPwt0J3FdQPULhJ5meNQXw
F8zeac3s5VXza6rzkQ/C3PtjzV0WjMlYXwn7Vd5hmZTGqnrrdSG2sAylkofXDMcn9NU/sQL4m9vE
aWe1EdBsW5cqV9HEotPjg+mAA4mcWT1RhPIgUWrZWg9JHqbyO3mH5IMGgAZOXAb32OZ8XV2dttXN
XiqPNMG59iDrqGIznQHGxF2LAVAOYZ2s9H7CXiRkOryc+ehPisnoUdPPJCoqP452rbfz1BBUflFy
41B2aaQ0ijjRHBq1jVGgdCVcd/zF3x3pGk7sB334u5k2dvHTDvDy4LmN27fKP3bDUxhgpyyqhO1y
vUtQeaKGJRj8gEDJQlgiRhokuHArQppGY2B45HUu4zn73XiRFwJLWEH1az/gTKtu0xKTLg/IbYC/
aHDvU938j1sp2jSZ9R9yVJwcVEpWRc/SW9wiL12NiVEqDCQsyAb6x+S/seQeJKiHkZnueUB0n0U/
aHLsN7Q2S7zinfeYVhiy+DWa3P+j9SybgTctdh2wunfHymI8xXbv0LhjK4J5iN/2eCd61Y9OKV3S
Y65o9mkNWvegkovAM+18RH93kXgPs5NVRyjBopZfIWTNb7Wm44hJDmFvwYe/4mA0sqRoKMhShYBY
WLwmxQZQM43Og0v7+TrzpJrupXvpgPPlEdxzU71RsSNcg3VXlxRXx+xxkW8OgpZYq0TPSmOfoAns
kdtngxnzmIERBMwBqFND8QivIXQm46E4Kx9jK/FQF2syzwQkeWw997DNRK+56Ajb7H+aUWKUTSPr
3LaoesUALxQbMPNjL7RwKxPBXuzqs7fGOBxbOJJu8IAoxnGqMV8EczROeIdUyFf/TAVvDEdK+kyo
fZNtWvs0hLcXDQP9HMig1ozQ8QW9pf7Kcm+x/OwL+AVCwWdGh16CzN1CSGWhsuB6Dxh0OXrJK39f
k73V4yaM300SBtngwiBsWZN61CL/w1lfLxfExG0Hg/T2NbfVu6uYFN9Lzb8VXqNB1F1WysevWi+j
ALmSc8L/skby5k9ZOjWUz0ltBAL5bifz73jLE7L/YB29/blLps20D/iJ+XC14QnteVYZ+bnKsEn/
Zf1kVCrDfeF9Bjj28RxYLaWYesik7W6RczRDQZRfGXkPgwjRT5Bi3dNk+fyaIQ/sLJrhMa9HhSuA
IZy8tVHvdPy+Q6yGqgjbMCj+bPZLEYacqKPM5b02BvTjHg7gLOiRgd+eChtlEXOB4CIM7PVQe3tI
txoWIJLyfI87lvR8Dz2P8SRR1JY4N/tZg46NyroPCvQ1Bn4RbtS4thWhoU6UrRBqbqmlmQkn2jF8
ccdXXLaOzorw0SQKSZknOgOPXJcbjDW6ICrGulS4idTY4knDpTYYLWoWKch7zoeFgTCiCEpPpNU5
PIMIvjYxGCxkIenPkBy+qZPONRJjLtk+WOE8TE4ebghc///RqL+TepcTZVhb4qLfssLZx4jHP4OI
sKttHoPgBQL/mVjp916C+1AmS9jgkE+ju5TSthywG3PWORyBohPAZUdwW1p9CNIspQBPUKTuBgwT
aMF4dGbytSWrFtsrckcJXYXpvVk5fqOPmtyZ7J1sX/SCfJxUMklWJ9m1VXB/mKd4FpX21tR8jfuB
6x2ymXnY4YBBA8UjoMujYMItDfh/aAvVuBlJqP+Ovjl+XhQOs/SCqIWCvWUPXN/no/Ar6GHzA4Sx
bc3dB9vNUbVft9P7UoLUw7n0XkLj5PcyqrAWSvrCxIQdJVs9gbfXLO/FE8wrD+wUEfHOryP+Nraa
gz5RvhkYfkEVdJLOE1BKuKRsnU9r8KDE29ImjCWkR989OhgXjZfxjDXTsWEb3hObSZACBc6cAtup
g+FM2iDojHKIbcIeKSWTwXai8ndyGzWYvM57EAVGpvkFkpwdMksbN+3B6mRLSFqgciVDmjOZd0hK
YpfaXCQ0dXLKMBXv9NYcTyOqHuaULTJCtQg48fwdCghpzDfFeezVbhlZRYk2hbqTBH0Nj2V929zZ
ECGJQP+Krn1F7LJmYYi2zlz0TFZS6SX0ukZXNNtw52cLin3zh7RQTY/aKC2M+echdjfoNnrMHbyN
Wk6YOVj22SZYyDddH3BY06+o3Uy3DDDmI5kUZC26J+n1M/lD7byY9V3J8cG/hGqE67iVFwnm9tg8
BUdSeHyqFghrlLbYd5700bh+72QMRWR2DkCYUaQLSQEbUvUgRWDq+ca/AOw6653IwtHPSgLRYCQB
e+/m1TLF1xwsjjUlxBTd0DAWWoGm6gjytMUtWRo/Tlb+sHfV7M+HKhFd79nt15uQx40TsJbfSskv
5GIO7Gci3mmHtU9ZactZ4XPR8rTiy65mXHJZ1aqRZaEVND5x3FnrwMo6ix+7KizUUZwKW/xmCPOo
41JQxEGaJHC8Xkb5XCc0wE5w2HiYPPlHPo1YTsSFIt6rD1DrLzGEELKnBQgluiPQQqmJS/6+Z6gi
op+bdWYzuuWXoybsJ03YwIVsLERtdQgsAD8Qn7NA2ebmPiv92Fn4xkp4TGIupqTgjpqC1aqU/f0P
f/YqX6PixhtrT/Gv/fWNIwN3hVc24Gp6r2XHkYVNUu85gCZEqO4ySiErzfA/MbsCWtDmLXkVj/SG
LGVKGc+xnVNx7ppMhbN/zweHlfsOSuVW/jJ0biogORRZe4qI1sqJKidvu4tZTKKWv8o8Fnewev/s
14Ku69gTG2viCpOF/4AYXfeiF44ECXhBzsPIeVhWH+nHUsAlxU7e0QSHBNNaWd0BUY7Ev+T1MlYo
Ma9CTudOWyqVSeEAObTKCKBgo+E4WsyRrLrMIE8ovTGpxopI6bMgIobpQVniAMUIvcJD4t7UE68A
VC1EJbyl12BW/KxA487tF0aqDJRJXNgXcLQltbKy3yXDd0/MKyXeqKq3MXeGzrH14kY6Zu6IgN15
Sz8GcZsKCOV2FF4kYEiHjXkDyj85eosMlLi3AcmVkjxcXCqO81qyY3lGCbLGPo0m0UeQvVowo9wM
JxDxgKfYg6NJfDZWns6xBeKqkm7cTkk2P70zHTwdO5Dg8rMYdb1V/QrgffeRQHngs+S3+sVTM9Zx
6gRiqLqyqLg60FQ86jmEn7iDmyfvGWiqvH/SVqiZF8YIwaJccVAn0NhfBrgabCg1DKAB2bKHVYiS
ppc2OFpJWPEQlza+01FiYsM6yMGzmdCVZHW4634LW7S+e4PUM91h4fo6ExYQohNENupr0pg02NzT
XMVin8PZmROiY9fA1T51FvZ7y8GUcb8qPFX8wL7RG7YyE3EBuDozThsQAEmQWFBcqmYMocCQi6IT
iJDeoi2t8DutWY3EEVCyEA2M+Zlhbej8e7IuQwTZo2yj0SD5UA2rs6haT6759ROuWbhprTBiZt1U
rsBROkH0QWwEtls2Aak7GJAOSp2q/PEDYUkO/O/YjCB8yXTdoSZrvTdz76HU0XmZNu3mrMc/2A2Y
Ljij0xahMrDyrEyavQLTa8d45/SkZ1SfM5hfM8g155melSzckNTS2gYuBBumsN55yBJyhM7SEfic
/Mv9BlTB+HkpnQ2PJ7I23wA0vZ7WnvxjxQvAP/oiplu0nCZBt5k43yAKCNkisJCA+x+CVCIKXWwi
7ar2zITtTxpl3obxFni2jzkLf1iopHpksYQFtv70dk9HU5BeYkqi4ggItHQXy+d1odO2nOMwTkHQ
ex+yb/tDZCdLNuyuDYCBNsWoHZ6FfecoPrk9gKmXwLz0+LrBodVtSjCu65u5LFqsNkAO9pxPgiUF
xo2Y+oqNIHBi9i7UJLAmrnrVEafLNNgYP94pr8ga7hpNJXPScC46705lqSPuUvLZnkN3U/j9RYg9
pTokG0NMn/KOMsB3xat3SOXOws+Hq1JSVIEIUEGuQrWjDlmHB+HKyZ76ppppsdE89kFYf90CpTl1
pyNwu66CHM+0EQpfiHlqNqJFNSB7QiNb9KcrERFV91BIctDgAQNqfXIrvkRZqdjH95s5rZbJ+0FZ
SUR6eG04BmqDJWwxdcGji529MyAzlA6TSTTMqwc+c1jgwu6veUbT/QLDFfAjnUIBQkrsc0HdETX0
+qzCx3xvMocuxEo0PDdQgCytvi4MUrMbrgOJoTk6syLy6A9iDyvxbMia+7W3Okq0LafDa75z3yVp
VkMJnW4osr+GKkpUxu3Qkl10bBbHwMx6X8/8+EHKPHY+7XKJkkHEXirwJD0ZIapfN5xBfHaaxSxf
4XhtBPF6T6lnWCKLOqOGFJNBdHd48Po0r4D6gjdOQpGJCB2Qcf6keT36tr+tMmmArj+EfOo+u5OM
OIEua7/szQ3oj82WdtDQ7rtbQs8TkJVQH/w9KhGtKujMuoDotbNyzYuze1XZ+Re6IvOemjw1dLaS
nw5IxOujdYZYJjcTwYg2b/mpstRo1x3yGcZkQTtGQv7Gl44LXKEqLVJCLOTQgfiH4MvEucxb+AxZ
QQDgDpxxRHKrMi48kp5sli04aa55ycHjVp9z0EUigC1YeFGgDVR+k44mgCBxKjPC79p9WozqGd1G
NNa6jiKB2f55nUySweuee2B2t4yr7pIy/3xVeW+2HIQr3R36Fiw6DZGwYfUsavlG3IGOu0wENv/3
+a7OSTcalwHcBLezzZ0WZGGp9cXK3HYxo9E7F64Ea4FfuZsIqb9GVZkgQkX/8Cl3/NclsG+SH/3F
lth0jR3Zihl8bPyTycgKd6IPQyNOamwX8HdTKt0kaFUAXfI8GDYmN4ExDceKVH1ckJ56Fhl3eKQX
Hgio4pRNiKB4OLETq3yrsUCzJjkgsMrORmXKM6CdMg1Clj0UrR9Dks6GSOxr0Kojhy4p+xKIuHn/
ZXz2KBY3dxq5+9+bkIAPsqlohxQQ4YzUA/pISxQ9ZkEj/jd2cEfy4qbdrTrBor3FqeWwWK5Xkfmf
cyoJ7B7q9XiRxRzMycS7KrWWATtk6Xir+wIcsPRMPAp6EvRgVPi0XtbEsgef5oFdLAoLnbkci5V8
axdNymVswL5OK64J64ZKX8hPoxQ4r79P8IFLuNQZ1+eErp/OMMxaxlGPOVMfTn/A992LeOFmzBVc
PYk6O1uxKLkbnVtUv1ZOhabUTqE0xXAfsGeydhHoNq2zHYldflydb4OIVO3nO8mxPvDkN5xSW0rd
OSVb/FU6v6H+Rs+2hObTivT2tQLilNX/z/Eky25ItpvB1SrTocry94ZQta3cGvpj+8MPz9i3OhkN
JbPYeZ07ETb53Gl/wOZdctr4pxPwpOWyAZVd6tA4koJ8OZLRQxAPDnFWMbkCBWbBns+4P1I4plFf
P9rbcVIzaS/OlHxeeAqgYZJbErz0mGRoXBZ1HG5/tOaVfaJpZA4qfHOD36Rg+SqR5zK5/zIAVDRh
Cp93BU2dEYfThhJ+zYxUKyST8/pYwEoYZ8J6WWLNaPWnO8DkvATBU3iRVSKkhukppNVPYS5woPWl
5ypKJurv2CbTlOVaeYfHCVElamkAqkLMPMUCoVdoEiL9HNINvjIOEnKfyWG3XILBiI+D2jBE4aYw
SRe0AZmTg8JASC+9+m4aAx2O5RG0DnjOMoHT9KclnpHpePivBaB0JdgISi7OyuuYKXPXvy9a4E3G
rzFMRnaWveUEymMAm8pTjEJ8tCZOGevmaHsLibVx98ibmcc/+zN6P7pQklUCQqHDlc6fR7l7bpZo
1ZWIS43lgKTYxfF03Nsbm0HqqWNkJ6chb5YV2A8UwqbGOOtu6z6s12EJ+N6YO1nIfQTkrK/XNeX1
jmRKSjW3W+lELqrfG17XzT++IG5z+jRosCMMv+tElZlpUFoN1GupuxK4QslJBxF8c8raB/RQcxvv
fZOzYKrDmBZe7s+AFeM0+DL8iwYVuV+h5ZtWQ4qYRMycQBgNyFyTq6JQyPS3A+WCytpHNokfL4Ig
u1I02UwzsEN6OV/rAe4VG1b3VRsCfB+LRCREo8dUFQ+txDyZjvUqVOi2v519vi+E6toHaw1wfppI
3eOkFTm3R6/q+crfGFUXqTsC8Z31HvSPfMIbR9RjnAE+169oX5LrCpi8HRHnbA1By9kuT2lI7uLg
H4otJw/SQG5itEn8bfWzgLHpFY/Z+y8vBK7gY+x+KXHktkNiGfHbEQ+BuceBfGXlcfunbfQzKfBj
eMRI06pG6iEiRqELANd8UKsl0vVoACY9Q5zTQn33FIIwBZYSOwx4w9YWkf3xKcAhRgPYlE1TQQn2
Oo2cIe/ZPNlNDAiauZLzKhYXM7L+C5DI5Ha8dgYLsgTb6JkaPUd4U2xfUH4oG6bNWwfjqZtoXfj9
b3UXe1O5Ht6Ji3PgVhdJ5z45HA1DxrEXCRrBRaz1stww4RuGVmE8LskVIYNDQKY+tNACdZPUBjKx
YX7mTinZlSTr7tFxfHsT6Is18rZVAqW3Rdl6yQtBtbaOg06UiJ3X7gIo6pukzbv6OFCrVOyQFTVn
P3vbrOkHTmx80bUyh39gVOnnCC9lxfTf7PIOOqAO9utNrg0z4sxsQ23lajRjc6W7CMoNOtdT0cmA
Ou6GNbHMjasghn/oepnAfNaqO5FN202eu3XfJuzJS63RGxY/YO0g4C1oZiT4h3/kZFOgSz+7xnEb
KHAEqkl/2/TuAu16umhtYPwIuY9zo7einP2UjBi2Ii5iuwdpo0h1JOcZgSLrWJdr69fnMS7SNg2B
F8yDK48jSqY9WcDedHfssa7vhBP16tT9sLmut3E1UPFomLmLGz7/4R/r9f4ZqOKBoE083bSHwG3d
VXrwgimOA+U0ewFM63hXrhaoseOaYI0qD5rHHAw9vrAW6lC/fQg1VnlkIK8cjkX78/Dx74k8KCGm
b+XtG2lckJUrFKj1uBHcOTT8nSAu0FHxVJtFivOvyeHZ6hFnOIbRx0hxitmm/qgRZRxrRlEp3GJZ
jGw15ZsGZpz2tSKnEGtKZlZ+XqrzM3Lv3FUmlKO4TgUvZJgF0t5mv1e28tLYv6TzGnfOFjwX8DWw
BYvdt3wfsywTDHgY6svMzoxH+//txo9MVHR8Nsqf2qHEQWAIeVbCAzmm5vDvsjrLYwSW689l0UPI
RgSKj4NiBj6rR2i1WEH4enH+UvXAhIHa/zbFAeRl7eD/mPcgTEC6/g+Ls0onxnIead7PQtbtQkQu
wwnEvkBJudr3gIbnvKHCUHI0ehXZZAwdGI5psT9ARQyEYznJrF5infHPiAD4oIm4XvDiMxTtNx5M
G4XQkqdmIDp01Addcxj6Wb3xBqwLgW+lI8qSDMRZU4sAmzBGJCtDE1XHdbo1bi+dqyCXXOLCkBO9
S966XIotLMEdPxtsH+efGrXLgwchwwbd37ir50vOuMO0EEkl+CfxWFpII6HPz/4KOIljdKF1ber2
UzycV/rC5s4eqPG7f9kXu7UlYpBPBwXMCjz+GLMulsHklTFTqdAIySheGE1GcaJwN/efEXY+/BDG
45fMwzsualfzLohF1AnDFNjpD3lTpfXc6nytXAfMZ7zF+EZDrNoc8o1Zc2dxP217ejgoVmUSqbo8
oYCSscQJIsC1Veboy0ygYSiu9YXDngWX9z7j56meGrLiI5Y3fd1MvYY7r6f/7j5agr3aRzylOqYL
axZfPm8ADiCVY/8TkVpYDh5FiaDR8GKwr1NZq4dhd+9Y7IIu4qcNDB0zU0nqCmBOM+f3f23DCBkq
M3gwhLJrtl6hb/cgph/hhfrtMhbG7b5djuPrcxPd5ocWd+gis7gJ5YBV+Y5YtgGndIAr5Ru8I9GE
U5327u7Ku+rJJXPWEvGzTOZilQZG+pwIy0UdiL64G+Awl5cqGGratw0HBVpNWZTiplgv+gLN2ny5
lv4ojxjmy9FkrJMrV8Ct2d7U4YLf/KkqhVXxBtSnM1C+CJNzcgpgn+7e2N2wupld8jyL6v0aMB62
D3mFQxPczAH6XmorzqCny2CYQ2z/ijOhs/BJ+xsFMoiC7ZleFo3jCW+DhVR60vrD4aGVbyGkHuVC
3/lZEN8fYgV8UCEvhuRPix3ffF8nmDPeg7HEC1Dmay/WgMEvLRnFcShszyzQlOcU3fm4G0qYuMUI
M+zLwZ3DbMpqQX3iBKHvSe+Ei1cjSE/cAv7PuOvJDFD9uxiyvd53lsT3/1+H0CPRam7OhSzyFZmx
VVvRe3lHNSZl2Mgy81FRGmKq7r8nymfn24zbbFKw+dd96zrI7gRLUHdix/APo/ub5gQYC/PXt/Eu
ZX0BE7CEenDR29+Q9pUwxIZkszOj/5R4MrpkgbdmiEaCHyfo30f/ToyVQm15j6BCmb0lapsXB4MG
xju0CKZajvBbp/02+Yeam4eaLcHG2bjnQ5WaVgUctGpzKzR06GoHzvDf760tlwcRlQ3kcKT9VAD7
x2eaqfYdYRDw6Vsj3zrMd1ihkC1t4HYeHhyaRW1Qk66OatLxJi3C0zc6QSkmb4TevbUaKhjnwbMW
J8vki4fhW6A+/q9sg6M3HrRLRnPLok2LynjlI6jyRV6qWOauotecW7hlVHhznxjQe60c0IlcY8nA
R51Hb+9d9MIrd0uFGNhnKT+k83Ra0+sPZSzyyzj3m5OAhkDPuScnq9VP/GgQDpifIbI4QPRZUIeK
qlu/NwoYghtp8bcVdluHRSfWAMcdQNEte+F4SB6/qtFMgRqRbphzHkgPdxFLbod60HSfwWQloFwA
vdobdqdaI+S807SwnGsHGcJzFRdwVSTEhpOgi0yYSEeCiyWknXAbYALcdSxxt6o3qSwyfZI68xbx
uYLEAB7vY7wuV2pw//C4pQkwqF65Oa4DUmrNy8ZzOKMaddeEhTZhGC5KrizJhPmrL4lrcTeruZYg
Qfe1clvunILIxuNZAC7uXG80nt3rq4zI5OTwqPA9B0AHSZ+BmbSrYnqqjruSkGlU0LIHscv9YSTP
vjPqiM72ECtNLjdDwLgq2nJd3N4coTCv8L2KYIF0ZboMgWv4GsIIL9WHO+X/Nlxj/u2p0nXcQwJ4
E2d2Gb6dknY7A6wHME7sPKgkO33RY3X8Bbcuh4px/L9qOQt89z8pH4TJ7VSVLUpDZNvfluBOSShc
r4v9RBlMAA/ZV4WYGXb1MTf2mOG6kxuLutIvHmsQfuIKZgIi9608ZE5a/a/2qPV6eFR0zKQw3QHa
gyx3Nxt7tnZxeSZ31dS8yr2I9wJi6HBTV1U8atXAAFaGzs4tb7132DBiVnMiGPMcPQ9BwWIBTybY
BbcJgsTIEe6UHAMBQLezpNYhEomrti3I5ljMkWhR/qdG1xsLIpMObr2Hhagf5Q8Jjg+Z+vAbRhhR
adIQKQmuslT2eUdyPu9mOVA5z380hC2he7i97QCRhHEB57BJjwQOtRvPHU8+ZoUC9cCYsIw8tPLQ
CiunolTqt+tN1FAXFQ+XKR1nkYDj569pzAaIDF2abuYGxAgq3+M7XJPAExFDs73cRkE+g8AE672x
WU4aOTn9/aYFlRb1kL8kLcHfbkKt3sjSXGNUv05r6MwXBCVS5rvqgzCmSaeInYfIPXwlGdfNV7Ak
UyRcOjLilZclq7nuGyoumj/e1ehIW3eWiKrf+0gOX92fkJICZKTtbq4L7TruYS2/sv91FD3t5FZa
xGd+ZXyHDXaj7bAIZTtPO4bLOOG6q+RwBM6TvYOJ4Rl19RrOebbSKgNQyJJYPyohtILsTwovfG29
xAvOp2Y9Phlo8bzoBa1q/u9LmaXimORbqt0xzI3MyDT2CyvKDnuASaenflLv8wOAJY76A1/d9V8/
UzV9uJGy9akWn4NNsBEOyYavEziEORe0h1duz9hbfR5P41hdlXMZijzwz5yZoCtmG7eiYzntj5po
0XhimF6Pj/Vu3F3IGFdjnz10eCmvtLtkxk7ETMxJMCqBSsLNDs/6VW8zaOsL5ncI2xCgq/onkitf
y7+4NCZYTsOm1UPO9+4XzWxNRvxCZT0UkmeRSfFGm9Q5POAXD6gzWkRwVVAOJjJJnv5Kdmr2ZJa4
Y0sNeKw1w3mDWCsI3AhGJrypEPwTx/3JP+ioJzggsc2WugiNiidAP7Z0Dy6s6KqBxXr5Hq9HV1NY
W8/K2xelD8CZ3RxhdsNrjtt0Zt+0RiMTPRO09w+hahUICZpHL4wiVrtvXcBDhmRIzgo8YhGXyd2b
Kq3CzOG26trBEVEiTgRu7b/4XxKPu0jd0ORFTzd1HxK16JmVzV6zN88SuBtsqHqnbV6hw0T3zlLE
1C0J+Pz9LeyIoG2RRr+b2TP//0C/hONrtQZXIT7RFXAnBDWFzAe34zXSVc0/ef0GBVeuUyKV0r25
ECWuX1czOHoqcp0I27xGV6yCF4VN4oMym2Vf2eXErc6B8hWjFiSRILUh9REPJwbJmA65u45baDJ+
7dg3isarsRc2y5PErsBQMci5HYa6/fpBni2aANyQJjUBjpYGrAWfuMmdSDh+Lx2I6nbhfWUKeUVw
T4NKqL01QSGq4fBmOV/KHLFXLuNCrt4RNL9igTH6vJqXv7qGYOwUAzRzs17uE+OFtsiiiQNY/rol
wH6CYMIupsCBEe1Z1epRMZHBJ1NEjRoXP6nU6gZm4aWvphRsRw2d7+ulkKdfbuHXaiP4DLIniCla
F4eJkv8MoyLDEQKeQHpnhrcB4AZ1MgwYc2OY4WLFi+Sffb3257GBXtRAfLjd1ruPogccb5JRraKz
t6yb1Tf/y6Vqf5ojRtG/KHYxRX7iHAyzEjUh6LsUcwJKvpsCS3ukKOUW/m7vVH8PqPJ2U7ueRrpD
0pmueyGyWxQaYyCtltgmVnzVn+l6KU1ZKTOSplYQSaq6dVSPFTM78w62DYhz566f4P4C+2wqCg7V
b2IDES5TBmghZyI7Z9+k/io87sEUSItrxf/QWZIMUuzY1MYFbvQUZ4W+uy8tpiGM/7sqj3RGUYc5
5P7cr4ZJpsKboUYJEANcEEN7qDYP6VYV3bP3XTG3L5mm6xNtTtNH69f84UchP6F06R1R/jIhzSk5
1rjirc9xHcjN05vt3Rb7sD7i8avBOHStwv69DLZ5PQDsDgmT5MA0KPDVtbkuisIqEuiN3ZTFBb+c
YOYQ0U+iOJstYhIwFdFr4iy3vMIclXHvoM16LEfUmvQt2sUXFxjeum2dXffIFfJCYFok7J8N6BK6
Dw5ZZUdiZlz4y/PvJVICDfx0e2IJZty+9PLPe3pFTbQTcgWvBFRsM1rARztUqJEhzUT+1Mw+YWSg
aPuwPjibycw1NX2AzBWY7bTogFIzhpYas6KiCi8IDfHpnCtIkLRVasqOnamwCIAubFwR6sPxJLDH
SW6YtMllNxhQReWL58OcB9IN/j5hqCpZ46wZD+rRpkVBInvn1QZ9bpsVKGwYnwcsO6ft1jqJ2ayG
oV+p9mnbwf32khOuXOVCJ6yk9NlG89lGWOHVFICkcxlxWscM3TRmS4zlcDuh+HbTFM7B5zeL4yPu
fo6CorvKaJBjstQJ7sFxTqHY6VoH/C2TspyiFjLsDsrv1saZL1D5zeB49pm7wzSjHLUKns76nPVk
l9yEW/mAU7rgO7TFZrhsy0ONxDoo84WNmOAtNf7Y8rDHfag8gnl9K6TY6DI6oULfUcrH6qeAfvL3
/f/Pw/VmRc0dsMQpSnE2rZRTxRD/FVNVhfEffTeHYGuU8eGZp4yXiWwJhwPzDOXk+9S9IaUw8G1y
lW6GROwVFD6XLhF31bLegz1sLLmDS/m6i+jk5E837CTxjQ193W7gke2isbiRLNalIsdxX02e9nH4
wdcWDUGYnv0W/gk8onz3RuzVlI0NBiY+Zftn2fSMr5XO/lH7MVtgy8J4IdroRMIdWdbvBLIp26VO
TsviWPl6yj6dMtCrvulDUD0VT/xrvw7rO6IArzCk/BcLkQBQ16i92KLnVUd7/IpRFaJU/nb9b5zR
xYy+3qz95U8Z9Tf0u79ZFGa+PDgZlP42FsDQ2ncK6QGguloh/i4Oq8nYJ//HAhFXT1Kx7wY9/22A
mibRwEpuDlZEuzWzPWrGn/sFY1yB3qaQIqv3GeEMfZ7tanu5/FE4AHSmt5dRS9vjVldal17oozlY
RnF1TCuTqIuPuiZi6t4dLN2eQ1S3Murt1adm2vdknDO0A6koMUHV7DY4PTIf3a2a9qoWwh8DF8h5
208s6tGBMOhh0HbYh5eIeLokzKRjiVEq0bWEgV53MHGWtr+PWLiyeJew/TQl6CjloY5KRLPsVsAX
j5zBGq1K8cu4j46mNK0ODI1y6ejlrUqtbPy0uMNPOdCelqJgqw6EAhRCcHv4Q1eze0sAeuJM3jZ0
ncW+iMMYpzKHRJpATYoWm1ubH1iViS1dfQOtlvGZGekrmhwpjdBfEjJThexFTUQGQDhrZG6POlci
n/mpCgjmn0awaaETYlXiWWW4DFE3JtysKON23ukdncgYoRf0kqHZKZXlbIYfjMmrBekncJlhOYyP
Kn6fQNcfWSGpGaHhU2a9AM+4MKy0mlcd3sUHW4ZPy5kXfrRAvOb7N3lwLkYe2+usLiGa0baiwXn8
f1EjSgBUuxBnSg/GiRWCxifpkG/7gZy/Ck7sD0Iyvcx6VGCWe4TU/Rt8hCKY2ViHgfHvMxA8Espw
VuW/Jsff3pvQONkrgrhs/43VnBxQMJl1s6vfEqsPA7NZ3W6t2Oi/71cE+tMUh3Ikbneqc4mlK+x1
WXAvo0uLgx1NxprkxahmkQ0vPBZH7UcxvgO807QwaIlUkltzoieE9yxAQr+r+2Q0a+0RQpDnNcZT
paOxWAlMcJ6Uj237k2AWh7x6pW1R2IaLcobQVhflD87xO5RWQ6jyiUMoCpxCJxnmEi0zaxx2ESRo
XhaLxidmvO0bJq7FRgcITIbE3mJJng2SSVTnKgJ3PiZsybJxizN0SY5v9uEhi0YTJpcBax0jEJ35
02KabrtavU2WtTxaLjzR9Ud9p9FsaGEij8+F4RApFfd2b6IFjR7/25iNDf9gZDorcKtbHzscWN5U
BGvqYWVWkJ4C3rjNK4QG/0IJTNYN4aiuBXnR/5ERQ7UGdp83UXYUS9kWYN43FzyD0I5XuO2vh9/s
UZ0g49yS2MXUHPTIxyyBMjTLh4mcfIq8eAnJz+M2N2E9IbhsW3AtVamlC7fYWnIjMIWe2gWbDBtV
BbuOibz93W1Ic7spv4bISbporGO4tPGYdZJmYrMI+LfczzxKHYksNIAnqNpk5JU82GWH4GSMrd0N
rjLRDj39+LsHN3rSN+QsFwUGQrNcq7ifowcFjIXiQW9k/W9XTlGGI+8YZaWwvKcKppAafKx3pAhZ
0sRlfOiuK1CHNtKRWIWJc5hV0rCNajgJoOzVhCcv+uF6dxTEwHL9H5Big0/K7ViWYnXmI2Hs9PbU
Ws8R7AiXjsEtEKB4PDczaoYEJV5+aak3rDv95wJLNHHPbwGerrfBs3oO2rswuvJcsyGd1Zhi1hft
CmVo/Nxf9i+QhlaDwz768EKeMCsTxHBjd5Jya80Z8gP9vqsRkmKSsSlax5ufFhHZ2wVWLd5Owakg
XgwUByxLdtus1fFqXrCfGOKIBCPk4ZJrmsAhTFZlsG6x8kJQOW/UZC9LdjS2P0a5Y68AnpI99MbD
RsohAmVkCCQUXw6Bd29hgAtKacGPkXAXzcV6hPiv2pGFMHX0FlkJcn5anlIDbfu4O7PEwC46I155
lofNa7Y1EwnrHTRNRSYWluQDlY40MGfOrOrzyBpHhMRHu1TbR3PMHusco8TsWF+NdS64qczdXj5f
ONWKIInYpH5DcZmw7X0Cab//qCcWH/ikEDPJ9CKHMdA8LjnwPNPVTIQOOtNDFo+eIjX0z5rjp59k
1IdZGzgcJdEg21+9wNAh36Pk55/0h6NU3ykvuRGqZkrYs/6RuqPvx5Y32ipNxcjxmR+gKsMVjdFA
Q9jXEQyHg82E9DzguHSPOSTL4XfZhZ3629yh3moQbca+TAlMhH6jGxHKxLpX6np9n2ZfUqxclEjh
hYg6YWseLsFRXgLhX1MpI+gLp8JI23OiRLbtY8Dtke6VzoTam4KKXCSabfakfdqRkfAOQE+a8hbp
ms7uypP/W7WuMiAe4N38RKjODK3y1lO0n4Jw7VwpmsD329Qs5mxEE/cFSMfcYgtJnmqElNKC7fpM
xiIT5IrBPo/rmJvfchZpE7GfuRLfzj7MDCAveSBIiOQNm+HSs7Nes/GsZqnUWiOaEQoC4x0W/2zV
Z5wpjtVlIzg3Z63kAXXitoVvzoP2wnZDtDZrTDeWe4n5D7+m7ZAHd3nSxQudhL5jfgEdTdRrsxrJ
T6HDPxSAATqRaSFeildlUeDjgPbZZLTZpoHcNW4hbp0W6b5cbDcI3nOOHYf5oiYTCRUwJ8iV7ydT
HkwNInMS3EVFBb2OfAe+HRhkuWArk1TxiI4dY4tEjwsePOYjCc3bYUksuJzeGhARTJHAQm7y3KV4
VeJ70Y6Fw6VUuR9VArJS3/zBqGFYiz0UIwSrghsWARr7OEiA2H4DAn2v/LbqDcuOnnnnElahz7yx
BP5hg9DLUMwnvPKkvSNKw868WafX8756ciRik2QdL5MaqNmS8cnCNrmPiVc8WtxKoSaP2MSkDEfq
b+sJOIKMlNmFurU5iDw/chgwF0eSHylB7jKJMngNNzlMp8G16AhoO1iYnWqVTTIFDOexMjOC0Vgd
nWxVquSc1/KDk8qgToAaiL0Gk/KivbDxcCYEgtKTgv9rlr0FyidsDyYL0TugP8SX790NGqe8/h/0
MBHGSMPpibTkIJbBJ21+FYOiZaeYpr1GtI7oBR1730kynE2ftytIq4s+J9N2QgoLVcli80HToAlK
D5iIlzOt5mPdbAj8je1g9eOLxsnXQHbLdlUf3lQDyuNUo1LEwtqDzf03lnmzLcoIpBGM/Z35TIZ4
bOBqLbvTR+TnIJxqS4YxRIY1qfr/bnfiiOEc4esOmVAxQE6iS2VsZr8UP+XcuIum24XY9TP2JmiV
rSi4dJD3d9Yfyv2gQLQGJxHTeDvSo/OqIo+hPrdyFdlDWVM619YeYF707tEdGQnEyouFf0Ob4sID
76yumliVRXmZBi8kwMo4iel64TIoe0H7z9zXE/65mUf5qI7CIeg5dLcvhID+Spa+wBuU1W7MCiNk
Qe/RcbxoZXl5ysizacu+o+tmnNX9Ukk+A82VyeM3L6Xvtm4/4oUa2PTXuhKUYbb6kdU2I5DEHuRo
DUO9IUFxGjHjlHCxyIMoUKgZkWHii6qJ9pKgUAGKWnWQTJdebQGsSAX/o6RWU/9VhAolJ1RSkc39
8Qt3Y//IbuRcIbDfgfl5GKuzeaOiWbBfjsrPZo7lFwjvhWIPxDevLXW8e/4nLFUr8rMeit4YQoIR
yKE2RAJHlVWCgTdVFYtvSYawBNqsuqlricP2j+6e4OH0nBQMM9WHnv9rb5dtUwy6JLkrRQ4FtIFJ
nugci3ayxVIkogzC3m+vTfAXWrp+3VXvte+OtkhJSMO4RqcDvfneGjUcfi5/zJsKfxXwFDR12+uq
4PFA3LfL64XPP7/UY3XlF5qoL2GJbtK3j+D29/jTFCXZex4ZpjdTwkZOKqTSKIJj7lEk1G+NX60p
x5LCjy7Sf2ZOa2611Fwgz+FhCpnLIunOCiOjeXju6eBbi2nEgG3iEm9Nq/s2U74UnCbaIyvO5zNm
q9zyWdECxF4iOy+m5r+DuBp5ZpTpD1PHduPMqzMjpkHHED5aIlE5hIy9Kjxu7X1/5WEosTmIE0oM
fRCGCNyN5JAl1SBMsLH62XaLw5J1hUggT/gX0H1UA/EfLmaPMaujYkP28SEIf8J0kuLQuxB7xLNC
Dw2K4NDzYwKV5Q6htiVTspBjAIsAvYZAdqndf5fk5Z9fmQnlDPOPwJpJr97otGlku96A2TQWLe9z
/+Mx10XmoQxCG46ZIzdo/CzqeA+jJ6qROAubgAP5+5FIsARQ7T8owwEXU8f0YwzmD9s/yslSt1oD
H9um6RcdeBaLCr7fxlF9nfveuR0jYv+VcnWH2uGutZjr2rBxW6FbCobFdAFw2SJBcGNPmiBTiJrs
IheODErDaDPnpWaOpTn0WAm95POiWvdmD4pK3CXEdQYRoeJh+AUeKpjOSwycb4egOcr00vdm4oCL
P5JKcuQ4RDF/m1gqwm93nWoFwMXSi2aS+BqR5rfVIWIrQiS5KqNLV5gis3B4lOLh2EeTsnn4vBUo
gtOa+vXbNfFYXOXSmr1BVdJUhUvbHBRvi7tRCFJVf02mL0BrkTLIhdeDRPmjGlbjucrXbIFWntk6
gmir0dco2OSLIIHFRQgoAor+fbHL3dTphUCD+/zLlUxHt1hehD6Ub8nwCOnaDZqVQ6tOzp3EyYi7
04elibFrZuK70tdw0bXscdY3WylwZIWenpZF4BeqmM2r/qI7ccDuHp+MPyk1cXozb1VRlTvR2r4W
c3sdrFOQon8LD5L6BKk24SzOrEQEVdeSKhXW8G9rsuvJKuWy4oGHzDW4kW2n4PzMDSDblRzI6zxL
Lq8MGBpnHr+B912wOBTmpLwbLYWEsQYe6cb++6XELIq9xn5thooSAxgHzqSHa70KfOMS4O1rgb1q
XihNNJRfDDYvEnpq4QhZVdAOmnltfzQqSWNLW1xC+ra+qYWaEkgevjDtIc0riJdMBrJ9pC692eqi
9zqKeKxhKLZLm6rlraQOGWs3pjQrowZxMr117kYyl8h/UlJNuPtEZpznyy3vy4PmSZaodIH3fHXn
Q1BGWAHl+vYuy8cxyLgD2BHnYj+drLI62ADG4jiwPNF4Bby77qSZAGKEAlPwk99++cpBFOutKrf2
7rto/277s4LLxctisuE6HeTd5uwGZU1gRtole7V887nzboobwmt3pgRD5Cslzkv9FmgFeWlcBaYm
G9wL0swDmG59h/oPEtP0p8igC2nBZe1bkJfC4h1mqSZf8LKYTuuBKL1ffdcYfNmuCyM8SqXuhJFh
Oft5Nxzs5IcM2eMxe3qjTtaODvGHoSd1L7N8uWwn9fID3DeS5LD8998aJOem+jB8257AKY6Tk3GS
VqZ8YHvHVTRZK09EGRYDNo2I9Z6qdD1bmoQ3mGsPonqPq42wRYNvvdgsfmllI+MS4wblg3Tmali9
yQg6iUT12QyTNuJ6nN6rElNpAoijmARFDkermTW/pU5xb/iOBNnXtqyzlnr7NCQGZhRWNU72eyEc
U6insQc39VWdA2xQMNyJ9v5v6DoTAGVOXPBwNDyW5fCDi3C18OTyF+nwU+n9wJAFf9jyGSdw7yvM
eLpDg5WgJ9kpasQpE4OgYcJ24XaQkSawv5HXwQY4cOETn50JooDNkI1YShmGiZLq93dnZmRQI4ZD
oMdXJf8sk4wfwPEbnAbQnCdsyQF6g8MpRmUA2WsCnB8UgmzhQybxh64/lzzdW+s59z/M9jbStOUy
huXtjM9eR4l4RNPT7vvKrQE+bxZPQOSvMl4nbdy/3r7qn8kNaKRLPNZJFE10TIqRdTA1ylLdxr0K
jpJuaJx7Es+k/5LQQd6J29jhjLGKmbBn8Ju/y6swGFdrIXp+mdnKmIRF4K50+CPoJ9wQpJz0cITd
BU+aXJhsrw8N8laWCWLH5o6RViaYKxW5uIUoMdm0ff3/UkuSu40ZzRSdvlOUoyBlpr8Sb4G3V5hk
9kYeHegUkViBKCnIFMt+hWiF/8ked3704SZxJUWsjG9jJxwAkyzRkgZFID0uP/1r9kJHZ29gMgAO
0ytX7/L/CtCCcAAscpst7k+MvPukm1Ap9QAlBPxp5V3J6bBY8lrH6dghgahZG/HyMt9xCBUNe9T/
NjmFG9GawwpF1XYodTxv1UlB63IvCVw1t2+ue+vTzOHwP5gsl2S1ehAW+MnkUD4wfvHsuj8S+Y9p
EVF5GTXsiCncl+1mb/f2C8MYTtceErGL2nIbD2MYuiKI09WB7cxIfTeReF6GAkvSZOy1t7lzZuIg
ERdaTlUL6TVCxVZHYk1Z2V+u8FS0ibEpEljw9wBBUsLWms9fMO/UhljnSN6KAgXL2oYrSOVpAp/R
hdkVPncV74VSMtESYAdFlUAAYHZyZsslSn9ZaFPbfKLbgJVmUnRMMUgWmQjV/MN7KG1Q3MWU20pR
1XdfXeT2ygRlzaW08s2dq3zh2lYgoiSeMpEVCPPcs1EUJYuLQHgCC/NOBjB346+6oD/Cd/kzZTxq
EqT/fHucZK3mzyE4R+gXFabNhw0SSbe+4lF0RXMQ4a0KRVCykYQ4Xj1V1KTl70ZxYsLHBbj1i3Wk
ENswrYAU+cxYYvMG+eUyCCxLr74ukwy3X6GzR5JwjmpIlxjfG8kYgNjNvuHxs+0GQxZ48XBvSNZ7
2uneN4FQtODDCxKGGHcVWSMA0P7xGhxD395dy/gfiiGsMRC0heI54cH7vHwhVOTa8gxlMcWBjmxz
Li2miMylQjaR7h0ewoM5LNYuAZv2pKzdWqPElhnMw6L8I41ecme13CQMBss0C72/o09Wn5bkkqjG
yLsU7/tjYXJztZNB9NPxRUlGLOjbhWEc3XLGphRkQkFcV2cvlu2sGopEh7cOZyrfORuNoTb+rH8D
ilDRISPZpBq5HjgUEXWsnmrr5F+qEmgGZ4YsVBWGp2oH+DOfx3HSVRswe6akdBxyWAK+W66Yk1d1
hyD5jygxJDLm6lH4M3Dt5s6pPTkKIn85DVS07bVZgEy+rzjKrrlZDYKU2kkO2FDqF0sm3NQVpQXU
bw1zXqJJgf/SLiwINhsW5Mm7mV09hal02A9sSkf28NLryhIGX8V7ZOxh1ItO18ohtnljPg5o68cQ
mQB8eOC6W88FzJ78Ia6+1Ez4rHAXc4Vr45LKpdRZPMT1zn0wBHY7ZK9+HaV5UeO5FmOKTrH3/fAf
OX0cNZojOa1hyI/1uV4NOsp/tJyxkf2kjn3hQzXlRZjygy9RXB0RYLKyDoaw7Y7Dr3ktw1qvuUKS
jqzjS+EcdTTCgTK9sZtCyroECQ4EJPLzObU1TfLPCNhxaAQdoEviShh79vkKc47qI+J9byfnfku0
WTVwg3r2iDPX1EyrPSjUy2F+x/UyOPt2k8IFlgxCXLdtLX2QVc9q61/aG6+fJo9RMd3e9L1/y5lc
OY4VMKYWaxj5WGYX5hBoWjaSpIu6M8+kIH58bGXcJdgfO33JftHCldHrRm/KQyCI6b2rO07h7Fzh
qyqZwTcg7H9c2W5kCgtwFTTcjAO0IkP9o/jVp+6/rcnEXcIAII/rcRPrLaFIUfwzbCAWXUd1idb0
AYNuyZlSVv5MxYGZYKHVV5+yk9QYDecxNG23wNIewdVcMNjgskKP1hQPIukaDsmE1v+LP1Shd1Qj
xwqiXUNveMa/wWH86m3bCDVonbCuRkHLPckDutv5Jx1wD4mt4rhhwkkspSAfvNokscaA+P3jL2hW
cTrcTl0lQ4n1TFU1gKC4NJw/+E/nyJuiUM3dZJnOTkkUKyDNadqgDcgflQt6pJ/BlhnDfbfn97HQ
Ga3Hw9tOl8BFmqXAQXW23bBMOEhyaBDDGlQXsyCCz2mH15zTC4Bhx8EUI8+OZGIu0je13aos8wWu
ydMtyJSY96MQSNeJgCqlFl1SmZii9dC9NtzXFgTg/Br1EmpXCEeFsanHU3ky3JDIA9+ksbBm08MR
ikuvE9mJXY4WUV8mKXioiukJAh8d98mfEmtbOOmCxRqc2u0W3j9DNC+7XEUISceVdAAARJ+kTHei
IhZF/tVU24XQis27qvE95KKXvLUR5/UAOFwtMFUPx2+fxMZ+rOFI3n2WPr1JfYqSqpPTaClspXPt
Y7BxW6ToDyu07oOEfjsYCqUUpc/zJYy6GmB/Bieln1Ar0U9+zp30RbvPOsxk8l6tuq6PAknvkMNL
HcNiz1ffaZgEZMrNxz6MDlM97vuh6gmoiP4UZEy/LBn2tMlgzE42TxVPMwcNEaGlmV9wfE95DCs6
ngSGjMCZiXw8Uhq9cqmX/HpofT/bajiQCDAlhdDM2bS9pZp41m5BISQpu6l/rdxMwzJIwgX5tffM
gj2Dh3k/bNUvWRZEZdGsCHhBYAfFErxYECuuGtSVS917IXhp/byetVpr2FtqC2ucy74mJ7z0WYub
9QE51jAS9VivNEVTa3yZVM0gvVpQYVlmSE6Qb2R0+I8Dfe7cekI5A9FsmQOz+x3OdtsEXUMpfw7F
VUEuLvRAO9fKUe+XFMtX8DYVrW5zMXD2FlYGWrQLSEh8GTbT4fPaE7FTRcUyUl5adGQQg0nLK+zM
ktoKoCoQJH3+cA1cbQpt786H66yXhlWTmGGcZoM7/uXfMMrPF+wiGnUdhuZGN+vIqzJvreoSkvjS
zPwzwZafpgOycNeeR1oVgz0Hw+OfTUz8ZXO9kETK6Vr+b0nVbItFrur3kwYKFE14qlr+9pVQyRKf
6fFuNsXUJmnG+7PE1OQX2yBMGZVAFCIteKweG2YCrRFjBFB7CLj+m/+Zmo9YshV303GybwrdGFfj
/WyJKIix11325GK+z6G7DLPZAcbesDS2ny+s6YyWt6AQ7VipvFnjI/ADZt+xZLQ1DxnHPy8sgCc2
5SLxsO9Ha7xWetugqhWHJ+ClVSQUaqraW1WiwfiU800GO1dZK63hd1ugyjR/NYCn18tcN4ShPM79
jBoV7p6bV3ertXzASpx65oikW7MXV7SrQUfaPcuYfinClfpOZho5+no3uhx4jd9E027w4rXNYxjQ
T/wC/Y6Gz6iDk1/eZfAVmXksULJFjVZpR1OZeHY/w17JXCXcjJc0GQ0q4U3Rq/NIbH6b4l5wBHXn
cTdHkz92LhNwaRk6SNZrnfoUmb1ZUMyOVZp/xJve8vsa7DHUOgNKSI38lfV+Gw6RkUNeHHukrKMx
pVd4J+qOeFYl9rJQUxLcRIdzZwe8O8KQ6CdBWhxUEV3nkkZ8kEe5JPKy1pU7bC2oiL5sZ4XafIbo
OViAKtRiW0sMQgPLroLqw1u8UTgSjVLxdRzKZ1XmumnMU2IHoBA6N3kVqy+1uE3oVNQv/UDQ1397
S+/LaORkTLrH2HPYK1HWXxEwyjikGxleao4EfjM/oH7Z9Qbmu/sDLCBrZ0kO8qg/KXxW914WYJqB
Ag+2Ik6PQDIxNJlY0WkmGWqxdsP9P0jdkh7JZBSfrbh9qV3x0zpFwWelZiQm7IBrWodT3txkzL3f
Asvtizo3OMMhrjwHd94qWzfV8IrIm6570DZPRCBsDhcwy8u8Sh0deUVUkcI9zUMJa3j93hKEY8rZ
2HAY0Sn3C3JkQDlm4LdL24Rv5CnG9NePwvJYFilV/Yl+lzsV+WZBBesCxgatuATWfEKmR4zjEKal
5xEpGDi+nnndcz8WvPI9WsaTZYRfRMAF78B/IdVpEAInpzKHe3RVNTEMywvfH9s5NmBG+X48nZTF
nG4bWwJieOkU53UA2sRej6oaHLoONq8TEqNhxvDJEClFoG50ldMOxhY9kdRGxKKK42yYbDPR9Oae
HLOU+EJG2YUPDNo8CnU36kogiwMximDBXP98IM2CMp5hNIWJQnwnGWAwOnAh5HqtAB19F1aK9f6r
FEgkExCBr/hEH+D/NyiPa+Htl5xxhLObuRygdUrZivCE8FSmGDkvQC4SimzPpgGWSR648Xn1SHN9
qtiiZVVpGKCy7L8ZuXK5Nne+AxFnjQDAiFYZ3JSzWpBMCt9Cih29rzcJM3UoQMFOEyVFgEB+PYcw
UGMAFc5IINapMGE5oDHJ83pSq/N7sr2Ev0VkXeNOXnW5+CNe7ZghXsYrWahdaBIK6pLiHXau7iNl
XnHnuvBsn9ZhYhCVBveE7wChoYRyZo4/kGJC+XG3o0W6uYdsxWV3nNI9tpS5PEnZ+T958S9AXJRk
rcD+zZ4Q+VlHOWoaOG5uApc2urg0peItEUD8paKGeIUhkN8XZF8jMYLSt10D3ZgcZY1NZR4+Mis3
2MxwKRbAN0REZGl3M74wNwlF5609Cj30fHOtlMDbmd0b6fSgJh9ggzgzwXypJ6P1q7vtMxKwdbAg
5SSSw8dtESYEKtiSpP8g4SJw5zfBQVFL1lCo+P6eTGEVF6K4DIvc/rdLzuD2TTuW7uDxfYeRdu/p
t8gdvm2M3CTMGh8i5iXCJP4bZ8wV5SL3ZI2qbENu7gedk4a8+va5OS8lJFMT1V6KC0l4XBno15DL
yQd1dY+FqGo/s9GR322jOZPCMh1vM3D67x+418MZYKOizGXi5QuFmrzx8HpQ9Z5Kks9O69ax6f+R
nYDvxPt+qvnDRS/QN95+eT8UzRXR/kcUCbdWBsEd6gpvGlBMKfZ50gAFvO7+hQL7Xz4QBBP+GRvg
1zGWG4G1r7rm3wwC1m8jjaKvSRcDoqV8ovwTpGQmGb3s3NrVLh7aKj/HFsdNdtI8pkLlTPRJFhG9
oK74TvRzcULzXXKaWJ9VZ+s6IfWsQXuAzH1DFbDoaxX7r6R0EcDPCYXwDttyhUn6oZPr4U5oA6MX
8do3RkigO3sykVWQUuD1sn2Abf1cJxYh08vuAyAKIdvXfgXyWPSNOD2E/mQD1Rx/99tBMyslZYz9
S9lGaRj1lnXb94l815tWkt2BPM/b//yr4aG71FI16YjuhjDWd7R0KJ17ovMe2V5ASxCFZql76+hb
szWpkm2M3jTgZmLHQ0WziB0p4f27d5GBZnR29Plq4c9CULLnMdCSmASvBhnUrfXgEmp1SuHS5c0G
oS4ZtoZAQQfUKIre0Vo0B/Irr3vSY3uWNCWuCzL4IGcxjLiftEVmF4kxRL5071fFKB/zDR0zIGov
e9frsMaKNMg1hnXSmA6aya9yaSS1ziUO11WCEeynExZlPzgLG8gEvt+pxe8SwRexwLYF9u/Yox3e
f00RaVQxgNxl7dRIminV/T0+jTyBQvxzCus309+/UnoYxGWYl9X/feZrqHRxWEJgrPSVvUgvCgm/
nlUvN9SAiFYtEx5dYiGglmQ2tuBVb1GOgeezfAAJsVZE5jtQjDfb0It3EdO3y8IYDyelg3cFMh17
ckkjvq/CQFoczZQ+MXL+idjlTjj5H6tjr7Sim1UfADhtzf1AGkIORHVZksui6rjcKS4QFObCFQFV
wjiJtP/7Cue/VJj37TowNa9B30Gk/DQkcrpHj0g4NsRTma3dGwn/mGAU/i2uaMvIa7aAs6lQy80z
HcQXGRKFULEOOnbNf/CBcxsbFjgD4fLzke9UoMJ8yGU1lOepl6/YyW4esUvj2s/hLa9ewGARu/eG
58Gz2IAkZ2FgSIZ23NTQfZiftiFC++u3h0snimT0B4JfIqvDR45khUfmnxIbZ0iSI+6XjqqhEZii
E062hqEV+8hS0ybL3Nwhf5EW+WOakXsNmra6SF/hBTs2REQ8FsmjOGGOnTR1A+i9X4Gvc6G90ECJ
jXipbBcODvq/+p9iLL9byOrMsQ5aYQyLxnAOK/RNPqQglZZ6w0bYXLSP4ZXmjXyTheIBkFrbzPbk
YpW/h67bigvlIr6IqJOLL4hh10pYMMmZfYOJ8UQcVqoqPeCrFcVIBYtX2q3QiAPBdxGjWm8vyC60
mVHoaJor9MPwXN7CYkJZQGOEhHCZSAsEHtizdNTVXkui5cI4CS6f2QUb1X3enrnlp8i84EwZ5XI4
prrHXmtNhnjwn7ADa2ztuZrhCbzor4vTRIjE2RVOFJY0b8wNiztArQ0CS5v0/8aopMSofQkTVGia
zJ/7sRVUtpDcl38/YuN8Jqw4AIjcTiJYw/Z2ntVWgE0Ey1Wx74vRbEHI08vDMk9YACtjCP5Rt/xf
fSFtgv3WYttgE8XFdLjx7z76a4yitqo7goebXm2XQZ0ioAh3LRoHNBc2SqZGNpV7AC8IvKy8aL9G
2hEZUgtOb+ltmjJ44IdsVWZMAgT+Pe9FMt4hbMttKQXM6IdqsJVyAAiM3LeOUcNWo7SoCqp19a5U
i6ZRTVXhRQ9izWP61H3MIp1pevCv6/MPWDV1X7ZMMs2s7NrqRLr7/dqXgAwP/rNtwPJc0ndFfAu0
rge3ssB/obV2AFAxH7Zjo46EAUGIudZ9bKYTpe3iunzVo059QBvqkZEJayGKEYp3HzPqrxplUGBe
GG3ksUNTG3BupgbZT7D0+ZW12dAM+LftJsf2TFQCKS1EJV3EObW7SRmuy8H+TzuNnvaql34AkKln
KqgfUzOHszda+IYYCU3Q+rVJCj56RpXZUKLf6fJ+vH+Kdprhg8FSaxD0l/cfpOa66HRMDft1TY4Y
hy1CqSljBs4xjvnWUy3Azl236gNiAj8fvcJ9YAPv2mFyGbBKKlM8NAmIDwer/Hk0ChkZaCpN6w+F
KmkscYgPAsYS3EfJ/W0u9OfqWQLWO6rIJEVHcLiaqNxmGLWhJJcHQJG+fQI2wFjiyMS1kDjM2/do
y7vAxJcAT25zOdIkickpvXq3nzdBcX95i/1mm9dv3vAahDki26KH2Vo6HZYi6mPue0OVWCdyZy+j
lmBQFVsy1TQ1wx+J3PDbdd5zjgYOpJOR+IwlVYxIMuGbeIbYYt0t2ttQYnuNzqICGF0mKUvVmB+2
rsmPg2UMTfux3B8AeWUpHhQsRHDLWH627GZyxF2dSLSWIL/48gtbgIdR/yAfkB+sTLddfV1CStNp
KklDxILa9ugbDr99VxMYvqeOcteDOKtcZWYac2JuuBJ+H9btyNPByNlugdkdYxXUeHUGn7cutzns
3zb4JyCKfpgn1HXLtXmwzlQTZPoXSKXsSOAIi/UoJUwwOTDGNoLBehhB6pkM7DJ0Hl5Gz0CeSPqL
1d4n3QirSJSYu7IvSqSwLApvB98ZUHd8LOzV0zXIZqQY5947HbS2QNm6Ykay0YDuhYh52DIRY46p
FRDSAeVxES+gYrVhvpP7rN2nE7qwh7wlupbSa9TnwF97bTBjGK//zQj0G9sLP3ytEsxuxYmfg/1r
IL/E6+MxK7+gGxM23txteFh6an5KJSigwJggm66H+Fys723W/oYcO6zQkYpAZOWe/8Kmu1N0jX2g
B7+88tvVJPiuA3bXSRtrQNNMOBWDc/gikil2xcSvP7i+gMbce6tC0XIlDCUt6BsZDcEqgYk+R4sK
5C5tfhhjT4K4bTtUsuRxr6iHYXovGsCwWT1a2xVjGyAyVnJz6xa65kAe5C9Qg9as/6YMbqtwCt4S
842DdhYDVx4EoyqPeQlfP3/Vv0B27ghZa7nOFdYQbli5FeYJjDUw4GNyp35iFLTZFQt2GJBAsaNj
yT+d4pyGVxj9xGFXnepLRQHPkub3hYvFtLT2FrbwA2MBPRIztcOVVGOKGhWY3WVJTHuwfT7Bqnty
g/PJLS07MvBceSNrmIXyzKfd2VCjD06ouigFTmEkY3Gigal4TBvc/SekGWB+Cx/M/OIsKSXP18Dw
jYI2Qy0y35HBFu3DJCC7TXdI46Q59jqXwGH6cg87xYXjgfCgSUXIsGppPcHLhVf7YHFfh6qZMAKT
1Y5geAziQv3uoU57lqxrWn1FWOYoy+shXJkr3hR4SlZLD0/3VFzhEyRkgVp9+l6iN5wAJexnmQ/Y
b+Z8CcwUF0xJf+msqu7FOC2IPkl2DW+amETzk6I0/V5T0MAt695lS2jjGszmRAK9Lnz/kf2ooBOr
syEMvdymMaP4/RO5yFiHGJYn6JYVeKgd4K9H2VTJ/+NonXZZJE/a78VZn6zY5AQagHb9iUh6RGau
xf/v3HLYGQ7eGyaP0oNO8T9k+AWAGjddgURySP97qfmrz5fghNMBCN0y1eTi8rV7rgBso/JUvu7n
4UsJibPC8+kLxUbuSiUGwLU7yS+0xZFl0W/cpLH47r8CbzZC7CT7UxxyIKWbd8wKupQBEtMlGtxS
8gPYEq2CW3JwekqbGm+l7PNPCXY43v7O+CQ9aRk2GcC3XwvFwBxChJVp7bgxzGb09T03gaJiiS5/
yHst9k8l53qMDTg53dp21ApbIuiSTbJRvEg6Hg/RI6/WUmTuhtr1G1SZAqhwhjA10/9Hw6fgPBlG
ENNNbX/Cs2o66tu4/EmPOjLPt5RLnD8UCwF0Vb7UtuMkq5VZh8f/E0qSqT6sv0AYPOPkjGTBSyyQ
LWIjgWvChW2fX+88L3uRdT9cwZaS95yIImJ+KAsnumczpg28OrmhI/5PQeyjiW3RHmInnN0wt2Bk
uic+SIoxp36wDwcGDyiv/HFFhk3UcOXF2D6+aTkiN3ODUJSy9SgZEnYBU7MlyqEtOXa3D/CQQBqI
5dKaDg206QxBFTJ5RYiuPCbyhsYMRtXq0OCRP5KJe5DMGIJSPzrdW/W0HORzT9narNfflnrBV4A4
yu73RXhJh3ed4I1Vk/okBL9eemSqf67BPLFMpJBkSkfYX87rlOnJhrmAUqTPfQhYXCE5fIddfq2/
GPi+q4PyJ8atUEqPiigsx/xmGeLdyAT+Q9n+HlhqYOG96AMaClgiSJu6eEHqSRFnOAN1k1S1YK+z
qX5RWP9WBpyOtuuyz/r5knzksXR6ouHhwmi2VSknF2T9SZaLxRcyHTFCizzatfv/W03Lat2fXpL/
WhDBucl0IcPgIm8mi12AwyvdOFuAn2NjVi4jLIbXtFG7lI1WO6/lMAeO6pxx/L1tEG0StRda2w/d
BmWXH3Y4yO8z+1NFLpWk9JxTWp58y0yBXUwyBIULsM1DLZsQledL3rHKLemUIASoMHv2wq7HpmF6
NOD5q7BJG7iTnT7VrCokRWTZoSwFHqcXEDx0Rrq3MYYK7AQ+xWJ/kabDopt+LbWsd3aQaeoWnXmx
fkCbFsiXBuAJYhJCP3tJ4nk0DfPSH81ZFgzNJQMQt4WVbL66FhQD7sdtyVRm/T2GFfiWxUkMg0Yi
UyacYvPeNVCsRpslNdB/gxSFxwnb1JXliIqxnSlY0FzNGwR3DGzfVabe263dzfOVXM4+IB9kmt8k
cg0v+mBS+Lxf8gGuoDM/SmFdjtG+U/snx9NB0hTTgleUZJgzYkVPG9rHrlhxXr9Spd41wHTtbhxU
YtsdNUuriMcKK9hhDf5u8qw2zKn/ywOgL7sUeICIi41poXeCMK1e67wVJKeApbUuNPVT2s1hruDz
SUPsfnrR+uK7X8R4e5lESJ99mNRDGD7TOgGAanWZ+s2YJFRAMlmuMycpjyHNMh6ddJ7E/H+izhQ1
yJaXHANTzyig9RzEiRE0tIVf02LWSdsBBg1aDVsJed6MYs6myW7ZVN33MDasv3mN/r1wBmcdxy/Y
fL1zhxBQtvd95xOpxF0SASLiu+dHnIIoZc/YwUETK7j4gHAJkaEBwSwLFzohyfV0fGFVJQKj9ave
WuqmmBulohDDFZnegeBF5+lz7LcDz8vKBCfDpQ61HwIsuEaaJmpoVtaIEfYKcKyoj1CU8q/onZaW
NYzyR8nP6mQVilO//qmqa7xt27bXXPt5EILwJNbbxsL7K1Pw4LZGTUdyo8reqrGFGnBpWFpYJj7f
xaO+ASK/bbHi3gijWkgbfmXkI3c2KvRGRDfANVxkaKtCMMrQQfKP+Lu8gFksK6YLUn4x18ltcMbz
KO18lpew/fmPTvy39g9/nOFETYSksU2bZttrjRVq4+v0qqQSwytNkqUDT8U84GOUo3BwMV1N4Drt
b8fHoYR9EQsvruTzTOraLBPf0h70UEkQ5gBJlKO+ERbRVo+SaTn7ribQhH39C+/cY7QC2gkIr1Pe
VIdg2Zi3tgqjJcBbQi5O/xHaBycJJWSHv5qE7vcgzM0eeHSI3q0mmP/BYU0+tRjg6+9zB3aT64Sv
3XnG4Wp4wt+/EnMQD+kBLz73Z/owbaVIIxE9w6neaglowqJnIoOwonC3pFoYGvDNdfqAStuzobS+
wKT7BmjcFfcxYM7o8byR769WKPmi+syVTgUm5TWmeCumY58HiTLFQaXFzvFZfRwxt98Z/kAfSFk3
FVycdpKD2+xaPm8fxMEFnK3Nrazdi+hIPskbvBw2L4PIOx1qWd7fTUz7lK5rXG26DNoJLVUUj13l
+2DgYYj5LzAb3I+rEy/5GoKzUHskcojUQBYMRi5ebUQ41eistWZG8Gu/5rE7bdpMu7NdP6eIhsFm
0LPbeIir9i/juu+hH2nGV/h//b/OcqHbeb9BGL+KwPOtp3FOyRPg2RJgvVpAVCGoerUe4qgNzxIf
I0X1W6yiPai5gVEALqLEvM4/45nM+IFxAq1+qDMqnl/sEs0MrZintCR3qXoJT4U86Cl53o/6/v7d
IlLE1jQjF5GhGLBD+B3FWwnPOg7A0wn4lGTYvRXJZKdluv+LBtKIo362N3fIX+rfjAC/AGKMlmME
742echGqaLjW1/DvZVwonXiksKzJ0CIeFDvzYSCQ6saC0mJRn4/FADwYUBLfdI09HEGdr9YnzByt
QFH2NW4AiST1iHjw+YzNkQj7ZkrKYYVCXTQGvhssnyWfM+NINSQB4O+VDOGwD8M6NKVCb639gVSe
iAHN4DtDFLUB+JzmzQkjCifQgltgWWhYtgwNCdlnW4Hg88Dj5JGa52Kco+bhQlmBgPXU25ie5FN2
9IsWvAKFPHht7+GN2cgGHJu2yZmbe9CIsQxLbhDaa3gNBy90W9KbBKogdGchfGysZrQIePtXyJpX
s3yPCFkqVbxgJDZNlpQXacvjzorYgcyw77zLA22PWWxinKcGAhTN/xdZTNA9pdzRkz1mqodN1cfW
Rz5LSTH6TXG1+o2eU8wmdOQDE+cCgaqswPQFjMDtyLkJYiiu6Jlyy6RJ/JrYZgV2Ox8a8Zpy9Xay
Ys7dZLebpLbcoMPUsUdFpfeKO1+Aeuoy4pgHmNRKNHns35AUZNNrmPsLBdOIV0Ikwwk/ESXgkEiF
zjiHUDV8uYoDPsoUEWUSkVcjsQQLi1ar2jANaTC/ncvmA6hZ0LnQdn6e2AjAo1P40b2C4NLKTvIE
48fponL397OR1Sz5Rm6m5VjFJKjtbudtiRZUBA63tQzNt3c7ZEZHiWBxolDmCmzECeiDPJDxDWsm
w/8+3ZYd0hLop/ooYKx8SZ9l9g2SpqGIC5l5JVMlqSacXK6w+pjV2iIW4EG4CnQ3Xqy1HWteD/91
hmKwI11YPoq8xP0svSWBDROFCSyr8va+O3aUayVpOGv9ZC4vlY1QdWEiRhdHsvDFBNILtAvLXDOl
GJF/CJoKeND82cWfTYpTrcFgm5/Dfbe1ySqgJ1/comdOHjH/jVr/JpyqGNhPdB09i1zjkA+0AAjX
GxaHkhf6CYWwDQgae2SSxEUDg4yqHnmVo/rT7v5VCDmMjXHgr8v0+7QNP/CTq8OWqZUAlXs+Qe7w
FVaIcKil4Yn0xDJjGcq4KDaaIsn8AfUD7kS3L8RWM8qSryTmOiC3WDnbe71CTSVJj8ryc/bC57b+
fhcRrzj2OrgraW7SuDrVYNVL/xG2iPfCb4w+kuXuzCxc2OfB541Kb816UExPl+uOKdgVXGNvONmd
YTgWvwySUYNNxReNocGOacHvsPRJOSyIYC8uYIzEAbq46VWaqrrplNdjVBpnINBTIjzLzZ9VQ8Zw
73LqqKTLke6FHLtFKcEbv3ZDaZD6/DQ3zj5gKku+jqw8JsL4UbCdTH3+52uWvtpj9VBX6K/zjx+7
OxVhvkGs2WNf7VjhG7dlC8R+6ImB5Iqnh9HQydRTIg5Rgmydwm+1ZYg9ztyiBK0jJS2bPhd0DJ8B
mTfGkuYrwuRiStK6AUHZ5TqT1W5kkuTg2uFVHzSF/UmmX1hcxd1sGK8tEaiIBQdrF/qVOsKoFALG
tLoTrtpYcmsFlFdHXV1fUosK3t7Ec75DJlKgCSwI7WCOq6wq7pNZMnF1VdmHKY2OwHvLZ0K9cybu
YyZ7OmDL6xI/+OHg43LduyPcDjf8r8ji1odTVzZ72UCfkAZyBuUuQ5OpwM1l7XmnWXUZBD1Uv440
Xf6GpA7Knmo3vaz1PJo5IDK0ZgQl683+DXyZEEWG6dGMcZZfH27fgHy9gTdMHDQh76IJHzPp2iDH
XabWsz+NM/KfIoZOvT2RAqHubpL1IvMJfARbXyDLZrtpYe3W3wRAaIXPHKfYtcJ3iM2XVw9Vkole
XRY8YBhd8+g5Jq9y2+Vv7ItOa9mC4zcmalWwb56udC7gM2KpcGTwiA95T1PNNFIwai0QZPSaY69s
7TBj1IaG5RCo7+HhVo9xI0Nopf4uS76jPLS2ntGwWdhmHX4QM3hP/xno3pc4IeLTbpdGWpYpxkDX
Ik14IzRhmKPMFxUYWzTeeAmHi4OQ7dyhT3yBd2eEXi1DkcPIAm9e408iPPGFOzPYk93EM86cx3mV
jV2iBb+plhJdgPTFVn5GPVzZCy0h1kWnY9jaCPIwnf5ZJDSil/Zy6vUHXwOzNanDxMajSAsJmD30
KpFveaIV/lrKjNmvEnpQgrQT0rMWAWb6gpthnLg0L0mXCl7xVKizmRWf9081lbcK70MtDGtzqTDJ
sxVUk+FmWzWDknZDWPtozqk91kwG58Qklh4BXFh3xBg9CrzVkYwXk/plljQD8h/CZPoNgakjuWpa
wp6knKrs7NntRJ0aJCGhD8ec2XACp9VCUEKaCEo0LaUPYt5m4nu8mHw6+PqqMzfZzHVmNEB16QZ+
oKRFx6OSP45k0XdjEKj5UguvR+jdz2r+tUCXRxQ9mM3Y52/4bVSFI08UemVEHEmNAycl3qEhnFTg
qgZZVnr46tiX8Z3kDrEioz0gqGgpgH3SNFQKC2k8MrbWT+t58uWvxSp/XFgxbm3z1NDb0LzzBbCh
QWNkmPR8n6c3zvGFIHEE3uupDqfsHVqy8Jcgrxd1w46CmIddB7Hy6iYcL5dIN82KuWgJwOaFKY4c
zT2XwBR/E3cs74W8WHaWAMBxajlJZeBm+oEXs7aDZ8RJ7odgloNHxgi/jksaxigdfzE5d/RFZuXl
PDBkXhXwvT+nkU46zBUocI1/bZcdUHdbZJChE5EsuKT60HqAdo/Upvnvq1FgenNMp+GD2Ra+B2qi
voxKrUXkxZ3PA26SVfghpHEYcTVINc7z9b/AMmiKpm1b5vaJfe62C0uZhdnM75KoG5unb97xfMOe
7HtN9O9kfETGP3UORI7gBC6e4KY+H6xiVYgmr38QrqMIshGjZEZowHFIV6B/Q8Nlt/aCkevOJsoV
Vlxj1p1fbHXJrKkspd6kCEnzAj4t1+PGt1EGoV9PEDh5uQXIy7w17I3Le0+oZusAWEudd3dr3fNB
P/mSumskFsnhCxAK7iZm4opL7FHRMmoOEQlLLKhRD4MSYNvlmyPLeZMzbcQOuyBVBmPlTzs70nIz
Ng9iZrXqhU00RNH96VAFfyLOoDNgz54vMXSQ32TMfCaIiv7pXjqoiaL25kPdn+RuusbJ3r6Jph0J
0RDsM3ajH6X5Jm5dsLd8A45dkQB/cQ57ZacAuSAAWt1c2tYfn6zCWODnsPnDAI0T49bjvPlXaOzs
TweBRcz4W+Q4aE80IUJOhvm2y8vheuXmZSfkPzGyb+vpQIHOuEUcZg4iPWHN9s26PY38YP30kpns
owFOeb5XrMehrDI11MAj9MGnyqjeQnk4FIva4TL1W0+zOfiFhY8XTvwARCLt9xX2AW0A2W4/cyrs
EoqcksPYIju/Yax+/TkoHmnamtm4z4x/7rm4dIAMIGThIAZFV5Vjzk8G4HQRi7cyi4B6oHo4NJXI
J3UQUEpPne3qnHSS/ja+sVSFW5jagrG9kC4b+m4ShD0Xta9mKZrUy7D6yySWoRNgYvej783SEg3o
IgAlRl4bwLnKjSUyPC/NTd6zYyHjEE+NFc132+LRsMYBicO5HKkh6/XILudAitAwFSXyb7CaDOOH
kReFnK2xi8553oA/fN9MH6PuHyYHLAw0poj3tCpJIi2oL2b2YA81kLQ3KjtZ3Wu53ELAxKbPEkEL
5H58N7mC2BzZhPa9mkSdCfq0O6PGo4kSEaumL0i+T2idiNh031yfROlmO5oRidD7Qi7NxVup1fPv
REN/zUE5AkyVgrkC5dt96WQnhuHyTmWgfdEBCYWhqe5zN8wZQlid82PhVe5ApQnDozhHn2zZ1SkF
rNk+Sp7AU5kWYlx/cTxoAGyqFJyEm4gRFBYgJI5hTLumFhMHyeVgM8DSyP7MxzxDD4SQJ9CUBUht
lwZOxdQuEXVJkUjM2ZPH6jERMcNGqK/7lPx/uzqmNgX+yTNya5fqdNJaFh/Dd9+AclmLZKtTcCBN
QpfZeLYOrIcjZKXo3KozTxbGxClI/YBRWXgFk0CWZmGhYuYHKuY/oTYwDFP0nnr7fyk/iRWX2T+o
Nb94iOX4Q0ne/TIJbRsckDNMBvgv59yiMY3Dl8YpCKPy+JpNANLtxo2/Cl7Acq0C88DNBk1xwazX
PQ7F3v6HFWKwCj5BsFNbAFO0yaCDqTXJEhVmQHiHwQhTfLTMTvM2oZEGmxJ59Nft2CCcGjBKNe1Z
PvaVQfzWtHE1gKmaTI5S6zldu4z59W+gCNZcUjnyFlTRMaKdwzXJ25Kz6GSXfNB7dAXxjJZ5Jmem
fCfslW/4uNrvyv2ZpQ36volz0agdflono4YCxTgLccBZM7Mu67XsRuF+qpAOoGUa62++lVhqrYDM
AN9vhYsejOjVN9tdqF4RWFZZq37asYyUxHJJhjl5p/Ta0X8sr9xjUdkvMYZo5keIIEn62P/i2h9F
4fmBN4CufMT/YRhx93MHvJFzu/ZHWMbEDRZ6jt6W7i7URogsjRHm/Ki7oYGk7beHFkW+qB8Bv3P+
im7A3BTrkgbIiaWX34TySAkSK5MpIgj+3F9z8bM6LJcf+i9+rKpTB2fYm20MPbfrML6wI9lQYdI5
GAFuvr1PBDMCcXFvmxojTh1rPFc+7DxGlr5e3CNajd2bXRZdxFWLk1p+wp3W+65OWOzKAvmC/910
ts3Gjui3HqU2vMxfQRRA4aMY12aOw3J1T+hybzhmhzvnjOwbLXruAcV1LMDbUv9wEihu+Jawafoe
qJ+XoMIoq1tZQbzZ84QtzO72zIcZvJUtALDZJvgVN4u387roPtl9X8KiAwfsLzyMxv6V6Y9kSQyg
y8iqNgAfLlB0of/ikG8PLOgIYovZmxW34N4Nbd+9u+qZrkJ2g1r1EzHugzd/ILoC1l0rXq9He5BG
6Q2BJkLDCnNtA1upqk2pdpVT/1y+zx0VFndkFW9wYugXvnguBKcDx9YEac+LRdLE6JmNGFKJlCLT
LQBK2ngWXXWNlNIzJdWrMrETKIgScsXpwumZ//hGJImX9DkF9BWZex02O+wX83g4T8dzQGVTfLaT
JNBYbltPMy1p8euYBeQFjJB6SOmUkDMadvyg7g2FB0WN3Bp8KdDCKE6BGrV7pfF0qSAA/M0Q9hB7
7hbJ/PouaLZFA50paUUpSMREjgSH+DZO2We2cmz9uNRLfbvyPF4qpJcqPu0Ffve58io41IuWE6sx
WBu6BPB17p2y7AgOBimvhVxrPOSzrKXPGC/Lkpuv50NlytY4pCx7TkgXKua1NM4C1kb2b49zku/U
pTV+fdbl34fdJYNHEc70ZFxy1pv3SBvtcFxCPcpMvdPIfGoyN66UFpPTzmCL1OBNEqac0qYcg5HA
Iq/YsuVZcSuu3ATlsYvvKJcZUg6s9LxB1K1M6n0204ZWm9SegcJXiR3wPRKeFYPyXxU+mSusMVaf
9Bzstm87P1D35YD8RN2G3VC9R9+6zfmyvGR7dL77vnOy0An3bbmeQSxNudGXwhl5kw/L+/blNUIo
VD4/6i9hH9oHghQChhUDFeJFvqOxnSQNbtYe8/FPzVrtm1u1ROxv/hklgUPJ9eezvJo1nsAkr4AS
RX41k0lHV6QRhsMG8CZ2rN+K1VrQhAoai9oqou4mZQQeu659Os9pcul/HrlCKHbfsOVmqNqYfiKS
gOm1G212y/uavmHm/rJfh/sKvvfFPWv3KbY22tfyVNsom4SfhFSKqBXmYwgl+mAkTkr9BkiZgS9q
tneecG4uL4WqmBEDa0tW5ssnIDWnEmBVAXbShtZ7Bku7+ZqC7sec2g3VL4WiALj6fKZUVAlucF/N
OjgEjHvkA+f/LhynKKlK7uPBsY7ho/5XsQA8x2RCChUKQqPQNp+lnZr+dFhGeS5uwQHitGTP7he7
swy+yYgRdwnme2hLOQEIGs5eesXCxzgi6O+vmlKMt/VFZu65jijpUPwUD+6iJb3B5dZSNquMKilN
1sqFgUW0SHaCeM4Ks8WPJMKbqyHajmzOGxLwqRYOKZF7te2zjkRlauAXHipW1Dl/9rGUiS68c3R4
15HY2CKDGoEGG/mjAYx0DzL7+s6qhEESrUtS0cMWQloFDHgRo/G+OyMIAxVzN7ak2HI7+/5x7Ltt
surb7y4DVj9AcNtwtWeGfNzKjtGjovIpJzDNPZhrTBzBzqRaj3rb9cyqn4LXQlv0bIJ5zcfnrpsX
6gZuLyIg3Y6q7pGbpAHkVGyj+eMwNsb2WdvQ1ZgypvOD4XVfIcKO+1eTuEjnxVSkyYQz+gDVk7+D
T9JyiSIxhJwuKkVeMscRVL1fFnUL67ieqBuBwUuFlGyqr90vHywNUUdDPAgFuhTC8rQZ4eB8qbUW
CDXfkPl8e3dRNm1ui4IZySy9pIoaGfgfHVHPX3KVUQ/C9y3NYSfHeQDwVvDFM9CD5uguNLhpPIl/
eTpwwVZW/G7NDqJVRf14w2TorF5AW4aZ48a2ccsssCRsJre2Fw/TCin1JLU68RUPEHJhv84gZ/EX
muPTxyAz0Dd8UFmzPUJzQKcTPiEtjTczPwowjQMdO3o4bz0RyIZW0jGaMam93ydhI90a97PTu+Z/
b+aAY9UzOQqI/Rr2M7jn4kcUdz1X6eUl+gjIwSWf1xg9ydj3+xXI9zNTWM3VLueVJQGOr8/cn/0d
P5lWCoSXTeo5XnGarbcZBakmWMTrtsQQopielfPD43tRtIri74d+brZ9xkgFaM3tkhOehcQ03XMY
ggeDlXZKq/dV/JsD49cjtqSttF4R6y9ZnosmOFMjWa/19FIZ3FRjuVkD+p9MvGL9vEfmSxTl6OIK
+8lx2DyZPesj9uff5MyCbdY7izX13o8It/PLCSjoharVZUresJJ0e6H0WKPVyK+ysNooRSw6BZ6+
iusEzKazUHtDwEafeu5fLNTGIZ0jjAFZm48LzLGjdzBGaTRvrr6QppDkEEXcRPSHCOnoFkKsJBkc
FAqAY7MuUdfOmsOE5wIb3mRY85Bxs6Q+if8+ceQMVCUkgV4kAzlkMT87rk0ahunDNOMJJ+3FwJB3
8Ono0E2DLtvu5zWuQnTaDGBX2gnOZnJw1uL3/f+eCuv//1KdFf/ojsjUmXkJss+KkQyeDUEzOPEW
UPMHJqBVg8j+wZjavLwC5fc+AmeecjBt3D3NKRzU7juNqL9Dm/fkmBRm4GeRZLSAz1Rd3GkJKTSb
Z2po/ki6sRciWm1/nbjSute1ywa5GkZqMYpnw1QJ0UbIBPC12qBOWa2rku+phjtOmGR+l79JcwtX
sE8KyFxO89UyK5wsZEwDp0bdtGkw6aujUOlO3hWgQloe/c5uxZx5IpZD3bjCp5kPFxgQxGQ0XSvO
YlVsHQrmBp4P0FNvl+S/ENlxe+eT0zP3I30uFbsiR5XmtdaWOyehGzup05msvU3RsAKY4C1yLdcm
CON2SR9AjJDgY1Kx7A80XIWdCg8m8akj9lD7BArlABFrbkbN8Ul0JLNaUqLUGDlKqqbGEwlqYib8
oopVVubpzoN9ys/ND9wfrszxwkaG4BX4BAHFtvyKGEtc2mvsAs0Pvu0z0hsKtRvk5MS4DSaFhugm
Kg1VDfUO1VywqPnrcjxpVVe0iVv9BynIHkCvBjOuB010NbM39E3Vw2K8Xu2GMQWVLrQeNrQPgJLs
zFZnr3eFm2kXochLP2UfJD/V6654XR1X8DGB/I+9gwXk4eu/5eAiQimqLivyPYgsWGoyyoOsxoUO
EQb0WXt3h78W0mko6XfPcHq80/rZwZZacePc5uPa1JLc9XROed0WG1+KQisgzSzRjOabOX6iU9Xj
GEPuWCZuFP25D3l1o9gwgDcTVDpvFxZSaIBQNfhdGULsJjsWN9n8t+F965b/cW3JZ2ZxBJaQnsvT
O4AFoexfVpHC0yO4Hq6wefV27P6sRbhtnF7Xo2lEwZWqlZvMzAVPy3C16ySH2IkbE/7B3SeXDdOA
6uv1zJZHgNgbO0EDI6ptK1UqKYwErFgQYnsXc3ped1naHQhZ+R5V9+bdcjVuyukyBnbfvvHunGj2
8OcBONDII1jlcFc3u5lMKlCl5NYce188+VnKNI5DpGLTeu4opUTyir98YNRCNSHd5BEU9Bg5uAre
6Squ6QZVTx1A28/Nj6O+wxuAZr7DHE+SqAtIFxSWGdF/C9l82OYcSWnxniYY2q/GQk1YRysADzuD
6VKH1NqYiB32dmznbM8k/Z1pqrDsDkHtrBsmXBXUcqDJitvr1ZoGE6Z2cfqViDZsmT4SudHdZyWo
aSF3grTnaaQA5knETLCl0MJPIlhNWNQFXOd7pY8RWFhirxB43Pr8aPIxYkxgtXMSK2dUNtkzEIEm
rGMcZBoDHRTO7VVS1uMbxuvYFwe8W/ZkDuUJnwc3jjLiIrNtaHZ1f+EtAGD5nt/nZJSoMsHkpr5e
5o7Vlit4Y9RBu6UV+Kpq8iWiL4teA2G3Fv75uzOIXxj4mwne4GvwxWxzGE4Y1Knpa6hNsqyYW+uO
wRnY9rOnKqMVUHSSSfu6wsHYSACEJNo7LzgAPAHR14P8zesiyhUmFv7d07E0F6yJUkWRo5RF7VQt
2e08PnW5qrLKrDBg9/ODdfR09pwpomeAjbRKvB8ZqPbUkQSzovjjyYUqtQavHNiUakdPoQVnnE2d
HanI/e5ZPj2ESDBwjC8nNjpvrQYmeXQYWyRiEwhck3sf7R6eXqNTVmdP/VQjhz3nEKW+MJ3vQEU8
JuhX7SY6OESi6fq4uzJwwf3SmOaXk0HHQlsHtXzvDcpYpYSkOMcoScf703GNC5TDxuMS7FcTXqcF
TzCAGPTrMiJnRPZ4aR03KNsuic1DtpqLFMszloyb02+vyzOZZkEnNQQpRtHkIXEosgeLl2khqEb9
v4GgTmA96DqFmqFhcciootj/fiq9B1p6YxXDj62suavN5HOYzkX6U/k1878/U2PduegNyewJIsXL
ocv1VfyKJLIPKhKF3GSFPocnPkQ/5032S9qdryIFTvvf7RJi/40HH6yt7g14SZSCfsojarZfn2eV
UP2byK1aLsvGmNbbxYcKrlravjVFYbO6G//jjZzFth8aR2uasz1C7YORMCr9tkeZ9/pShICYb9Nb
sG4vr6gVGRZgdJfQ+DLDfvb3wdrOr4pkIR3iDagVwRqXu84jZNCD8DQX3svt8YJSN0v9VeLbijmg
XFemGihYeScBKMeSFwgKLKQ/fzJkKxxTBRxcYi4FyPLyeMUc9QYcghv72MGzhHXOUFFSRgI98tQ7
k7BIDPxvl+g0h665jq6/y4HkX2JW99zrR51TqgqpmvO+J4I6+GUXdqwyUTn08q3FZUiqAUtOM73g
oZtaXkj9y5j4WTucR070/NPH6db7VV+hxXAnxQ6MHhi+hqhiZEm9LvRmQ6xWGs2h1xn+fXvGkZmA
3a5CLOeI42Z/JoOJp0o/nJWOaVuXqQlhNuDTRw+0+T1JjH03VXuC7uY//JGOmIVIqJ4CzQVl95Uc
pJO0t0ZkOWpFSscOcytw9kK3nmTzu2vMkR2iponMHWBhwGz98PLgpbwbE9MI3RgUUTkgYP5COHjh
w5rHx87RNpdbw3a/BMbTSkbrJUp263AOi4uOcM5wctzSg2ThbmLbNp8YaIv/Ebyn/1xo6ODf6E4G
QLzeNHMOsanWQ7NEZj0LYt5rjbA2/wRJxf/vx6OgTAEo/ZBwAdEwnR0NDv19jomyUMjeEtalsXBH
YCiYBjwbDV/G2MxMh2K7Ub95kaR97YfSGZgaFvUACMEYw8wI6DFy+pvqZ8yIOKdmnbvv9/gq8BqH
m6d4eEqaLOr5DRffTqC1rSzVrdK+uYUNxEh59xc7yqsmzdX1nYjuS4BiHQ7igpUtp5b2KAC8DQnT
ZRUxCbzeXli3yk6FVqAJRLddRpwn/6xqrMPuu7+l7IGZU2F1smZQEFDbiZHbaVJVgQH4Tvdy8kXm
i6f2JJ13hwyPQlrt+phjezBK+I+0SbZAUKbBVhIYd2AL0HtydpaYlsOFyN7IrMN5S9HDroLdD5bU
YBL7CqHaMZsV+IfzJQpBCsIUT3w3rkTWnIJ8nL1o/H+mhgr0scVQvpmsYiAUEwUV6OxehZPHCsj0
RKX57zYfMMja9qvkmd3XuMX6jdKeuxwDDE7Q8zNkSJ4QKIEOzn/2p9x8UT9p+5V/s0NhPC++EJxi
rRLDClB7aM+KmZ04EqVhcJzcy37o5+XXq7z/u70HygR3a4N7ry06W0C2oMIFyluUUyOPSrcIrMJ/
qr1Et41YI0/gfI5C+eybYCG72Q6W7LLvP/b95R+8/PKec1i8Qom/pYr272MFLaG+ki4hN1zc2n2J
yVKBRPxzdDNPMkqU0OUTA8zqd3RBXraW4RmfVpupv+VHvAB/Cng4fzvf4sb+Y2ITd0OrGccPIHFo
X0gZy02SIdqyKoajlP72Pqt8gCiwuiwaks9e2KNE+uCYAI3xrpr+i9iGi1DLSJkpBoi53foeV+bS
xqEW3N+QuRml/5Ajqj70c0bTBLeFy9bdVuN5e67N1cYMiIGx7jeLFrc4zsKYoUZjTkVl36fJjQ4M
X6OiDknAeFgm7PfntIeEIj90xrzg/0m6U8nCe+pv/hDPAkbXQarZ9do1BIvfjFR6cWkMqxNZW+ue
94XiGGoxqmOczcgHGyH2824x5rQh/EtYBZQXx/EMYP88ihREzEXJSnkZ3u19NjD6aJ18YN8pMIN3
jEErKnwIzEhtKPU3h1hLMq3ehHDYmFAIkUlbFG7ossVI9G5h7+ExDAJC4rSGDJ18ZAw3SQcNq0+x
VYNQBNDLR4zB9yMhbDSqoZ0/S6ZnGCuF67RSXcI5HipR/coc+tvolU2caBiy3bw6DPZPEdMHaxpn
5vOnjRa6NsLrDbvQ27o0+3IHYA40cHPfnuMWTNGDsbaTeN3Y67uUQVC0SD4OYvw+jw1rFFZCzFlP
qPzBtAXno25leYV5nNpYQHBePqcXxkt+ebrMf7Rz6vvpUns3Cme8epIdlcURI6zYAb3tXRGi8pTx
Kze0szam/83M0raRZe1yR0CYsTVVHJfNGGTYCUm9pb3/bkjvj0a4yuKdvBUjHdBeNH5+VK93mGUB
e2jWyLgl3CL/qBlygR9cxboAK4G6KM3Xhn+Xe5DtsWlzdvosJt6BehKNI6guSmRFSsinPbt2skpL
fNVKDcdziHPSpCDEcIjdhjFVWlEdPDuIdXUMPAOz00lGw4Sev3GEPG15BOZfk5gjAMo9Nf+CcrBR
iAGHs9uUvdeUKi9a5JedkxIRrfZ7ARD1ROAvMv/lIWu9HYRcNEQQwuMkOw6oxkL9ITmIv6DWNcfO
+Fs9N9hWR7SXxuucRSCWxHro1tvgU4RkPELwy1222WIubkz0cjgTMBrHsPX1qkb4ffv1r6nXw+ds
tRnfOvQy4NfGf9Mq/X9MTl3+q74ZLSaTVg8xAbLbYtU0R5HnF88s0EiF4RsI+ERBP7cEV5yNPUO2
Rai1jEVFxnLiZPNecQxAHZy3Aer2neRvl06DaWey32XPkui9lPQgy+zY0g2ullC5OIgUJ4J48QKD
q6cazg2VEu9Y5FZWivFulXnVoBVEKAhzbmQM8xjumdFIeXisr+2elC+pMUSROX0gdJO7mYk2eCHU
/MZhwXNkvnaE+bIPXjlHQ2KWiZxMHfNByFrEtVcKm0vUBWEKL8lyjSLppucq5K4g7wo4fVZGqURL
wELLpmXXlvvAT1CRkVnTEc34fVB9DueCO8drHqqQdmtl5HwA06k7t9T4Hh2/OKTkC/nfSNzh+rq/
1WVBTgwEDzPQ5c6q5Znf7jNzCkB/LhTVd2sM9gcB1SP1gIxW8zdBbHYcHBlKf07le1P9GNGAndnP
oz+gazcDGia8AG8YBts8uFkTvDsTVuIUK4Ofd3i5gXPnVseDaFLo4eEHEm9AHlP2RbW0OYdAbGIa
b6kCQo0sNrjaF/yq1j32Kunhl4fYoyxvqXgTnKG9cwO/RXYUSakvgiEXMcz7FUhoPQGw7BRK7xdb
b71nB+uIx2fdknac2hqk2q5uzQSK7Q9F7iWLaT99X+SqPvS2nheymayxH791gzdcHyxNLiNLC2Uf
nCFCO9HD30P+3igLYB9h+lGzDKNuPAEoxF6ptGTaa5TYqvARvzL6ojrVjG1yCBytXjLN6pOSLR4K
b6kLtxECWZ8apRxKXSL6bds5/qj0Do55ydg13+KkU0S1E4W+0kjMGCHDvE1XEjXoJA5qBWgwPzrv
ON15UI5IlAQtjRRxDjHD5nWEjLa2cG8HWSxOAbhmQW56x25kuAECk90mXNg7RYGuXoz1RMES4roU
n+jNfXDdi34Y+H2N2lK3RkPN4E842t2a+pO1nuh9zXns0Mfb8ftk06MyOABEMS6hH45KAaPTPp88
21nbVF8tiIaH32hYj+nnNR4fMMy0EmS7zMIxnRFDjcx5EY27fo82JnTZqWYDigleDx7lg1PqC1/1
S0uQZ4RYBOiGnFXWFKCtjau8rdIQe2Z9s1ZSZ3M0asWZn6C5pNg9YjN2HU690rLWLz1RfvM8F113
IUyP6BPkpxowRpqXAV4S55qzPybmDIryMLKk2Artfk9sR7Cdmi9/ddWTPTsW0vzfRs4Ys7P1BZLG
w38PntpqFvcFn3cjQnGDP9shcYJDzXjyplmC7cb08imTKk0AkEuM72N8cc2IZMC5hAYOZ8JH4wFo
ZF4RZiG7PGf7rGDsa8OSAKIDsjqNnh/JQRwKcRx/kZS9bvkQMCPUX8fCrUalTgl6uaDLXRKBU2EY
mcu6Sdjx0y5ZtqkTok4g/Og+VKYhH+T+8RVQ2JZqHCEjNH/a4z2k8mcfnngtis30TSKyjiPC0kTA
h8AXnCp27XHs8LCXYyWZsZ4R80C+XkIRHrPID/MwLJUNoZrBtOd34xUnlR9UaCpwGQ4AIDRScwRF
iEpuSAdwH13+FPu857YC1XbelIvLFuWYw0ryvb5i0L5L966I055jvJsSEPRB+6KNQVNde286muQD
4j4OvNhS1ai9Q7pVYCsAQKi7TqKxH3X3h/l1VrRW2O0egVY/mjdz8N8k17q/ahckOCR4uIUPnT7x
o3R9arRSH3hAKJl4Oo4IeGaRvf7en2s9AbC96vjTSMLcvwTgtCrdiBLgasGV9/Vcb4KExRTYzh+M
kmiCJYgXduWAmgHmvB5PHvdlIAlKS1d1hEOhqSIAIlTjiTaxuuGVegmlpNM5uH7UmxtoST997C3k
QnpXf43rgNX+/nfwEyecRcUqNJKBgM9hQIYAgn9mFnPGv95QXXP47rbQVbm//hSTJywCMg5bMEeM
BuyjhGeJw1PgJpBGSsMkoTaa7p8dBuDBwWEbniG9Nb6pNtrYHhW7+vu/bgFhTkxinWFWnWGQyoRu
OhveNjeXfp3nHQj1Sq08hjK9V0Cl4M4a+vI0p+qyCU3ADNoxub9UokaS+iTH016FMYhFgPyV99p6
tTrUeQbOOPy6isE9QoPcMix5n8YrfAUAEISu/LPoi8YDPWGNfEOo33bFmtJdAAxfrK7cgOQWMMs/
UOJsx9xtOrdlVDChpgrL7YkceOddimHy39xOD7j6Gq+1v2nWPdqin6XW1HlwfR8eSC7m2fiL4NU2
6qI6IwnTvMI8bF6naRYTx0EVFn1pgvfnKGrHYHTi7VzNwvTxnx11GhzGgk5fBvdBBr/wQQrpOgpH
ymd21m/aw3m6pGQ/7uoCwtauDXbZ8yfhfMEmckjCfTlNp0nvLAhXf5yqGrh3dfveIP1n/fdQ5Riw
wXehOTjQstVlgTtIAntOQ/AAplAwq0em2i6tnaYvQKxuFFUytj9VXKjVTiuiCVUqO/ec87QU74yl
Dvla5uxTy2xGqSBMPG4tgCc6dwICFYZkMLzxmkXsMlsSimZV6c/n8rc9C7V0WeghzDh/woNV8NTE
3y5tV8Y3oEGMgXuldhG3G12hrXUDvb4zhtFGMjYqi8ecckZASJ2w1MQybNy2lwJqtcYf/dAM0FF9
OQBjQusMyOavA28r9EqEbdXpT3Sj2kzFLxCC3PfpBANRmOhZaNHwuF3WjzOIlaoeD5GhWRkWrSZQ
tfkYctdrO7diGryrq30NexAnQ+BI/mZY37yg1m7FDIDcqyHRqQ4iSmNN+84x8EZGs5wuF/Kq064N
IyB94oPNAXfVkO7t1HWS7zDH2ifmn6K13wCUz2ryWYY6joRyk+ZNXdC6DClaNbM9Rk6Rltqpu72u
rkCfU9yWKRDd0GdwtAhEp8ImD0ysYsrvV49/tG88ZAfgAayaI5yPLi3H8Y8BnypZvmwl12s9GeOo
Ff09wmOBgFzCGK71zP6tDkviPUpw/MboFtSuIVd9P1lpghLLybYYZeKPjN1psTwfan2/ByVAroMn
t5HRfVc+fhj2WJajObUBf0HYNb+cEGLGmvqIxdKqlHE/ezIzCWgrVoY2rfC2votVapqK/hsaaO/n
8yjCNF8KwR6GTEbh+veWvqdWP2NRFPu9xhwPX8tKgCg3WbgI2NC4iIhred3aCJoW6/idgvJf2SVV
RBBPxcOrdnmXBfex2gxperw6YCxFtM/y91ij62O6SKJ9cO3Ky0sP8+x4hBE2iVpA6swGQT+tDLFC
QVdqVaXgA8N5bmOM/prcf3XlJ2icQ4kf9zSTzSZbXkfQYfsZm4fSKFhSAAdlka6wO0K4Hc48RRMV
/Nikh+UprQPql9qimrb3Bnf4VQlI2y51aeMjKE1fWnZ2ofL3WexaY7wlzI8H7a5jxGo11kqHm955
CNNchTYyPx09fzJVLOGasIyCCTrBY5VMO1HZI0Sg4mqoFUA6+nRVjqB/kZnGzigkoTNix3ObgCWn
GZ9wPo13qlRfMdKVnAOM/YXcuQw/om7IyhGNLCChq1myeaPQaiBXpb4WyETvs3uI8fts6zgRp53c
bFKhtfLvgq1Rg/nCOePUCwo5bNBeQAT+keSOxdr4wiLBK4qiaq+NFkYChQta6fv3zCFXNth6aT69
llsu4c5HBTi5njH9jmxWZ8gDhgYGTHYMghn0eoJ+E6g9+fUsNkyvaAje0VdYEygvazVCDu1JSpFG
xflWNA1zSyQT+HxL4SNtdodp6Mf52HOrtKswFnXqIjASvilAPVdWWjMf6/8eLjoaROhADB6p7epf
zxs08e9AZXzhjfNg2gwbpXQ3AisgCj1W5hLBGtC7U2Sby8XJnbmmOWj9cBMZET4PiqFtJYSNegaD
UvBU30xNGCpm0hMkL49elYuE/COT7fZjEum4LBkmtDF1h+ilE6g2PhEFqcagAb3D3A0i9ZlWKurN
k/UKoupFWs+aCdPMkfuk7YcgVCJdl7JTQgmi1cqkjQhLuNPvDFN3tAVyLDQOMq8/PXvIZBpSdQBt
jpCcTjyiz4TRuMUvHv4QBWPwWuJo6VTEZ9ng9wx2fiwoexh/dpGNkgogUqk5HfQmOcgcLMCGhJ3Y
OedcWCLwWAT5pkSVyER5HklM8EJmgLhP45jaWZ48e/0yh/cumcgbn+LmwdzDY+D9rVaGBIhLmK74
knNOsfuIqG4SRjwQ6tDdauei3XDCoJcHtRI4x/M03O0iKmxmeRmaAWhBlz4w9YaIL716bRfXJBd8
HK2l+ipOF+bXqoUXGso/a3XR43cHnng+ch7p2EiYmq+mEpf8C3N7Dzi4j/ZpQpUtWqkuqaYdWDW0
iASGdvC19iQwWlzomzSl35LT6U2L7hWmUHCIWwhfK2STcajgv6rcnIhBXRHXvrGYaq8iawp6aySF
jK6XoaQChpOFXSQkOnggwEhoQJ7AecbSSbsnnP5U5owpQvtIKfs2copc6TCaLycRtnTTzjiJoeaX
jtk0D6P4qdUX2IjcAD25ZunCjWGCfbFMYscY0QVqQq0fID/8+ZKSRiwpwWOnl+KH4IJdNZXtXvIf
K7wZ/lfmpMxh5srrj2u0l9d5F8shUSdOFitc7FGNFgKmauKYo/UQ8pXUifzbrjWU3ACYHQGdtYn2
m4zaSM7IQmrJOZCFWHnOzzdzADe1PVO6lc2TUGZKCRkJtehV4OKNPQ9f2KZkF3PjiVlqMBSITUcW
9me4zQc97DXHXt2YxWU6NcYLn+SzWT1rE5v6stJ5Tj2uz7V63keZRbgF6XEnSvwJyFxBHHVgPQEh
ReOIWjxQShfOS7wkvCVKYxFMt3g0KBu/30QWth/BfpyV35BYsqm0OCe6/63NG98v5nT8rAIayll5
3V2ec1PJeOPNk4n0YXnqoamirir/ZZv6afISeg1kPHw020KB7LM7Xv8tgJ5C02g7Qcd/yLgitW8B
/AWStelUeHQ0qizdP4PQpI0x19lNkbFG4EVsHFTasoXMZCgmfDkZkLMGuEK6rr7fgC0vrTcTq5Bk
f4nUqqlGL1lUXr5F48PdTzJC4UIhzeC0uhfE2J/Eim9f72sDheQHSy2LNkSyH9qK+Coc2JDD/jik
GF9Sp3CEosqZNUm81BrAUKOgLgFNXztvgu1OQzzOyKEVDs8YwdBP5JXSTIMVXqsofCLiIsrDnBg2
xzyL5dr5IwOqFiAw61hcQOLNtzDNiCf28wktN36KTzw0N3NxPZFN5djzurEFgQfLjwlLDXKb/hho
ojoRfE7W9qIJ8lG4uW2rwS38LcADxzi5up3LG6UZK5y2x4HFOH0lPiNDp4i4dddFZyox36DNdyau
+oA0hWJ/uaUJ7CN5Vsr1/qTgCeh+O9a+H9SHTPbXGK2fFamegxGxhGzbIwI1Ax6O9Pg+mZo8Q73R
/AsJRIwkkojgh01J1FtpbYvVS+7SM8sYFy5mL8T/NtmmK2YOLgg/dXVHQrqgtgMWs3MNV64zzYMf
ehdD4rG9yamGToQk9IX6bK2/4dMyXyNJy8pxiwVFo37SFexkc4nidu0n+vvx3ICB0S57r27d4cbZ
ouIA982+RttT89U82AcTCaWI8QTb2zMY0zgIz9aF1YbkRCwtlAiGhLoPEzLZLxkKBon9p2Imzd3x
lpAdxd0/mK4nLKgye9m0L6nUhbrg+5+u/IRL+j7mCM9oHku7BU3XPuOpwclzTJIed5RvwzBa0BzW
iS3tkgSesgXCIr0zPY3MGCb4769kExyjE3kiaF5NdyEec4VCfhgrOZgjvlnFDZeQEoEasZcipdYj
2ylw7wjIaUUnsrJM07B1fm0kh8Qi+5P7HKVZc6SLKGUArH5cjmePyX5lWQLBzldoqAVV2U1dCk4X
0em7lq1Jd0tX27+9EXEi2oOSHkcX1iWzDcg6iuEHL6wxdQaUml1LtjO3eiXxxv38HDjl77202dAf
BqDmtWgsA1lNcHuY0hn2jcByzqW+lAV/EJoxDBd+4UodixnGMvdVTtOrEl9hDXqWhIxy/kma7pD4
Jyk5X+xl07krTtTWGEyzeE55miFLJDI30ErNIQxL+RYrCL3dntbnAyjIEf6Edzn4Dy4fnpKwjt13
b6kNP9U4mQnV2zYgEnB3umouUFpGwqb0jEMMrvJuez1oIJxJ37tC4+8FV2cZ92ung3BTv+U71Iw2
gx/iIUZlKUWq2dNjpKI8L+XhgnyXMssIAUMTtJWKQK09VJCVz5e7MOQZ/lQmWHeOZvpHfnkHst6x
viWycI5QVFJAHQV3LBr/93wcBL90M6ZwI7qKoCMVmIk1ZbtFaI2SEwR1t+V18+a0sG1sS7dyqokJ
2qs4DL6406aqWwLOSSwMvN6Zr/h2c0iRpftfOlTN+622DDD42PPhQoHaV6/Dq2rnU7EUk/3nAejS
mTzFGFQQcf9ad2IigJvmMy13wCwZjgcegu0/Ue4eqOXjfrIJTJLohxYrne3RYeLHiavjFYA3U7T0
3WIVHQR7B3LjeRhP3ZrO5FzhHzAeedAoc0kKt4gOOatC6cvGN9eF04DYBl5wnRQAllqrFyboPdjL
rc+asUyrvI5aM1OFUMLzygZFTlEeQ0l9iCyzLaXGGIij3RoD7nQznRoBveTBzd+5U3FOKZxls7Gz
plfBVYmoMsVaE9ekNWO0EpiAjj4NevdlThWthKvRQRvGl2yKF9eFX6nLgX7DselpJikXOYHxTZND
XQTeXKLX9qAO02HB0T0sLD5DvH2zOXheMfbppGZmzozsmnvt4wfGvTY436jdjdVQuPRQHs7jTEnW
2JviyKod9ccow9j4j7HOioYYdH4eY/2npy7ylgmlvUPCWIwKF8nYjfLY7H3dj1JbChYGvSaxIJdu
HBwsFGDRDEMergOo4Hyl7p6CvrhRzyj7jQP/RSa2Ai1IDHyV/ayrp2Mh84+bFEFsLMMI0X9MEG0Z
qHEbalnPbPOsmbeb15YU9X2YQ2wn3zMKdZHcfm9bSTmdX1k6uqLJYD9uLl9q3ttIojP8tk7QkcA2
DXw021LgLrKESx7yFRZMifu2UU7FNnqks4NeRq6Cqk2+bjb4d5blJJxKFT3mbcN2qXjdbgI27qaf
fSUSVVHvWRLG9gIgoKBzW0qQ2rbLzavX2bydg3/cO0vhCBv+jtzSYENgSsJe97n8zAoZBVRps9l3
oNcPBL3pXrw7UNTK76p2PdF6XGezeHmxfZRCBEQn4mIBuXaPWk2e077hYzOE0zsbA8uVQjEj/1h2
UzXApV1Ga7wY0rl5s83lmj8vd3LReUqpiHpDVz4MU9epSDytJ/lLAL4G4+jQksGjtQ+VAV1a9R7f
qdwlYMR/p/L5bOyoQAW+dhCV4s0FGs5dKxPAOzmQWTkFzFm8K/sIUGDA1RYAf/i1jEnh/bsmplKf
WmtCDT1gswx+oot27joiQ8sAGLEwlsHOpzzGXbG/FdFxLzBgu7oqJGYVSxf8axqJ2frrXpKxEcUF
wdYlYjAs2UKJ2KWesX/5z8ncqoWIhKXwefrxXn8uw9GuRQGpbGcoSkxhIEBHueASR8NKPFDtP/rV
F6vy/6pRw/xuS1NIho5a4V7tovMrVL+BeKVykf5M8FWvhltYTIjdlJimTAg6zYUM1k2pF7L81N1+
g6rZIc5lukhNIFjxRsPrNLAoRwxI1YsAl733IDyDbSIx1GTh58vSRhrO1cx/U4VDhlGfZczzV7I5
tjDxhQiWSJZM6B9EtGkXqbMkP6Uf7Zr9UlgXD6GkiUBqgbRUGWevWdcRL9R8MqzgCHz/BJM4nxjy
ENXKQ8AuKyqYRoXM72rJuWa4QLaJGRdxeJ/0UTY/EOWio7Z8Zf6woi+XvqWtJY+AmLsfhpYyZkWx
yuqp38Hh/whouTpJ0967YnXyhY2zUlgmVsrrINCfwggnw7j2kG+2mNPcxba/+niyv1p6U3sMQZkw
7BgFdp95MedTZO/X2BTcig7SarP10159QYTv+rZPPGrthX5KX/ADpJ7bwrvV+GY4ZeKAG3uBm0iy
O4EwJWJEXxP69/MNJgO5xxRuCpvtuWVJ8oosizUHGQkj7DxuYyqCrWwZJbJCF6H8HQX/IQ+PS9mE
q8oYw9BF+R8FR3A5KYSXonuAAOKkfZHlttVpegbSLRgfFT3FyoIT0CCQdnRY7mqGkkoUEuUHE24h
/DkoJXbP+zB9yZwJrj1VC68kxdWYgfGM1kTzlAFzdYeHya8Ozf8iB+NvTLISbP91yyPCGormVlWN
yJAx08tJwKanT80gU4fASSrpFbsPt4cAy1JTmG94uC2K920nEUcN23qIxhqBEpbXWYIAE185MclX
wVjKD5vpkFH9beyL9we1Q2vtHx6xEw422/QlOZpogF9bEYDUyvaa2g3/6qOA/dR24y8qLqNJ8J60
9j2DmI6hXAoojyriX3le5DjgxFAnR0oZBJDL/M+nVgL5Ig0cjznzkLBCxPWG8P3SWA9qbSThuNZm
jhoPtWaro+P3e8w2pfiUty5yEWknadJ3s9HhvO2kb4kGzyKP2of5wDxalur+RIHjupa0UAq+4yOt
yWzvq27q5H2JKW4Mjezcj9QatLd9eIX5/yLwePXGvyEwcIQCcTQyc7u6k21anYGeyuzqjaiNkuPz
IMcINNLK+CWR8t/H2hI6YnUPSaQ3SXksrmDbo6rqSAQXLEKsLFTHh9dK2N40oC7FxXRO2/RHiGFf
lHoqLmltoyicPyHLX6sXbdftjBzzhJnd0k4ktzc1uKko6JkggOC/6c6Tfe5xb54t7l76XgnOLv0p
nBBfqo/EQG0+5X7gGxQkWyS1W9eaBJKOTS5tbX0UCuJ/mF7GQtTjJ0H/1EJBs+x38yXQM7b5A6UU
sfWIva66Sv59vmukk1VILJazGPuWlvBtXZUqQw9mAHGs+PHRCCMbF/1OFxFM4thZnvvKjVm3Szxj
BC/qw24dLKM368zXjrGA3rUUCBR4FIq8Q5IabHtjGcv0wEqCOuTd1PPyF+Ceylqi5Q6pb3E7c/CQ
ZXHFVnugkjqYWWPpKNdhtK7j3V6rcLGDi964SbW33w17BJgLjVZ7z2nMPz1GmogKQtWP9smQ2TFe
uQo8bu9MPrd56Y9LmgdrTozEHzbvhK1NBJk6mwU4QwWzxuShYuufCgjmPYnMi/I13IiFnuVgqNp9
Wbyb5gYOn9n1Ox0qKVZjn6WM+FziHaYGwFaMgof+sK9SeJ0Ik3gTk7EJ69PF7cpcx0z4qskF47nl
vryg+C6XPRr/+aszr5U59vajCVDMhAhr4RgPrhOuJ4aZnqM704E4xrni1VbnPhZZcQSdfH4UKzgj
KDNqR81K0BcJwxHTr5q6OftROdwibeeV2YP53R6eDWHzfdRV8F9S1pEZK7kvwpb1atkdfeSD2N01
YuwJWqlXmFfHXm7hTwdu+Kytbm5GsO/6xEzYwLgCGm7TtK4LcFT9Qx99WXMwcE3igTOWy7Gtb0fC
sE0g8RLlCUSO1m6p1HjktzeLsHip6Xb1EfdxHTgYR189k0fZbPU96pynRAi5UlXjaavjkdCH07Mm
Wtw81Sq2PdgIntAiwwaiLEepRFIWwP+2uMhyf+qO3AIa1IpIMxeyfzcAw0UWohecP/P7ZZCY+sMU
0cHctNmfVeJVNSitSOL0IjvSYG0GUUkJwKEypqsttIxinmOjosVFN1ScbuUdM6tCQKj5r9V0iw8L
KS+/HLUimW/OpuSLuH7WN4C06tk9tMn9GHzYLsLfURbPLZKkJDiGuBtOCVdvEpm0snngbfZ1Zgc3
CGb+YS7KNNON1AsVxmnQJMdiiYM/XMMCghEGSCmrQNVrJHPn1F/jEHJvkvC3BY4ifKTo611VKCWt
Yjn/+EKoJ1fsnIfKIqXXsHFluxfPusyzlD8rEZsPKioPlwMbKor1UMCQPNS5C2jnPc/zj/A2Pu4J
v5kdFcEfdiEiaAWwFTB79MFpjjp1CNWcRrw6gj9d3uInmNlgSF2eElWrozJdiSrQFZTnCp3dn2+U
7VhvMB5NXaG1inrXP51MdoUCPd298UrCUrRCccFR+thNLVfMDwYDZQgG3fNpmjeDrHQgxIlNZfCf
Gp3xafE9tnFtfEHtpjOfgyNYP+wlZC5M4AnbeLGNhmvORsjmIVj9NpoA6zWVwQOo5leYdIJwfGQw
eHd62ug1k4PWnmwvuW6ea0hl0JrkcIaP67kA3DCuAlpDJY8vf4b1eZbfSJHIGydo25q7tmLEmYBR
a5Qwl5/puiTC84xYo5b/PtpWCSDO3Am8JeKsUjgF6edLVefHZsg+WVhLcAT9KQoaEiJExDMQCQCf
ztjicXj91l+IYxas/7qKl7HgJ938fzFoLMrhs3rXwrYK/7U5if1/T0zvGNiA4iWAaKZSZEE9scac
oGRa0pxYjIFjJxDEqAppiVV0WxsaL5EbAIw/fuk4cfYJTUqoQRc9sWz4LA7EkFo5S+4lWCRaIaCe
Vu5qDA9jjuxgDqwYgutgGcBk4GWffSCu3K+Hh03VrcMLD2c/249WSc0h81P9I/m+tYJjSxk5F+8F
e2Xnr4NG9H1aIlFu+MwuDiAW6yasMCoHk4i9NC5jjrn1jmMkQjSjQU8FuKnoEnOOw48/00cYFkLU
xFVEDmy4We+mnaAam+JR1Ql8J8GkmkL4x9VToA+uNAQkcZl9STesyOaNd6ZDjyLh9JlqRk8PZKC0
1kf16l26skY/HRXgwSWRqU9foudsK1vXQKlBVCgZSstPHnDnjChuhIES2ioK9uB0ER29gM3E1voX
SUOBiMLB+t+qH74vh0OmBTzonkQyPbT9A05K8/Hm72Hs0e/fDm0Q8PqtOU3vSvAzYAzO67GB1Aqi
198sqFdEV8kuBzJOh9CyPwFTEgYjxQDrcUkKbKVmrSH9AZmKwbcpwjJ2uJuVJ8QuaJqVGWr8xcn8
CxJgfOWPl3mxLhqSshnEaxYXRtQpa8CKchy1uSIRGnG2qzvfzjRHLN+K5ig8ELa06Uj4EKZriiUC
m2Fcuaump8ImkkZetHRnHh8XV10lOfwwqQTixQnSlz/JT2FyyDbYvY4zEBXkdPif68I5eO7sDIIi
+YzAJ+WA/qP/ODI7bs9A8oAaBGgst3wOSCLfYN5aaMEI0wh84QALpXlkdSBAvYl5aZH3VR7GExt0
LeW3j5BoXIblTtIEtucSPeDA74dH+6+w4YlJKUpUetoAcM5U/Seyv9pom5V1/fCfb4klquXxBRZm
tuzJHSBpOwnH2V1bqZveK9B5CKr9vEQsHL6EVFos3gHkHOvYqcMgz1zQ0Z4q12Rxnij/nwhF4gaH
S7nslj66rChOd4tfwtrhzw2k0qYO44m/B8o+kQbOsAP7TX0hD0BUEMLOH8MyqLw4qKhvgAcLQ2Uz
DlP0QIq98yyF6gmO+o9NhIF9lpWvaXAjSdJGxl3d3eJs1J2eA2MJLkK+hQCK96zm905RIsHQaT8A
l1YZ+FUQP+yyh43AXGFVBomo1rsWX/GqAy+LmGOOB510bZ+pAcNjgJLgTk3OjZeL7vCZr0o6vC+T
A4tC612bch2sX3PDwGKMY6Y9F3L9geqeAsPxNQjOkDvAJfEN+w/mM2jWSDw8U/ab6vp8P6et8DWq
fC1RjwVUQL+EJAXh3ugip+VMyHaYfIBbr0FcMOTPKEy1qHlQe8l+miAIC8e/2I8SMDXHQno7I4Rb
7jdZ0PU1GAi379KcWHoH1bMQdbj332cD5E4tPPzmL5G5Lm3ah7VtxMIza40W9A4qTQ53V8Ai1kVY
zN/oQXysIOaCcsLweFak0NKUrqWFD/fkJiVQQ3VhtPMvF8cdVVhng2hwz08n5ouFpXDH0v0YJRXF
KiE6Q0IVxSNepJvP9ZZF8xOZfJGWwRMQ8hYBfprKR4sKusZFisGw2FV+7V2NWBUp3ylDQcb7/ijw
NqUV9eGEzc6dwRi2AyAQ3ebbsKzAOUNrB54dtZ8nOqHSbhlX8+5mJD8gyWmFuayLPoEbIMAXf8s5
ra+hQDAwToBXJWXLjkQqHvtVxdc+6bM8wPMmDwe+t0dwKXg2y4z49nCsxqow1kMo86UzJP9p+Hw3
dYZb0Hmjn81hRlXcHEFPxGH5YKKKz8q1TpZVved3E90s/o0xEp5JegWRH/lMmQu6iu1+h+ICNPgH
Ja1tTojF5T/ZNU4DLQ0oJbxkWEYLilNUVPq0cJEPhCbv5UvAsFCEywFR6nLyFG1VHp7V7t439nNv
6JrmRcxYeVURb52mHxEQ1vczONN+w+0fJyCE6uHXhNYyw+DAdrO5nMCBwWCn20ISVEn+6Mhok1ab
40gyNvNvLPisF1AVKAIEyVf8pMv+xV1KlRyTcytYBmrxmoNvwvp4jk3DVu3sXdv2P1BQ36si6JWb
rX3WYN9Ok+x6bJIIVUCxcdbuZPQYhBHm8lpuQU9vQFiElEZyQXbyVbvbFM6Om48xY1Lr44OtxswI
iW26AugXTD5tQdiMiwaAnEIeXIZE8S6/ofT/pITlKq2dqJ+uzEQsTXSPgKPh+iUbwyGpFcR4Chpy
0Nik5WvksbwvDkRnOm3ldgBK8Xj3nIhPqRfcj0rB0q8XHhaYSu8QY4tTM7vmnqG1QTrNDCjlSvrs
ZkinN06b6LYXQbzVm5aZBo/wRGFNYt9sz/ebBJDRlf3sg+HBVXa555CcEPtzOczEtrPCK8jXC3O1
x6vHDYjO9Qu4U3sDbvTVDyh6M6/yn1VK8zEovy8fpaCnqmwNzTrPIceBVDNh464KPMe79+r5AmkN
D3iZS4TqvfqrBXKaA3GxGabpINa1E1/sDw+Mh6KvJQfHdvA3J8+Q35kIeWe3B0tIuA660X3WME55
SKjpLpsE2eFzjRwidDU13oM0w197OWyhlTD1abisXmb6CZRl0/fKLJ292igB38SKdt2DyzwSpzxE
apLNHIIjFcdkF2uhlvC+Ds1QhMiv3fuxSrZp/4EERGnMWyKv9uEyLsZR/RAKSZ7u/MwjbA9cXMbv
GJg2t1E0lyd83/IbWxcpWJvZX2TMe7oKrTTAt6G5o8XqCq+cJjLkKLUznyO0P0lwhAcVUNXxelh0
uGrOwZ1Rc2VBpQ/zU0jD0lRdJ11KJA7qbcHGMhE3LxFGAvS9i6aehWYRF8yp7z1ge5tayd64sig6
TLCoOsM26dvx52cgvj58loLVYy7ahWK9pGDb3St0IFsKpU3jZl6eZY48JwR4X3WPieNrPuAdLj+Z
yeRPk3g3/aE0BHtBiXOIHnnLJdF4O26RPI2WXUX8hNmDtwMdNCQBXR+Ot72yX5dY4lZaMisP44Zk
2MAKowhTW0n0EdOY2f14KjcOmGXSETs0MjoWjit47sTVOdOygTj4cLp0Fjc0+GxdOtOUG1awd5hz
OFrF5IsJeYSN6gKHVyJMyGXPkwBz8s+0Oc8/k0YU4u1gmyH18sKwb5A2AowqOHMKfZyCN01WQT9s
1ayFdhKn+nwYizPH6UTTXkwaT46YgD8FYXdft7U4/OCsNHtuUJSEpcOdHeMZF1iBxcfhsqjzE/FB
qPhkPza3r7Bsp3ICuGfzpxJpfc8dEhxluRn81YnKtBIYPejT88q6rEEW0+aWYG2lD5br7t9avZ1x
i42oNWbV3KdJGNeXjWeIpCGq56XvkiP1RVYeeqtY5MEhtV9AFQBSdZRf8ugXNG4Hbh9Y6cDttqDo
iAX6s0gpGGAqrmX1g4Hsh7xKBV/A+vXI4ktydnk8hNq9MB2J65dhDSU0OaJCueWxL9dsLYzY4gMy
yezDu+CQXM6eLpvBgkeTlPgGoqKSjlHxVksYgvewkGt2zxawHXRlfSwFg1pV/BgtJ+ee89DOpini
G19j/dJq3qvEc8DQGeuM8wPSxdRAcxjylnL/fg9VuWo9WCMXvCFUF0ZPFech0dWyXJeazMv9okFG
bCrHXtBsoGkcM9eYbtpiwYAHDEGTnQZT1GOwFbuqpdOTh+9Mf7WXHmbEGMYgjNTiI/M+HhBoLXXq
PsLzy4crjuIQNp+aO06TP8PbIsWBoWx59B2fJVWvo8+xuvY8Mwgs5L/YkEsfR/dKPle3JQnXvWgY
EXy2JnkclGPHSSWKWS0+G4Au0kCjO62DcqjD20tab5dwSS8ByQhjPhFDF/9Vy5Romhy3Cw6Cmv29
P3Ous8xCBZMwxjCXYNUY4Qam1MSXbKi9hoScekVOPwGYstABGv042TODiVbVYaz8Njf06u1sBQV4
kl81ZWZny4h8J3e/O620+GOerlTXR1p96zP9wQI33GoJnRVGDnM8Vkqi+GCG3WRcPw2RQKNLqWoS
gTqb2fEU0OnsMkcbJXrpWWs75ef50dqzFuGhoX/pRPBTV48jj89zzUJ6zQQUPYyqlXuHiekLItR+
DStVM6iBsUZC50Z/PcBiHMlIPBC9WqdqRZRCVr8lWKn6rGk4FyA3JY/ojzTure7mn7iqQ86qx66g
D5xRmIF6EAkZQXK98w/Hc/yhZAXaoibeMRqEtKI9yFSOP83gKbx7bbPXIEZbNGw1lD/H9rItyS5Y
DR4JeHMP4ITFQ3vVQPqK86kosbEFMKxnxDXOs633MqMI2wNbcC77yJdYa88f1NGf7Q9Lix65cbN6
QKwwXntJg19zINw3O0bdsttAe2r4/aH5WhVf67OkZhvgNrsAEVIXnyNdTmisnZOt2Icdi/UzDHJ+
9So44gRbke1QxJC/PiL7IxEeW9sy21zcuCQPnG+JX2TJVxMhguSPljLFOw1kQQVrPYtgyw8rKN+M
NbREBiCPXd0ONVkXrw7GGc2rZw6JK+SKs6g2jPHJOdkGOAHhR/WP89j8pYyn7wOpmVhKXbEhjtdU
xtzFVgcH3XGjc6M86ynwB4T+OQwVaGpJIf7YfQ+8+Y8TIMOSZJ8gBW8gjiu26wT38C7qVckg8lvF
P6R0jn4OkUzpCgso12UF7475yEy4ag0UtYXDNdBGLnUx9zVhuPvhZkUTLiXvoMggtfe7RiLeeEy6
ySzDlRoim29A4UoK8oaSe59BAxLkNqVVv9q0/IbeNnK6hXU8UK5d3dw/rSkLbM0dgiElQ8yjInDp
fWUPrzpkyNh7dSLaqZff+w7oI965/DxuylmVy00jR03lzO+AWueIeDTyfL1cFTqLJhhYSfAdLIZm
t/uN9fEqNX3b30NVR+AyYXboJfpMXv4iPceUmKA0ff7YaSj0iTjC3t3W4pkqXUhfIy0lJhyfaS99
HiMMwpWlD07huj7TcWmGJjLykT44Y8acNWfaK9v193Qaor27CsDNg6BtWrunFE8xNmelJ66AswyS
dFpw/UfsFtccM5yZJm9Z05/xWTOwLQhDu06FdFU0tWr0m1dPxPqfBLxOmfJiNU+BX4wbR68ZAgZ8
m/Xzsm1Mgowm7uat16XtEYKzv5QeBWKmUI96VkSIva1PTCgl7vrM6bZCRjZTeSLj8qbzKgnyTI/U
BWIUdK4ASvl4lGUkA2RXfhJ/5XQ5DpM+pRu6wFNrsAD2dj9Tt91Ug+UF3hBh4cqgibxdC/i0qJ3y
BvlAdO+BbtpR+mUVhudW+5+d1nvZtHmbNRpud2imlKtgEmx/gahjI+kvn98AkixT1Jdj5UIqjj6K
ip2br3B6BFRh2aFWBTjLMsnr+iWzXMAgHT+N/spNx63UmcaX08pE5A+t6NXgkZ6RnYAduht/TYkB
7pb1adXyldIMZFvNPGBFi8pIZO1/v2CKkcmSiSAln3+tIebeIizSxEsaFWsoect7Pq7E2IrFcCJ8
PEYeuI3F7E3iatEQ3MhV1Jp+M6+cvK1zuOLnsoa4cNVqbymQddWeWwhiQ3IPULi2uw6FC5m4NKXb
lXSnam+yZT3WPxaaj5bJvDRwZy0Gke8OwJvic9gmiwQMSRdTr+TxTeVWbT6QUyeAmZOjlF+ZHg1X
ju2mhkLpc5lz5N7NLA6P4LGpXouZzRggjqN07ktgC97xPna+mEdY59wKfTuD0YplOpA2eQf7FFP5
T0RJzURIJruWIeICKzJQAYzDrkDZ/+dvKag1NAjJWUxEDkO9VsvFBKs8j0AD2BIGt/h5O9pc+BwQ
rPCzQXWNIWd2tf428GiDVKG1XRYkrsZmfQuOgLK8PK3ivxh983mljIM0rSX1IBYArr7KxkSypfR2
ZLO3ZlMvJ09gyqSsrhQaHZtMcWJNh+2JCR83CZGOXbUUMfZlqdyBMrTFymhV39MO1JiOtSJ7FSom
VDIMW7KlZ+Ev9p1/ugPilkMTbH5FDYzAPFUDE7rHoOOg+MkLl50a5ANjuGaxdDuG2Vx+3bBGh4Yd
UY9fUVax7YSCCSkGHovofsmaAIRUe40G7qZOtjQfP3ZK4s638YK9BI5hfSCyFnmB5VilXiU9WBCH
A4Bb+022sit6gg2VJKHpc8BQ+avIZoJgIMOOS65PqyCiPT1hDG0tNvgv8km+ceB+NOWLCQcWhsbC
exi8va6c9K6Ms40VZ2qnOzTN+18SZ2TF2/u+42EL42WJIXGC1ktOF+UBPgHk4rz2b9eZi+xp/Xoj
IgYl1RDdSRc5w8I2dR/iiTy+aIw3vNKnnkTB8x5gGDO6LzSafFixfHZ7BFO8JPIzN2IzM+87oMmm
Ax9zyYBb69LHgaFaoJQmrEmG/LMB2dwTCM2GssC2VouDrsZ3nKkoikLgMYeo4Yxl3mbNxGIeXJ9K
gQYmImNDHgYp8sh3MmVHT68EUh/441J4SuXN2jA+MGYOtGDVy5lTkqn8pWlE5mWCvfouLC3rHWdQ
eodjR2mkLcfLKixsepQidd3mpGI2Y1ews1503T/3Y5EnZ/xgNQQrnqh6T3aX76vPAjPoyKYyjnEu
iNCpq7VP2phHNAVGGpoBjXaQlFO9/gUSirwW7e7fheq+6aAcI8oRjTH1oQWsW61LJnClVRApl9P6
UNe7vZkaRCSTriEMQuJkkBY+byS34mOWATTsbXOlRYPn+IDOMQN/ToSMFjpPMlR6rVjwTAy9iFr6
lKqG9981exvU+vGu9wW0KMTiiREq5AluBLkM9PdS6o6Fzgk7UotZub0lUHoj3qmATO8zyCtYI8U0
FAFPOdyW4Z4OSpdbNtuh8mU0FC6wZ6y3ORkcH4LnYakariBPhekkxeInwIRT08YOKZgyXxbhFjxn
/bwcYUXQhuWzObQYtPfDgTK2qe5Lea3nUxQzEl1YZ7riE9gLq5Nm++MRRqdSklBarXS0M1OEKX0+
VpsLuog4EV5s8r5KGX5fxwcucqCEF3cSa+Wmpalfx3p5VlIqh/z8UEt+lnTigaHU4qu2aQ3Dy5OY
VBLfhaGxLrmYmjkwL3iEU2ez8VRDUqkbinoh5sLlxCyofc4wY3CoCsnf/gZUxANOHNmSHa6RQBos
LfBtlbVazwtDmQmbJYewsWca/lFdxDTfbsXC1MyZ3kNHteQUShhHfzsASwOn7ND3NyjzijOylrBQ
HGsOsJTj5Tg5Oe7w5lvCPauJTeBg8qX5TTSuWdJR0NQq6Bw/+sr14aMxsLXDYhkGwd1JhAa4Px2f
VUJuaK3JvIL+tBmLHG37Bv3k10e/A13DaBbcg6fWs0pCNdtoIk1b2gMZEgcaMFiH16iVbflkx+HF
ZD8FOgF+veTKimX2HGg4Dts2sySWxIFMkbGLON3RFtqCfiZqujg6jh9nfyMK3XSrWbWHOrJ2QRA9
gdpQ+OCUSZ3e70ba1wJJ6R+OnGo4ukr7/ZXFmunO1sL7QzcO9kNOshLK9vdrjCDJivr7w4d9XIbu
4K7pdGreoKYUZOrd/hXGdWDhztzGpNBbvD96gHEpeK7WDl152J9qVLTrWXtZhRcyOpeTtPhYCTCH
UoPtc7DlHqrUEpG5cD77FJekoETxIDCx7Wc17ywhF1w6AOF84roBzml3Q0JZ87OBS2LkU/80jPLM
HnnWzmVq+daL9hirjrIXs2qIvI9CwkcUWFcJFSQFYPQYeOM+lae3yMgYUPIO3SD2CcYi/O9Cu0+H
O0w7q+7TiYlFtllYoBRPyHpcOERqkEtmIBV2Cg2Cmn/PkoLfVOb4k7q9aSSE15bp9KqwIB8fGKZE
GXifC7avJPXrV5PxJcw2k+mTp9yQyFHC4wvk3VAHzWz8DdoXnadirQbr0Oxy+ZHLOjBSVxaG+XL2
bci3mZ5q1YN0L2dUkuVR6S3NJrsLAXceZXW8w5O4D8+VJ+Q7Kylualaw8lrFgx8crTy7K5gJIUbD
G3IfUuPPaeQAYoR+se/ylXqLmkdp+BsH7GLtHs8zEvg+krQjXeTEDsJHACeeFBOmYvQ6XgfqdyE9
vD7MgpSRGky1SVAInIizzoF+0LwJ4rfL8upe1fk72Pf1HDyQladwzLjI1GJZIfZavK/YByamYNlI
+foBsbGK00dZtCr1lYTFovEtVixxndaPHs9ORKAZjhWlmqX/zlxvlcuEUrInhm16qidkrFPda7PW
tFUoiqCv4vj9Nkp4h5KO1xRbQD8n+RWiE+3Bh6W+h/Z5v1g9vu8GahBoNdWkEXdSIJIDRuNO1R8E
5GjA6zSlJmNSTqzpU69FGQGRIftaGnEFczWrFZKmXGHWKzOrmz4y1QJB/17YCTc1t9G176Bfdhwl
tREMkowNKN9sGjCslm/uQN/6fLJ/l0wB7x2VZc5RFGhdIdM+fjpnhTmvKNvYlsjHkiSCoEgdOfCz
qS85nni3CXKWlmHIxkxAN/VlUZuNI9PkCJkmHX9lZHFH1BZXbRMMkUttmE1dh56oZOWWmix7tMEf
0OrM4oweSqmXzUKCl44wEzzd0je0ZMupREejtWwqikQXnFbWqir9samZCBfKPAPiKOleBq6zt+ju
qP9poW/RAD7v7HFtZ+B2bs1aZXQ6A4lWEwFwSJ/6ksRM9Y66TDRpzpHG0Ku2X2/+8WXN9Fnd9o/t
aR679MwZWZmS3ysCGkNbPq5ILXCpObw0qNekbNAh78eHBSEBoCRDQzP7gw/Gr7zp+A+Tzg8t3/FM
7hHrvMsn5ewWs0mEqu/SnCvjCg33qAoNnURpbHRmOXKYGjTcajBnv5NUvp6zXHgJ3qp7y783jDkp
GTzbzQVtnPUUfU+MkBMfqQ2Rv0XlVgFIfXjYiEOBTticlZsLDAyp8XL5pReVzH25DpETyO4S2gnx
cs1C8XrO6tnZNSPReclSulEE+kplqMyLLLm4YTIlsITRwm3VFDpBx9vaI/F0dJaTt+/1AjcXNCOt
mRhhy2RPKtK92tYFVjQbUK0VpAan9B9ccStZZBv+xyxx33BHIYHSE1lhm41BSq69KqhRNS5qj3zK
hotnwt51uJDImlKXgy3iUo8yGygQDtxuZp5LSSmy9A1QzT7L50CjvzgLkXMZy9aNFw4MGEeLDD9k
UzyBkS2T/85dYsLUbmUO8VFaKH8bTNCCwQx0KViLm304RgK61R3+0VEaA4paqDvss5tyEGxdc1qm
pc9vjbQpeHzodKD1RDXuPo5HkoTi2TQT4S0G9PI6zL1VGxcbNpPgjhh2LNJFUaFGxabTzus7aD9l
Gsw+IzVhSOqXSdEm4x0dkAEj2kgXVafP/DxQGpaZgc80hDBAlp0IZgeGtzLne8KX8+B1YWdi3nGP
FeFFgnhdfnB9Mqwjmn0Oqqi6sttK/a6q/IbBQkj31rS6wix72inXR0abH8+8uKp7gycVU+Ij6its
WedXpJVxW2eBGsauPoPgOxgrP98/T0aCDw/Z8cWNiQvD/5Tj82R9U1r5LlE7gLpFPaly+A3fnznh
7fnD/ATpUvOD5fBj7W6SXhFPOoD/1GDs8vHbqWduH0u7r4ffsqZ7BV4thSppHts16YB0BXYpL7Sg
8D//qTuh2SxmkD2YsQt4tY/T7qh6ib+VG5ZQpGfkrW9Yx7Tl3HJnl4yG3vlaiLpIRL8kM3SpyVMS
UgXN41v4xNBv9QTduaDU8alQd2cGAk1+3hXWBvh95yvogg9gPGsBXFlMIfUx9mGN5QY97bL46Lwq
QSyK4mvSQZc1cRd7e0Xx1BG1L9MCLgUhYdI6X+Orsn+EHKm2CX4tLkny98CZtf5m0Yrr2bGDgkXS
iINfcM+bJhNTPuug2h+inyuc46zMYCoYb2qxUOgsWUW7aAMbtOtP2szIky/ekcPRSrPvTiW/t2gs
k+EskMo1WeWZHQRgMeRrV2+uAbGdohVMSfw9dM99dJ+pOezcertktC30bOlssdzF5ia6+VRYCiZI
gu2F9AOeiFeIgyRTD/MUF6eoaDkZ6zYE52J/aRK/eGSU2V9GFvNC8tKIyqZ1oeXATmqwsXmovm0l
BPQqwouMSh7q50sZ/KPVxw/NoO02S9jDLRlp3muc+RIYY1oFspmYNSHJ4xXyLI/kc5P7EnQAIlyB
YFFE00sVoUm0dHm6VZw6yy5H7WVfFJnQnJny3HHr5Et+XurfwAvKOUbJ1HEiprwXd0j9B1wEPX8v
M9yM1t4Fdsh9JSBVYzd5oKv9FQKes32VdkoPsBmUZI0nPvS8NuT34zYwOcjotwRbELRIfgdUnQPC
Jm+c2XJSzVLBatPShzuloqneA2eCc6gjzWhLFA+57rPACX5vLkh7lzwzvExEEsLxt2ceud69wERW
f/Ftdh5jCzZoaXqfRZ30O6q0HSj+Hq9DoQIzCJonSAn//v9AjK6kZhqBvKwPB+MUJ+4Y1mMcKuj1
QTlCik0fDXYF69ICGnRd6RJ88WPvrYlvA5Wu4BnOVm+NExCGhuES1w/3MBUjqUvjvfkaV16pBNUS
pZn/Ed3wS8mr+ypu2SadXiR23w81m4WF4E6QSke5e6ll5tD2Xl410tqPBCASp0iUMhM3MVFzQ/Ya
72dBqwA5oBDHdn0dVMfuSzedr93QkC8BJdzu0uSS8mul/wKxtk0wRwCEcYng3BaZLHbbghQoLb8O
lIHpU6wTOYoAmyRCyL92uUihKIgQpeCPTDYZMAo7bpVr4AoTc1Ops8XWYwtaZHfuTyPYvcG/CCfd
yQv07myhT3HA+2MJcA/S3sJtsWQIdJVGroTXIcot+ILTlWWeKjFC030QVzp3dyqQ14lNfboSveBI
HufTb4tbdtcK5GM9lchzv9MGEH195gYHHpzWve+Y6Y2nLftcRur5TfOr5p1by+L0Q9M7IYVXusI8
4AwBk7cbvXpa0Ik18kr/6lVoirRtkgI6zKCAojkDgmrvGAtwRrvz3wuoE69csGfp1kHdV1eyYM0J
k0DxdMfy3qQy1+f7OXb3bhPT1DQdKbAMzdBvIdBU7I1VQthXKYjeKxyno1a+tPhlK4GM4emV5wdy
7PLRIKuaXbwXuc0W8snHPE9v0zC9Ab35ds93XwKA5GBpkPsKB8pckcPhwiWUKyv609wdPoovmbvv
gF1DoXORPLyNx9PZP1LqkYjGWDehbBcZAWCtTjD3P5SjINdV+JCyvy4DcVARctBpUNMNgNPQaQ4a
r9F+2qVWTMFhPYbobu8uFUkL/iRAfU8NM+Xo0ANH4qE+WM+5vb9An+9mdMNeR9D4WYurir8OUREG
MWvpOAHLl2aimD37YvnaJOs2Nnl6QldACg+glc8l3c+Jr/L4Y84HA/oyfYhGKwEr/a5r4w2m10BD
q9BlkjZiZiWNFtwkXa5/ds9ULLTMiOdHnzUS+JM79q7CoEHG66Odv9qL0KjrZbraBwkpswDOeutL
Z7c4ltpafgg1jaDuMntu+Z5HuphsKJwPUU3SIKwmWi0FMANrWL6tmdDOZBm1FphJp8vGVPyY91xD
2ZzzkNkLnDBn0xOtNLv6b879fSSzycLxujj4NWGl8PWor4ztriT+iWNAbyh+906P5leJtl7uTZJn
R4WD1e2Kv59Oy98AnESrL5rXgKBl3rcQXlb7e2HQeGqQCj1EYAvYhmo34kmHmgBkAaZ8xk2QA8GF
DJYIZh+FCMwiGRDVJh5wdyDD49k5vLAMGC2HGXy1WbMsJY0ON25ewuhVmn937CdnEO7fBUJKojaK
TWSfO2pYp2syWcy0O9Puj/+HZ4PJVfgyvLEdekezawT+XpRZEgMbmn1EtfpeqZvP+wdfNrDfAJw6
2BrKWFQgkE0y9smyHTU+S/gACJSJNeuzP4Z7J/lKe9vm5XHrpTjQKtTrJqTxY3RhPPD2wIp6ZfvA
FVcN9ue+l6VH3NeyI8uQkWS/PCgKIbfQwxDPDsOX+NRMbfdl5huQ+AjLbMqCOaK1AAKrGhXYI5ah
u4ElPNB0EaDBtB8K+cDMf0qhDdVjR1UgDJmQVlSpdh5P0EGvRPi86H1wN9wSGxjnvzxRbRHwCviE
KXHA/LXpVXcwYj+wz35LEqomQohBIaBZzRbei/58LHkSBkcBmEO0B0+n0bCIbMbhq7OK7Ixl7dQo
ogyv2VE1M7xfcae9jRQL0hyWhDyrFAD9NNki2HI2fMRo8xn+jq4M3sqwPvbDGinTkER4qruyyp62
NVligU92UV2vh5RmbC1xnOYwgBs/SUF5F5+oTwm/tE+Nlu4cppaypTzZJBLVwSIVluNAeYILlUW2
S2U4gI034SF1t/VKyzkF/Hsu6X6PIsZh8t3c+2iJv5doJi2e7G+Z1jsMW9PXswPUcuRjhceIo8DN
myVnnZfxWNabzb0HydB69IzpiGWOdD8G6YpV9RY8VKiazEGckeMdOh4D9BnQwWhnTy67wb+5XzMS
ZdkUjmAbgVQyVi51P5wNuL6YTeEiVVaplmY3A6lJYUXWx85eEuqZayN3I0oxIRmuNsUYMA1WK+Kh
9xb+98U+wKsPxyKfU2rlSFGxXZmmnC8STsU5MetG9OmUOC62c9CtEpY/YQNkHMRhbcotmy5WYb8L
uGkk37xGaxiuI+yMX/J6vz4RqufAr/m6HiCGecAOm5e58G/ghw4r2j4/ksiUcj0H5PljUyb5IBpl
eloFADc70aCAY8QfbUQ7TJv8BMaP3UmZDhCeCahQX92rW+QXHDjVWRxfTHh/9t4W99Ufi1U1MWRN
do1q1haHAhsHPKDGuDXtbuGVMrWAJchbd6gI1IRA5M3dLG/AEuUqsK9GFS66UdOLpEZQHiyVggu6
EyuXJjm/T/hPlXehePbrcO4mdJLuVCwJkvv5YKK/c6RcItTFtjgcIsYzsBN71FfCcgIgGqmWLmmK
VZLheL0MfYzTXqo8YDM4fZTbvnEOcn0KcACM9VUeu/OtNPbcpn1Edarx20Gv3IdAnoyhC+I9uzqS
RzdvrldLzeohNylwNDiISHUlRrURPINC0V2/NhfcCylOOryn10S1bV42pssF4bYLxKkNiWlloG7f
NJiak5tstQGnCvAE6iApIyzWeRlqAZmEkRxW8bD0GKupRQIo8y745amRZLLJ0AO8fxVy7JAdvmSZ
DCqJFW1Ad1BYdCOpFzo6ZkPRnaZYmrGadoQRVUCqbJ1mLJKndr9PjMxEv43s314QJYe5v6s+NHI5
vS3VP1BKKT0Jy0pw5bcgswBO2+bceRt25jkSvJoi47B31LArw3BM7XgOMpe6Ecq1D39K+JAw9L0r
eyzre4UE2P6jW/IWaaGEuIBFWzWKIIYjLC16qbWHbrXqdO2TcLi6Bs7OG7V80ucLcGEbpOpdkBtg
aNKunnG+J4kH+jhw53Aykivgm4UfAUnNBajScpWi7tlP0hybgSQOnV7dEKvJz6t0FATdwK49rK9t
rJ925acsKBGJYUT7xoc4HCtHoWDhVy4TlL3VScHoSdlZyOOcKV9h8b4DbytSz11OQr4VP1ftIU/g
YwVv7bBrtSaKhXObRzhb+NWt4bsvO2F4gnaSA2hWztKkkXdfB2yEG+yy6krtySlG30EoOfFtcdch
5pQv7/A4Sx111ogrmCZLNNLl9QrZbzF1U+60UHKbSheH6tsX2S4HKWBmLts3g/EO5sq6FBtgz1LJ
QWJpcYi63YE6c+l+3HjcfbSJ/4Ir5csQ/RWNY9W9IjJolvqZUgkqktus6oRXChGEvigNLqODfp7/
JQ4joqZJKEquNNFZuC4P3GleFfQXz9RKCE6ZySPerww/PAXZGPO8fPFlb1c5QTFFChdYy7txQYsB
/XVi+F728WDwiVlQRA2YZTPc7/Znr1PSamEdNr1Qtwu3UOV5WIlWXujC2LWL1dBioABJPlNfPlAh
GSYDbIo+y+SfkvBHHadhXGSE3kEZTRRVwnLBnsEhVjBePPKMFUAeSEQ2zeVwvoFYeBd/osnjGXFQ
M2KhIHHXWBfuUntcZKGd8z/zbAz2USEnjMC+dLAHZi3kp0hmljdBklnPUnGFkHmJBmIHH0tFTqnO
8BifmhiA6mvkQ+y4b9pexLeUAnr+FYQqcxT+loQ/yWUtloEVgI3yBZ6HujatwWt1NtBghzT1CTn4
ZwRb5euXD9HeoiJk6hyjQNlHRJRP0ZYP4oaCQ0R+2TBOr+DO+6EfT5bcfBj9kOg5QRYnKbq2VBiq
lXE4J7CY+V1Mq2C5vANF3JSu7MPNSn/509P10vXnl3sJp41R4BlItIgwsmVcpnSN1eBRTMcko5eF
EG5XLws2M2aO+zjUHECEnDNyZ0sRnE9Frd4n9QfyCyBEME1ylUfCkiD5rN8UswFDUN2r5/Trm3XP
1u5GRQO4lvSGtTHjrje5459caUinCpU3VnPcId9Lq3bg/2uIzc04dGoiIXeQRdL/8I/fKx2ch7I9
nvdWPvdMONspClbLKa3Ev5so/QJ5+3N8EUgVjoNXc+W6SS9pFOufvu9Ymoo1JX2dp7tvfE1SoPPV
f3SY84B4GF6l6xhQCmRjdmex7YMJZR2Lf9xLE4zib2fK+5IGvljx+wxb6Y0lD32Qoya1kwD2CSey
AqyEzcvh2OioQ2l0gt9x0rKNwk4FFElt+9QI8jio+bZ4H/2bwY5d3EFzei4Dus98lLBamNjQbBck
TJVuietH+4Aihb70yyXYuOghAbOfabCyC+EVPI6SA90JCYzBquQh2CK07JhgAorDKEwzb4FnuXLF
m7JwEc5RTYs5xCUg7M4BZb1ZOO29Lz/fd2zVB7mMsDVhpdefsAkibTd5J/xTnMBX6/G8mp1L94vX
L/wv7xWr4MJkjIFjjBTo9sooX2sdT4VTiqEnzFRM2eT5cgZ9GFr474oMBgXMqjS5lHMetuEHqw/4
n6Sn/qqS7S4U44ULvGu9JJJuZIitV3ShPSAocLiJgVVinpDeAyNh9ZijoBUGZtqepCdYCvasbXuB
PpIadd67/u1CkMfdvxRPus22+kv9/3lFIvF661lvXEhpvPQb7grClYdy763O5i7mgZF3fsnqga4C
vRuAMESukf6LuivpgRoT+OKD17QjA47mkW0c8fstCjzJNkTVgcWG8OWADmb5OP9jIXud0upjG3pE
SHzmdopdIEEa+RwFu3u9Pb/PVoTvVjUQ0d68myPZUlfUvdSArronMgiP6GzPkaKjbZ4Zeposols5
HSAFhy7eZ41NHEeeZ59U5+ZSuouuZB7oex8emmO3I18b3xHtXvXpJeQpI63pLM2O4sQloDvwcIJN
MgStQQKYwKgwbtb2lR+b7Qw4Zl3kTkr7f3oBsL46UnHXHcsh9vyRDiZR4bdcJtSRct7CK2vMw2tg
MEBI1WcUOBbfr5k54gnLtwUEDbnJ23XSjBgREdqAMMipAp7LHa42G+qWqYqZ4oTSE0piPXGWWtCy
pKXzOKB5eo6ZDwFVDOMR0luIt0/Btkq1psNvKeCpZ4HkQRoZFFy/QKQpSKSxUuPTZ67frQmE/OyQ
kUwTf2pNG0GdVxyg9VvA3P8TxPhHi+HrydKDo9zgNj3VsH5rIA/xwG8UnOenohjgE9gZdqrcRz5p
6LR0BknE1eDgtA0eFAlBS5d8+n7VOHInQgWI0Cn2yVCQHzFTu7a45gBC5OUOKRLlL4M1Aw4MAKv3
lwrIJBKlYUbkkgT+wBvQxxC+7HsSfxMnPqVNnojdoHH2pXCbOOTX4kFvShjiGNkaj1yZ1K9TB64V
Jl1ifYRt3C4Gqrcps9hMb4l2zRnkscooeB9dLNuEZdEXQDDgqRH0U2owqz9ZAGNrdTGASGXS1aY2
Uz2S2DxkiDthMqqYS70S6fDGsSDTDRALS8Oq4CF0VREW7i3rCaDq6i3AC78frmw6UKqNGDNoL/7G
qE006fKx8Mb05wodiDW8VE45FUCxO0Fc9GjHqtKnySp82ysJZZiQYYHZW+wFtGqYXnBnCu9iku0O
ryAwwWw55Hnsmk9miEGNPUrdTSWULk9F8l1fl3Tb+K2NgPbs12sHoFT2kcKyVPYNoRURucj4QCHv
x+hMghAhf86tktyj2rJV4yNrmuSdL3bqErB/aEGHO2FnaNbecdUdJJOsON84J1IV01LXU0QHyasm
k5Zvs+oiBv+Q8oTwADf0gnjf+kXMUzflEc/OKE8JD32MCA+zSxTGVUPpDw/rcW0l4I/brBeB5u/S
Cykf6ikK3Ag6a+3vYz9ljVauqy/fXnu/PkdPrCExUtTazzv+Xzl5ppZh+ljSls6bTPXLCwBxV+aF
FTnnF08PQotrSGUGTVHbmIygEgWifkGzQJBFQRx/ZmEd8aYCmQfWLKC83WPuE/DVHBzDjo0elK6e
WPvJnfsmKKxUrw1VMR0arFobkVLzGihsA1fG4t+4IAPl2BgA7ZJAJ7ZnaeDwzGXqUTUDGkEG4cJr
/PtWy5X7XKOdEwmJTvCJwvAMGfYHOC0Ke0p+JI+mg5LgwjmT0HUNFxa04yxJ5xVDzJJRR4rD5EmB
iUNx6F3YiG3SF3N2wlRbncVbwYZO5yoJ59PQn/I364bGUXGyPMbWzt1usdwXbUDa4iof+tft1EEh
X04nrx5+9AbR335DRvnaQTDMQIzz49MF0RmCaR43HuxyBf6Gh9h7Sdbue/y3w29RiPGZ1BbkX6Yv
qwh2qC6lidOTa+AxvkDE+RVkKpld4heksM4SwscgzlXs8mNCZxXNwHYJvbh5kJHpW5ePtlD3Iu33
gOPnIMM1U3lMCAQEY/2VCgEBRdYSulNwAJT9spRIq91eRcOecLwMlc1Unt2NvbGmp7keH6fwzsu2
0MZVFPj00LNnq4oA9uzoH0L3BonMHEqOCUOmki54g41oTdiyCVdM2fL4hLrglVeW+XQyM3s3wg85
z6uVwMaThhJIy/fSRVMIzjR2P6UtzqJMuLhlYQ16dxv4QDMfyUHyadnMCu/Eps0a3IGezxJ5Ud9v
D6n1bRbnQVpH/FhixZbhpc4dGzYe9joqWiGc1edDbn0e1sT/3C5sCNW+Q2P6VtDfrnmKe8tasa1R
Tjp5sbDo/adoGow6LV0Bxvx33k+JRtc7WK6lWmT5kPwWFLqolxPAIExfJQvr224mLBlvwYUtYCdx
1BtcLIBoGPjGCvO2uxXF9pVdePJ1Q4R94XhXQmAH/6FtW943XpZf/JEqTXuB/UYYzevlUGvbYxDW
26Yj9LP6BHxlucTEMi8g3jrjBGuk95pcNbm2KMTsrbKkq4TFZxG29wNPfIVhqDEocBQ3fkIXj1Jp
SwJRbujC1iH9fWOkaBkefvxBAmk/OPseScY77vTPtwE5gde0Nz0z8qBm/KCyEtz/ltiopAMBl/xv
eN9hTjyEn5twrGskfLrugN18KJ32jZ2MpFbdX12LhmFH6PflXxqRMIiel/JPd3MjfzCxvqEhXnlK
NLaW06Mw51/jmH+WXSfzFTayA5S/v491P9KO2GUCj/wMVqO+cQpJh2fGuGop7FEl37VT6qKFwmv3
IGwbo0uenVR/FgWxxfSvQw3vbrDJ3D5QuRV+ipcO9yOSRe/MP5+9AcLXHnNEvuDCKAWJuyMQl3nc
q47mlIw4QpBsB4+p7RTGOVJAnTBBO4fPLrdNk261oWIXgFnDmFNwKIhmUi6fAVzkWaEoVRxvzdZd
1gyrUN3ZU58kQqaR3Tl8W9GNDJPMtK98mLTCcQPv3P/VbohXsPPrvA7DLYl1J48OMGSrJD1p40um
4fZM6I+SLgfknIkug95GN+dTUQJxzyC5/rncuLVeSyhnAWbS1UBhsP9OsqVb0M8mQgsxYyYHEvnQ
DXQRqCmR63M5+5oGeuA787Vyq2NmD9Q5ApcS/tXBpJVvsjhddtGYgiCY7PkCRKhpIrSoFxcSKThm
abNHJzmUZ5dS9oZLc1Ymaw8jnQQoRlG+dSF8KpmCHlmEeAC8pmhv/cTOnrvyzC8vo0ICgMBkTxGf
ZE/AuLK4l9ZtXbUAVG+ufoiV5GjMLhjswPvAiApZ76F93KvA7S47CE1ZaCWWjyFIzeaKM1iScxWR
nC3MLMe0ugW3YolNWuSiRoiTi+XDwCPL7/GbVCL253K2kZ0cMZFFJKoWgHMUr3D+ylQeuvTk0JIf
v7jR8UuM9UM5rUGy/5OWddSFW7y0friVVLWmG3VNbTbe1DhaYtOoHpAHpHXyJ+jEmnc5lpOzG+Y7
/ldW+OfSpwBXutiqqBfQWK+zqhZuXbAcNlmOq1vb0K9lOrX0w+7A7rEdUzSf0LCfV0Ff+m036lqS
zM37ofPG545JYp/kPJ6D1GJ6fVjWCdvkZ1Rm8JIXP75UWtgLqDovOQehUSTH89xDdMpp1pfNRo5F
2mdj1Fe6NHHaBA6WGquYXfEvEA4QJqY/R+lVLcSZuQeGfH54Aq750hTsO0YcbZllABzp96/yZ5y5
zLKi15yp7xl4EL8vVDPMV2nMkan0e3qEdZaw5o+66xd+QCtaMlCfmHyKaGWQx3dyggszGL1pv/hO
H7TzT9OhF8pXUaJZc5/SvvPXB4YxjDJRSjG/+Vb6R664zdVUA/e2QFpx1vw52GUAqMy/qrYqVNed
n8+b/vnnGvWBcqvDY4wFpMCfuXyqSNHg568YV5Q8gPSxa4oi4Wo5YstrI1F/cyTbGxTk9FjgPm1g
c1arq7XE9mh8thFDoWUSGK9retYXt/SsBmWAw6CdkWJSOr2mpU3+9tJbekOgYQhgumo3AtFfJfam
iTSMfYJ//8UwVpuuIWJy9mx+ld9o7/3JJT8y+bwWYLqiBWvp+vomWFyJE5l5R5rsLsbujO3tMzBd
adytYB/69WkVTEclg2nR//6JO+aQWEJri7Q57DqvnUjwEM3zXVlUOu5V0RBvIa4OD+RlX214lB84
BmJVWD2TieFGP+HK5qqDaC1TxrImZOLon2PbraF1uR5LUcJptf0bKpWwVIYHkw1Ad++kCq4ctBj/
E5PaAASo3EquzEdCf8/jcGVZgoSPiHzIk/lcGOBvfqa5XJSOwWtUnUsp5tapnrcYUqg58S57kglq
bHLJ8NXrqylu8IiAlvhPbOwDYKXMw146504gFzMqF6lSocquwQbvzQJUyGb5bQ0ikfkGkrn5qQLH
Wm9LAeCWn55NXI6qPxW4noQKHXBvVhQt/umdznTC3jL7O0RP2U24EHqDWD/HGDYImJq/g6MMFqxf
oxm3VFbbfHt7ZwXEk690up39xFm1e30Unc3BOwZn17g7rG0LBX6ONtr5tlH8wHnFRHM3Y0Tf1Bqz
LZuXeCNM9HLfJQMAPMK6RI+JIdH2sprsV5CKl4MHmqxiCj+WQIKWDlOtnEr0hCcahsnSPl0myoWW
C/585LK/yGYOYp53fl1mu3UWoEBCXECzAhERK+/Yn2KZ9S0PPHHndNp2cZH8nDsgreUVxGQ1tIrq
BYiKNHsRKDdBqQODr+2KCmLmTT/ws97Qg7YH2/fQ5KX+UyB7A3AQA2l0sMBs7fLgBrwT8x7Z+k0L
hN8pnTeWEvYcc1gGtgQ7sGCVqG+iGB5/l28nzps5RGfYDsH5jGL5WXV8vjynsfW4fZYkHpY+agQ/
tLJkGRq/91t+QEI4XaHZZ9oy7si1+5WAfuF76HSNLMbOk1A8jdlg9oae64jgry24KUc+ZzZc1gkk
qMMB/l+N2SbhsabzX2AaBEq8t4/sKTF4jCCzBAGHuWtC8Mpn4z73YzWEexv0wQgDjRIKXlEFuy8C
YLT665usxvBXvOgaFVt+WgtPGb8C/O0FPV5Rre6s/YMfL0yICdQFNkAt9Igw8oKE/ftdGWyvi8LQ
imE12hk8alo2WMjlQolWetvtvufAyN1+EWJKG+/OXjKEks65l/iARHhUU4qvXu9B3UHb8BgGtzCG
NkVpchjnic6gs7ED/dCH1CUp2sUXgqFSzssmhwoHP5KceKmZfgjQ8ogIwEjePfCACazAr+DxpGoq
orDyBXK0K5Oyw+4edd3hTNgAeua2+b3vkWk0EA5chIjsou3PBOsxyPvbSGGjqAsruuzU7hXkLSFU
J9etEyeNkxj9TXB6aekDgElK/odjn1k1MqrqJiEW9v93lob9BYtAZtYrN07yWRqFNSXbwVyXi/4C
Q2pKcmoAWjj2xJRLucgMyQTMRJpggDere08xiJLkm6qtS2p9HERHbR4bzVXTLpeyadu63fqgCVDr
jDqRHf7O1DC/NOZlNzuSrv5ybnq5MNnSNkFoQeaKlNRrEHe/oBZP1HRTtzmg/wP+YmfSKgWWgdGv
9vRKLvzEjKKUoDu+S3Ssr0vMp1vEEztC4YxCJQW8fTMihM5eOqz3mesCQCIh/LpUVdAcVb6+7N2U
mZ+rlebhl2SQIj1gkK057pTC8xSqSavjW7IFu1eMYHa1V/JNCik8O2QYn4b0SXOE63h/7UnPl8RV
KrqdYOOInyHvKVqAA4GA6ytjQArRhW7gjDPkW2Fo7EZ2KvwSWvP3dHSBPN5gbMDjHp/yMscBhfU3
PSSHq/DwKurZv7KeGiGy6LW2wCxvPEedFlRKoHHjtkZ0VRAn+dmfhjfGGvwcTgkTIixLb0Wm9gtW
N+X6WXEOgqxv11N0GtWpUecS0zsHA9xMxsciOZAAk9ee4C/gnjLcvj8hkUD6osaUB1mUXYkWZD5d
cNUNTwy5VHTvNZW0kMNeCU1pP5P4qgkDlIVf9xzJLnR74xy1WzEgd8/jpNclvUI/USH1Zzzf1gkz
IivqMy2798hKPGclun6H4lYgQYTZz46dTcBuo9vkzv6hDnpCr0pTG/ZUeftHyv8xvQNg2r26vNlA
KRg9VmPVCiILsXgrybMSAERAn8adVvxbNrAEx3GtUcwFF0YHFEJNcSZV/v4xg1n/6j207vq1TeX3
uRvj3Yd2zd4RjKT3wt3dMyd57MTN3RgCSpo47l1cork+YT2YctYd/x7rfblcoc2g5djXQ0RipHs1
rpJbZwmZIUwiZtbm2wke0LRNLwz7wQSWmaf4rzzR++7pLhjmFl/VTt/GjJpyACdSrdCz9Y1BN/lh
7NrUuEz1ILPFkOqn2qb+ou6IOZn3MPb1TIPSGrIRtGYg5d/OpOs2soQRO8/bwixhB0hcufIYcm4w
W7YO0nMmhN9dkw7Vh/YPJ1TC/YXgZRFYNjNXxggNijsNVqNHRti0vuFvp9n3gkcKOQms9MEg4eqQ
vekan7HNQ+YkxrXqt1Aq6+nZShLC/ap9UTvxOsdjUSpYswFzDvw6hmg0LD0cWQuY0NOeLRCvEZp+
6c6Xor2HYOYsDS/JIWkNri83p0KPgZYR4oMXchJLUZQBllkNPxJQ+yRRnyn1HX3IwMH0fc91Rnk9
Z9zUZem/+uh1b8VHjN43+H1fMRPKgj8AtzyWxqKT/RwgXE3u962XFvguUUWOUEIbvy+reF/oyFPN
htaZFEd9c0+PoERjSDpVRZtg5QCIhF2uBiuO+q6KpsI23ruBesg4G37/IgQJ3byYs2i9GqRjbvM1
otCCvErYbK8OzKaNIMs/oGlTcAMhPw+qNXSQJaO+Jp5YKBjVTho9N8FoI7sU6kosPfOVR1fO/DHT
J4iev055fuzXO+8bP63e2YmiGI8GiKain9tppnvqrmKlrRnEAvVVniiCE2ss7X8mgqwOpXtZ/EYp
HXiNKfJj6f/6SQ5gG+BMV8V8DXVshSNzadwksqEvu/SMjY7n88bgjpIVaeUC46c+04MQpQCmZ73H
fVUBYtptmjaiIW3vZdMvid9LlVKYM9Pt+de7pRZlg+6iv5sA3DqbzUUvroY7Ya72Rdkc1Uyg22Lk
le1CFn+KBtKPQ6uKCPf07i63/jnyhpot5kwzREKzeZJQVhlzPfga7gt2RT81zJ2cuueD2gF7IVaO
78EAmRS3AwkgwM1TagQeJ4n2mnChvaQKYIXjTB6G1Bqewp5gWi9V3XzTK6opgqEIvJvmqT/Zaghx
Z4dxUDO0ja3CBIYRIkepUWnWSzdGMk69gQJQoeKcuQlxaq+BexbLdt7qlZt56tF1+k8vsh8cXGbY
jzLD4IpFOCMljNvhNcMy5XE77Iq25r3Vcg/90JsGnc3Z2ziYtn5MsnVWHqoK779GyV/9GwpLUAaA
AD+t8+Dulsunt/jK32RwwtBv2uX16iHFxLG9WUnc13BAA7433xoVcMiUBhe/1u0nV8iB1nlWAf2d
akpvgUpLI2xivuxjk9lO9kg+oWD5lT1avr3zygotzKjex+qsqT58rutvIUBUWwN+B9UwEXmNW9yP
uDw+dbg+cJUR23LO92iXsXlTNzWeKpNMUy3cm8tXVpq87y1szfMdZyCWdpG4X3UnshXSpejOSWN3
jB70VW5J9facdJC6s4cMmiGC4AMBTWZ0zrJGZIRSjw6RKGZDZGq2guWQ3qfWCESokLrEWkLICUKd
WOnJOXADxImHgZhbYy8ojM5eoKSGNcmb7GGzZ4KyXpHJcWGP0PFaW/ywk6JqrLEl4slj2dzmWgWa
4TvPPgQx2jLK7BXOZkwGIEDRx9ejKmW8GYuypeXsbj04CdTibE7BBq+bBUduQyjZaPY4JbFTN8IH
ZSTrOW3eGS7BIhGbi7sI+EslphQDA9ACp8SmtWwy8DC+P5tcEBVGyq9hHN8KLdu3DDG27PQcAUhk
hXR8BaXqYRU/B0CVkeExGC7jxik5ZCkMDf8NBtxjgLGureY8lKSRAC9NYmRN2dhcj5KvMKr55EJ0
VvaaOmNZ2HcWG7hKt3mndMtdTR0WUlMkKdcU1MuVyQZCj88ubc8aHVvZDxpzFAOx5YEAK54BJWGa
72W8Aa6xvyhUJlf5y1uEgUMbaAQm7bVInCLm/HqNvMOxUt2AlYGjLT2H0/f7ZOmX8tKUXIjyaXVD
Ga8CIXTJgmrfHP+kGpG3OaIca/Lf7hEAPNSpxFETqZn89uk5NQt7rrSYqUQ3egYtRchuT55zFTdS
4kyNc+12H0TrRA04kb4kHbP4aJVIiUmbHKVrqV1CmsrNV6zKEeYQ5aqqj92AXn/hrNf/l6uH3P95
IPsHE5weOEsfQgfVagxjypqaCS3f4cWwXctC/8Rd4zxPaLGRctpU67OLcJMKCVy/jNigyZBs7C/V
7N/SuK7ecfo/S87kCOrAaEMQ5sVmBNOAI5i+hFpfYOLacLhX8s9lBWYHGTe3vuFkEJej+BmcSd6V
hMdIhgf0lotX42/s/vX1tjNrFVFrKvsbX5oaiLlveVlGBV4KOvWaE1Hn+2ozon9ESTJhyjToBU9b
jE6JL5+XYgLMCNYT8Z/b6fJ9QjrRN5vpMKeFYyyrnMnKe2tsKj6Ql5ac6kxTJCeBF+GOQn2dkEmv
MLHCJgodMP6fsetRuNg9KXIlO5iL/OoRHJ9uB1JP1YsvzHwHzW+g/OXki+JyodXF01NHJxJWhFcN
nu4SDpJ0Z3TGU2xdtDYL0j9TAMTSAh8SFR+JNoZYnYxvmB5LStIcgXaCuppm6umFOHBg7lgaRNWQ
Wpc946rlvUgSKPywhquicQepZXnliMzwOqb+jX7OAm3tU9BMsSbRCplGr5LnCkQdracesTsGbkjd
rt/aKWZJO6oGuSIfSKP3yDZ2ArXbgHzMLsk1xIUj5m+RGjDfHODYENsUevGLsOxRGEybmKBf4RCh
Sb8/2fDwhb/roVEccH8OBjcVxyoIFKjetw0UNzj8zAQzw7KUS8oWX3OAgievZ48x+PUvc3tS+CAK
1r5I4YT3CA4NckK2HOHVCE2RF1VZnEGOnVI0EDWM/PzrFqFn26kvBRz3EiN8PMX1jbb9bBXfW0/M
P7/BtbbOfpNyobi8zcgK/aWVdatYKriGWWBHFyoFFQuC86nuKb5dyS6Mp+YpzZW/Vrzh6vVxGK6b
vkHhj3+cldYoWVh3R9fr2lpZ7SUGlBB0M8Vr1vHoxnacXwBdjtBPprypbqAeO6aIVNJ1vw2bhBtj
BtTNdMz7WpZYF6YyIxC3ZkXEGU0xl1K6cKeeg4Ow+QavM6PnFpfkQ6cVNBEuMe07ZRvckRXf9JJK
gD/UlJA/JLhVhlDmjII9kVlSqmrhO6TrwqEQ6Rx6szrY2Zn1HU6OYoOBL0vMCIUr4GG1XE4HxonF
V6nO3Sbpj3+iW93VIFEdzA01PF6DshxlM2PkWLzNw49cTnR8IFByMhF+ZoUu9Im5IfOytEUoEGvY
CQq51EsOny7gXKUu7kO9ziRuGbwsBHRwafHgC8TYgqyE/5zMCU408aUCzFsCNBcXoKmD6lvplTyH
/tC5sK5LWLOEoxjzg27CnliS0XuB3HwWhwmRUfP9hzNgdFibw+IVAab4U6JzkkBdGALn4+tr1M2L
7ujuvc1L1VWj/VM/hoM1Nq9guKuRGj70ZGv6n5EkqkU0HDDcWQrSStkO8/hmwnZK7cfskoxHki3C
aei5HJZQQpVPrfa3/07UH13bMdRCtOVyI7PH42IzmY+xXvV0FQ5z5bppkLaSjzFNt/siOwHf3fb3
NOLoYpRyBnB3oBNXKRmf4N44G0KKzo279GMsgFU1OAsGYW69Qx2fGHhrVQ6bIJ/F6F/OJG1xMLAk
CCr0m+pvhJfsw0aLKGrxkVRBw7/iJ+B/jYm/9GSHl5ZLKcQbmvQKQQxFNwOp5EifmWSqaVV2HKy6
ExuxVDxqTgqY4QO7sIbucyiBpHcHNp/E+arRpH+e6Lxgb6s6PpfSBAfKu0E8FLJVRyQMB+Dd3rZ5
2omLPJPjVM8iMXS31vovMJ7tD5KgyQBqZTGjcG9Cw8rzvsvzFUIiS1lBJ2FttI5xgnwPkSmrqrNA
5vcKFdxUIvCCDZkbnST/2YRMaCCrL6bNHRi2RbLAuoKAxjk+OZbiMu28BTLqWzCiUiz8gvN5g8kG
JGZsK4KXZg+QaHEmPFXaaZmksXGChel32Y9+k7lXfjFIXJ3NNpiLDevB57bFW8U0etiWhItvF4Pc
cD0Jby4+gk377XW0csOhHttd1LylAfp+wzMjWWtTJRIsWvcOZ31I0qY4OjytsyHDEeJvQ2d1a2wJ
hnQAjvCrYAZ5dTyilQdCJ2d/kY4eAyLhVirqx7cFxr7Q1EfJ42ajeUVvwQbfDnX/8d5blQtyKHsi
g+zB0aEtTUfqYlW9ck9CBIYgdUw4KsGCO0npCEM/grLjgTeMlfUkKNuaAGu31651LYdjgDx4AyJi
ktfQHIGcdugQf7cQEmU1rDIs0QGBK7G22nCZLTfag2PVORAbSZWGZ3upvKLhUZW+IcZgyi6tBzwY
nL+UGxD46p46+ZGf3Q6tQO/S+OLUxCehIgIlCGs9FHCSjCXhuWCj6rpEyt6XqSMNCN0NzSyniCE4
PqvH1JVOL95uNx5NnUVKwfBf9j8+imutTZaNkFEefrBSQwxx/jPnlMLPhx1r3B38klHA8RcK/hJ4
fNvVq0g91dkdYPEpBPaRhx0eK8lGhxZbpOAw9EuuXy6pLDogypRrv5phEbGncH5RPc6YN10RN8Dk
mYSOr2MZQcdLm4swXaKhs9eizs5xN6u7OIwQBQgj0dJBPMklGg1SawfbOIRuydmXF33nMAcy9HE8
rcjnIE3vxZZWp7ET2ztQ+ZNj45HLYNGCknIM4o8mO/V0xb0bKizyiLtbQtpfzb3D4ZFQLqYkA+IW
nn5pG6rA6q1iZGYOqrl6ciBX5pdnU9/RfUC/qOH6YzLgdP7I5ezL0UVNtx1IZ5JZ7i38cJYD0gwu
qiq/S4rzyzsUTQDgYAK+/lvfeMZzG0SCHlNlXf7NBAwKSLxSj0W2qbxlTnsscZ8Isxktp6Yx8AUW
ei4OD1N7TIbcUrg2mHFzHfC3d19s5b6RIPsaUk44Oz2MuClYh7m/HnKlScJg2voSqV+lQGvz4Hy9
alSmpYXgL1IA0HF2eKZVRHXuPbPCmDibsKwhUzzH486MkkOhTsEC1qGVHOf+27d9SdiszhfmCsBr
sLmf4lbLPnPwxnlFzcZVPNWMLfuj4YEjXSCWeCAepwq/WDQDX1D6r/rbUK5frGpArwGsfk30lmCT
Q7QRSRusHrqoEx5qRxVkimvNGndtdZXtbxrMr5WVSI9SJ6LIx8UMBMzRuB+AaDMUQz0YNfNjeYXw
JtJZiElYV4N/2rcHJC6YsW1CjIWTcbaPOghKZPYStaxCnq/60eCPOIiVZlshpgIfqzknXDY4Ddt/
vTyyXQc10XEkwfRwo66mUwi8Hd38wa2njJVpnDSEjXx0x22ZaH6AGqfT01l8mGXlQSM/411VRwL5
+Smeesyj5b84WLL7T+AJCZqsXcbbVdppS5sqeBaCuKN8J6S5sxrqk7B6JIcF3kTYZGzjkW8pkNGe
oyO4uqt6GvE68Q7fZx7NlYTaDzQBh+0pR3Epgheck0xao9DzCjHohioDu5yV3OXz02dWSyo8802D
MGuvOcKISjYm2x3kwvewg5lQl118OR2SPJWrdrxb36zTjajLam+fPxQ7g9nmY11u6WkwW9cqqh9c
F59vogKCrEuULQXWGmjbiDiH2mF4nnwZfJY+m86I3vXRigADLWze4bzNYdXTMCHJfLLfxkPUugjg
u9evNvTrl5mt1CdwmOWG4HuMvoVH33t2IXYmv8pO3HAxut3QDhzRdxmshC1nQOlGK95RuQ7ztoPP
/np9YCJ9iNIFNJXOpnnGkQtC/rpS9HTLl7AzAFiEx1oR2x9PLKJN7Vxbj0//FO7YBIGa2NVQ2Eo+
D3+4VRCVgGtPACm5TeAlcbirfv9zLfjyybCsxjnSWNB1qVvASBeAlGWUAFpjVQRnUB+K+8Apv8zp
h+y6h7yN9TueoVMpnoGBuSZllx9wKi5XrrDnVc4af6jY1DDANSvzdpMP970mRNsv7W1BQZbs7/if
dLpcA06U7NUTtV0Z5bTAB+wpx44vUYFNci0jxBexrrSDpULaZZ0nbm7gjQKCyFXfC0H7UDjQXi2s
NRtB/sEu5XzHc87Fu0PLlo8wiWSnj0OIojuX2w3i05qZ6T+9Cp6pKvzk5tvOKxsjm4OzFKaeyuHN
3ynvVSM5yD54DZ9WDfu5UVYhamgpIp/iXsy0BqTM7gsOQ6MQxXY1OhlhcVd1IJanTI6dUCVl4sG/
ms++SWs5ASR4jqdUxWZB8CMaldAJj+kt+HloPZHQot6Y3bpJ5oHI+N10jvw2+4EIrB7in2ONufmf
BeVKA2eFVwg5e5NUX21BO8DcZxmdff1YjsrqFoMCYwcnnzmf0oaCK3lrBGL2uVY8jP+rSO4N/nX+
D35f0hSa27A/aJrs1JIy1p6kHkXkYtvP9K7GEw4Le6H6iD5QOBBvd0QUqsjzvqvPDeRCcKqzl9Tj
tjbvtlH5LPkpgTCA/niOZ/awDixtFivwMLzcPIIlw5DRlaCHALfstq+crz3RzSC0C8P5PizVhon3
VeiFdGXBYF0i6h+VPssldnPH19c6Wr5IANtwL+0ypojbqwNjm1oX4j2uhhQriIE7zehIIqMbBzQi
UT1iK7tgcgMQiHLLE3xf9toVLztahXVZAAbvWjaXt4RKE47RKD3T/K0d+QWZ11RcbRbDTSdK5yFD
ETOHBldWWXaghgDoQXT8cDzqF07SYfg5fmT0Lq+Xjsx74SaJJMtnl7Fu7IwyFuOMtWdYBevyCN7z
Bc6EEK69TAY4MmBnw6QNwp1Tf5b9zrmbahgXEWlJNs7jEttXDmMzf2vC9fyYFDJDZqMXEPyuA/IO
mDSaU4vG4S8nayRkYcfilFelkk1X2+bSLUBZQKR7chrjvqVeaUJNw1rOGXln/BBOLfdzy8aNM1+6
8oUImSc4nESa5JsEOBXvAtOk8ev4/CVjtEZuAACYSZ0g9cWMmactooMhiGM9ivJOIEvV7Qumnwyk
8hxR0JOIsoDk9iyh9R2DeMVrbacMISK68cSZpVFHRkfauYrjc3QkOZL6wmG7Q2ysLychBOJN0FCO
djvg3o6XNFl/DLjSfIZvS//Q4vQWtpfphxgztwHPnQIGta1cEFFg7MacC5MHssLvFo8GaCVOVc/i
L7DhW5xjkpLyUzC2BitYmJ3c2fVTa+i+zlJVKxBq9Uor1nUC9PGsXMOwi8pRG1SG1Gyh+/ziT6lY
VOftD/w/4BApJYXItQcIwF9eUmrol1ZZhD+5HcNnjbcR4aP9XHonaKqlghImFhnrNU87MdSokffe
jjZtiUnFib0wkFrG2wQBXZ8/mpxjKHkxbmPCsB6DGeETdSkTvUW82oBDkIUROge5UNP39r0B+dx7
NzW4XqrD6jDbLki3kYCOtRi7cVO83ShpIIvvUSKAWikE8J+pSsmRusw+xt3aDigXGhVXcZEpPcXi
yMmygFfWqTsiOz3fip9Hwg18rEzEwga1PSISsTyMFQqtEG3YK/QZbYeLXZ6JmM16U5szzzf5xwq4
FFwNLLQT0jzs7QoGIBbLpjQBp/eAkZ3Nf9rnsVE7rWzl105W5JUeaG/9+bzNF6HY+rAzsDSUljfR
kwmB8wNneM7rwWeOmNvjqTTpnD2cmDxPp4UIVuYCVvIKS029HE6Wb0peBViT2VD/YJWKm8fk4hZW
KOLsmjZYxMwxxk91CRE5t4gDWLkL6lEbpZPtaJqFW3B+r3a9Uk/SOt3pC0jyxgW3b/mNMXmL//9i
0WXSwUU3M/nPojZomRJTM7MwxYxM/3Kut1IegH3UrMJuSnCTdDx0UPKXD0++nhPonhx9mhq6kpOs
I/2F0dtMJ9Qk02tJjp8Wcgu3zFZigcI03PcZFDbjn6J3wf8HcMVET6NZPPqvYf00JZFwhigQAc4e
fiVRI15fzvZ/ayZljZmItBxHLL2zLiAOYVWzZygAg/UbGgQuGdRQJjrU4wOjVdbiNRP9vpZgOP6A
Bv2ZssaEj5ggUJOziQdT6ZxnUiJAiOzNE0e82JoajTN6Y6/59cnL0NWGAjXwBttxzy+qfMq9hekv
3b8+gYJpcgD7LB3w1N8eBKqa06pZvY7BO3FxO+v6fqSSkTVKfBddNVrcqW7K/Ezpb+OfLY5vdp8X
oLE9eY1GpuncqkGYDPXrz+A9j3wCR73ApRLUJhjyuOep9PCApiRyCXAdXpqBr795XduTkWw3EQhy
kHxLZUqH4EAq3V0pt8gzdRcPzzQ+TdFkOUuWQ6yX/cYj5+v3pdFvZxWliCwvefcOl233L10YMGk2
hThV1HxrzuniRnCTOL/k2y+SIu/nEzazC75SGaJcFLreQo5NF1+/Trj44WWCYQPH1xh0CBhnkX0e
+wWbqwjg0hlZsH77ehcFv4mS3ZZwJQS8ffyMNBVU6Szm94RGxr+j2xX8uCGsudvmRFBtb+V49Y6B
IcCevWyFikQoKXoAY2TqZdqz/AiVntLkONSmyiexlm4f6hz/4vf+HEDf05XkPjauLKdUbeTmzcD5
sN9rdoam0Iof4jcPeRuYrf17pGNboGdgDZWLvtaZaGjNUVjjjDBXHf1h9WEgwolKvKkKZ2SQSJUt
8HWH2jMdEoWDPDySYHs2PhQKbmhXWNq/1EJva2vIgKzlMM7fflSVjIEpn3LAY84C8JiZ1Yp/dIlU
MTPwJFsFoO5j9HtZj6+6wfTANMK1kvtowjprXsIe7C2+z1yZAaDaN7UeVmXz8qUQy09HIm7jk7cf
hvknZoIqQlHcRSD/pltleeWmB7Uk2mkjKACxU45xuu/EP3vLZykhgSzhNPM+VlFzl8xIuBL+VDoX
oaer8YK8ZWwRRf5qUdW7NtQLd1wPrS0evr+LsTCQX1spIXDD2a7dqVyz0hhGZkUhc/OBJwn2VKJy
zy2USNcCEcl7CyQSUJ2szCS9a9CSL30hoUqi4OMdzFAENke/zXDRtE+skBFlHodQKvsWSfEcIWr7
D158y2iRW1PX04yPsz22j3Fdff70JFKePzi/NuDybD/H/gIFseJBcHSLcM6ZAdvlrAABCSZvCVzP
bLxeyHOjIynKrgIn2Es6xp4MLKRuoAccg2vbYZB6oM/E7d+kGYkJlh2Ll2qkpMn9egtCQerUGs/u
kttaiFthhIgYQZ4ycWfUbLZOTZV9FqXuELNJ4xODubzsefRldjYlHpqk/1jDvF3EQwVZqYMUM68K
rtr2h/P4JiA20hBdtPNLG1UbRghaPdJ1hhe8c2SemKBRumukghLYVPTanCy7ixCUdJqM9WH1lxQ4
c7CMr+QaWD6CMVcu/2hMC7YlPr60MATTcwVhuDM9ESiwz1hNnZidOMT+IDjD1/JkGojeNL17ivWK
jDdv80LvD+vA5rOQKH+h83cKEsVOC+0FdOXwGTqc6NNNUvcp2v53XqeHg1bjf7CYWux1xjDYrbys
FhuWcR3c3yvCHbDnfzYV94ficX5OuqXuAec8YJzrFXCffq7t05pofKArh5sTkgldLJoQ+l5jZb9L
5XykdK9erRnqdQ+a6wkJhtzLVJ7bJnPE5JUwsZZTRx8sjzrYforLUv7nMPSJstOemxzMrrR3odod
F7lDfL8yYTt+SQFycGsDwE5ZKo8ggZRXdHAib198+jTe8kFzqzzPuwpj0DkSJD4e1rYFO4BVrseH
eRzkvIOdcrCw2jMWIJ/SdhUTqWwcmBpUW/r3X6R1uto0SzLdoFAlnJDXenE2dB+Q5jxdWRRo9IFe
FloipzPZNzwzmMRrH0YknXvdTxHhkQaAZtXAx5IFgGnZ15YNEiGoA9AK8XEEKNP2w51p1hTanmgY
j6bwimZaX0ooqi/zo5tuVrltYgHiUpT94dGgsujMNfJl5JF6nuB8zoLOCVbU0zBYNPPRx5MgAJ6v
1qAHQ6HVIn88M22kcJc5/3O7DHsJeyNox8yXXS1OmfmCZHpjoSLe1qR3JU5nIueM/RUTDaLwWf3W
i4e2fRZ91YzB2d/VpLzEoN1dP+apkbaoTDg64ttO616RwHxU7kxYKmrtW+sK/0+p0Q+aBrWtZAdD
ZJaaVi1/QpPKbwXlT992/+KW7eXRov3rSniIXcjdFTFTVa5VccDSheUJ+tYK1AfKn4fAI63Y2DSW
MM6W54he5DvfS7unXyMERV1TnXBeB1ntNBDjc4JZ1tegx7Wkw92X626el9Grv/MU+QRBm5lm3gnd
ePGjKcsQe6qGmd6dqCq0vWqnOdlgQx0Du4ZyQ6UMwsFsxTm6gOQZ03/tHbxolySqbC4wW896W8Xl
XX0Rm3hvSCnFT8r0vMIKWnfZym6K7f8T7RkPsv8KOMkn2m9yVspTiAvf7gal6Vrz25qzyj6q3I5O
+oeUq6VzWHdE/Y68M/FAeZQGF8Rtl/pS1QxX/pkrc9Sl84tGQKAHgT/BzuqKJAE2yc2Iypm9qX6l
6tyTPfHJKmzQ3GqYlRBVq+nuWEdV2W1wZmvU+OKTtNvqfz8DZxR+s1rVtJy6KZ0nZIrf5RyEyacQ
rmjPiexyh1aDzM7KNG13XmKhoEHnAnE5Ro3fNkrxhsz6SObs7LzKWz5vQAeh/UC32Oiu+k1lvS0F
PURkjIFhoUVXRfq0lXtH+q/85bTSKI+VAWh6AfYJFv5vRASAhXoSI3wPuxol1tnvImrj1xXgFW4g
odImB/FqUlJgVnhvrs56NOYk6dpAE0CxeZbM8fSGKe6sCSIF+rpWfKKi24ZkmoWJIp6WMcIrLzwM
K3B3ho4RXWlXdOhPEsQcigmswf8FyMDVW3+KUGa+zkfAHcaJXpa7ryd1MBTKyPCWSMtYqBvuwdtD
1D7WAC9qlj+VVf+lccNBHRnNTNNjyk2GGb9zIOWiz9Ej9cS0eHVt/vi7tPYaNtdjpPQpXESOQrWJ
tQ6rNmdKGRliT5DXAjBFGQyxMDbgyJ3kybo9dyoRtVkUYkZxphGcvFi22Pp6/u3KK2E75qXPpkM6
XaEFksr72VFTs1o6XmVv3LPcWkgEuiwO8GZFm9xFyZfb05BOKqPKxJeLWW4iRPK36c9epLQAQtTn
EdovmxyoEskEkCpX6aAYkeQodf4YKBrAlGDefQPyoIpB3mR5pjZtfA3dB0fOf8hXkz844jYoIZgO
lF0NyW9bz9EpfSEj7MIyS2OvA3PWe/DSMLQ5Kq6c7MjJOgS3XNTHR089/DIOZM1DwivBx0z1UKUR
nSSxiMxe7NlTCicu+1JbAsv3y0JUGb1kvZU4Hzu/EKVZomu/WpODkgCzpBvnm9osbO+4LM/1uQp0
fFbA84GO1fXGv8twTqiTEm9QZUUdPSGWOj2/bLTj9Rl0FaT0lsktunGzSzbh8ULhqnmocJoo1scA
j3IaUcN7qU3WCv42iRrzkp02tPBdb6HlQLl/mUyB4hb18T114pnPrrr5I2PD7PRRTjaEoHbOwr0m
1BQc7NzOh4+Ma0vlsX6zf42buqUyx8dc17DrCRhI7wWlOv406gK5AO/o3udE19qbrch+KrUiZfE2
jcoG05qzA+Xs/DY5vNdlvl6X0HJREW4Q6jxJGU0I+h6Rj5wZrK7ZBeZACCYozlYsooS0g6xsnbVt
LgURgzBtCDQ/Fzrh9DXCrzQ8kqlReX8InuXPQlLOX0rQRgZIGEhnnJMP2FrA+EKFrgqi7qVxHx5e
ythY47RmP9LUsiM+/J000FGtkXPtXNzz+MCgEWgIq1l8QaBZNDzMnWgbpVwaq1haJi5q0Y3gKofd
hac482byULU6l+mrFBbM4mSZIHzMufte8SOOJwOxE4TeFZKLmZbm9ZfjUjf//rDb6Ghcm7DCFO5Y
hhRGyA8dEm6GAEm7lpoYz/yOW61aEirfivjkG7MHI2ziaypiW+D6vsD5hd7Nc+b8kqF7r9mHsGMy
9RlPVGcrXq7KXdGXflygMT/wq8+KWyiA0bZQptT9iDs8+kLM/h9z0fyKdTtU6HU0IFIvM490h6aI
/Ji4ISx4COhY4rDqe1aKPRw+FzTjhLOfdbmRWWQJIe+QO3a04xMEiuuDelRI4K0o5uxKvW4zlpBN
sYkjplFf5uRT9YGs/yOc3kEL4QXvhZ1bdZcllQdRjSN2TP+YFaubh/nnoySWb3Wyx4bgzvOF7ZqQ
6brojQbgc7ljglPJp+aZb6oC2gvp2huNdL7rYw2wQmc61tJKE3CngaomZPrasOJ8SI0+7X/2NR3n
xRXij+1Slxyo/om40UnWfqBTQukd3ijsO5XwayaBcCQL77grAqdlyr52hCrHPKEuoV08rff3xb9w
eOg8faZQXYsLyBWmcjvv/tHtISfhMwM/cPbcKVpuksdGMGJZ/YTgc9tjIvXp9hdRF7Ui61TetKnV
mJsEhQ6pnn7oBW9YrCmLRu+7dt/qZN35tMhKnaJYILn2sJdXLT41UCSbk1KMYE4oP+eAGijjvB/R
w2LeLrnjxyExjre9Y2x5qVtCtRFfkoB3Tcx9P07fbfLFjGH2DtUJqMzT70Zsd9ePBFpgy/pjvdGP
D95o09xfzN96vFaNIUi2hZXqyPI2CG9IuXiBolyFsLExMoLrbcy3+jZKs+StbNRW8eajicbX76ut
4vkBJhWOSVUqI3gpbR+SLt/Zo4T/LDYY3La2C9ejhJmZ0l1PCQ3lGPo6t6EzpujFfJHN6VR/yue+
lPR8LPi3FtpKutM4PdOvUlS33fuU/dM3TRjaYqzO9PwZHj1AT173Yn0ascMve6D5bn5Q9Z6Thyyz
f0F+8R0Aop/YvJUR5e5Wc3uXTFiXIZFVYhGeqofT7dRGCMiMXMG5CgTxdOMzzBsBDjaRG5HcD0/P
9WRcNQoMDQsJrjzrsBAZXXSryiw3jCV/VLzwrReCpa0KVHdckEKLgvUq4o7uY6WzEexejVWVutS4
SIwusDq7CldY2UurB0GTbuAuYUim6JsNGGf6Fp90EJ50/Ho82z0KO1SnOLDmX0TqVjfkoNvc5WZW
nojjX+O7rLeIvnKTHzQYjgae7SflOVtwXDGEM9nWbjkBD4je1+JaKRcRgBOZy0Uu0/LT/0yB/ibF
13Rrq1n/JX5IGzO+pz6Vn7+wcxd85ejB+m1UdIJxMJxlEyumfu6x5MoP8s3UprE380YkfLasB/HS
IkzpdSZZAM37QOezgI/wtPAx6u2odtCmc+lLueckf4Ji3WgmIsejZPn3Eqsu/9LKSz1+XOk2pxRQ
Fm95F3d/alzMAtb+k6wnuHwuWDl3sGy/xCPUNA4o7KsdAkGki0d1yZmT3YSgUrX/fBfqxxmIMmnz
fZJXFgN9jhVBNVZc2KxGl/YRX7A7yCqGDFyh4clmsiBwyWCp8khcu0KxmVH75CRaFc9dzTk0YKJL
6yHg01aUnLlWit44yxje2pAjO1PSTBJ8SfjgzrQPw4bF+3sg5Y7O/n+EcTSnpLcYxu02GiuwRs5/
yCfLOOIfPZEMnGBZKeHqvMhHInWc0zhdIz1Wm/kfd1l6cEap4W6k26z23zwVaZct9qYPJHoUxFTa
x+g5bgeMRMs/PkEY4lwiYwp4aj+Nk6SCyVnpM/IhAivzx3Z/qF3dTlpIcRd+RpD6DxGdgib/LkaL
oA1Lt1UE4vI820yHhErOdygsA2GEo21iaex+XBVv+FHPaYBJ99qjqWelPKijDs2uvV0gNsdC2zU6
s97F1TEQTcGMMtlo6ds6uSXC7Tw/EH5aI31GyM+PEhyvv8LKfvhdPKmHwr5c3vLQ+YqEyEarq3NE
AgSIXdyYEJR6mguozcsW35GZ4IqeEUdr5lUlFaImuLg54DMD1WXjTLHi4I/14719Qud1z3KG7OaT
d1qUQBAmfx6CpE7LSWf2eG1Ck5cWMhOjrluUoqnmOg9Q3wVEQUc1r4yEQGWd+mtApRpsA1shzaWF
fKCus1tdtaPDHZOUUu+y68bZpvbr8cH+4RXSDSvv6ce/Ab8lFPYLDL+mTsxjJKWWqomvnHQ5HlTd
SGJrmYGXM+XnmMjN89YAK29Wu9kSyC9ZjDnN5VBYBAHmJAaUvywj2DgssN+7H8pxdcq5ICS69BaU
1m2Isb09jlnJwtis3O6hcO+fRFJmySCiLMyKp/bACUpfE1HPYo6TVgwlcZTDZGc6FxQ7AyWOTBOK
MjgtURDvhZQ04LgxgXO7g6ZSNo/KARHyBrvjFmfU8aabxMSrNxzvCqUwjAMYYwJzJQol7i+F5Xa8
ax19ay+vOEeUdxN3DEJFXOqnKaoqQuetsG7PZrMNcApMcO5Hc40XJMKuIRqfM3ZEmD0ujSdeD+K4
kAFotKokhoL35Vk61RXDvtYnyE1Tohv725wpBNWpcvqgojr//JWZXW/iB9Y2EFRvq01k6ejQpaTV
PvLTpMalnL0qNmYVR+gmpEsruCfEMKcHzphMXqSGEZX/2fWpRSGsoGEmVTH+Xhqim8WdNzFH8V3M
DaQ8IPG4cW62qpcsW9LyMAeINHXJgoTErOE0dM/kvismiRqEqY2UM358Pl67H1mAcVEqVFGLCNY2
JstuKGKuB8TmHFrE3h+SC3FW2JCJHnrYJ5K2KcFuImylcGckRK4Y2cZNrZ52kFqXtqw2uT85Cj8S
JyJoB/NYeNf5pb3JwGc2IL3lUn8fsmZAVuVYZ81WKgvC9FDvYEmDxkT2GpHzG+aomcJatxdgv3EG
vC5N42oGjc0sfslF0JKF2Ij9+QipdsVtDIOMiffPwN6Cna/LTT4i/gKbIMtAAdx4igMEaCiZMt6l
hRG9+Ai9uvrKrC4GcnljaI+DPIds8F0jGWat0WtfLzJ8SCxTIDbEMLQ5F/rn5/UQkQSFOdZHv6Tt
7QDw4X2tdn6gdKFCFApYivHo6qCtsCZQOEUkLh1vmfqIimAiR3ErT0Nn4B8895mOijuSn23+0TUu
x+d6PSzYfbn3BOtJjULix7KEwa/vZwDGj7k4rekXGfonNOikUXx1s8qKRYrM3PPI9NpgGYJHmzX3
Rs5yMBDnEDrGyzyKtNrT/8ivbIqHWxRjPGsuxoe19aYre5yJoloV7uhXW1re8e/VBHr5JT1gyOA7
AicT9HqUh+mp/kS+KJ956hDyEGd0d37I60lZwHkaqPA1YKIBUvhm+hZHPLcPLO7GG5Bwsw0+Ugep
1WugJdC/8h7xdAlklurO6QtvQY+GE7iNycV/k0tzDHYWZSvbDWyP5EDG2NrX5qbt1SKveQiIOmzU
AT1otR+SumzEQOwdQkcezrm7mk566/rMj8YOTvj96e8vg4B9CWDgksb+fICMi7R9aXpCXJDOmeNd
oiLGoIx4UsLeiDpT0omxl1LvwwPwfSNYw7NS5MW9apreqig3e7dQpSy+2ZtKpYZInv8z22WWr8nb
hrz03IKXTxrz9spkT+baz7L2NdDpRfGr19gMug6iT/Cj+LZP2yXTTkCiU6EIE7/QUxroZUJv3Fnw
ocDPNBtWTXscUNaD+pTttNALBI3CoorK6bGZGL9RI5/CHUzuf7tbSPS44JZ9iKGkod5WNqiMyqGV
54GGPFRqb0iFax865oQy4wRrjkNvB4aj2J9JONjffS2YRZaUNLzM4wOg5akVWOIx8F8aZH2tc60v
PlvyHiu5L5QsYwsc87/CEGYJ9DjmTOb3w9mV36vLD32mHGQFPkq7HdC/oBI+NF0vR8YBJ3w2NiDk
WVJH+MEevVFIOCXt/jKPLcBwvXetPsSZxna44tQoNf4sIBf7EQ/Z4mYQeSSrtjl48sL/RxKl1KAN
drPV3KXSLI8m5gu+/L8Oo4O97nrVZjUEN83zJ51yrKiln1RKuJj1/ymWbdGqJjI7//fLpdYegF5w
SBDr1scYzUuTMmvP2GONnolLlpChgcDLdnvebREPQ4iR/QnEX409jJ2qdXt0LUMZIJAvTXQNNxeD
s+17WdTrRoBWGtaopyHFh7OKlimnsbgW4FtMmZrBmukQoEpbdNn0tVCbXiKLyZmNoSULuR08PgfK
/NfWgxDMJ4rRfO339afFA+mNFXmAqYf7zEmwq3dZCpB8/k/6jUEwLmAz9lscSuhy6xTw5og2eqYP
aydWH3L1WWfbE0CbyUihUq0R/B0gkCC2Alm/0lGJXWMfGUngR9VG/kwF0yoHHl12qtkD7gbdv6rg
jwnAxTfAXKVeFFQ/zr2dGsDN5zpOyaLlzQDc4URRGMrllyXBSWu03tQKwQ57HLnKTVpTaUpz/ujO
5amhEBlPGU4bW2VJ3Ul7nQBTzvNkfjjOvzEvViylOv94gFX+JDyXADk+M1Qqpz3K8k4+59Iub0aK
J+UGEj7FNCuj6fQQ6YUggw35rHchDE9+WEOzeeg42nFt9h6TEV6SfOwyW/SQ4BH5jNkMiYViU6KE
lR96JqV0dvKx8zRgLLY+GaCL+PwTY8PvhWnAPtN8PSpb9Ko9z7zWE0cbmO1+TOjv4HVo0GQaBJs5
n3BnsjnxO7zuKp27htgqarDQnquKO2aERp0x+HyYYmKXJcEfXMgN55W3U1ll/YSb1fPfAaZZ473w
bt6sy1eqynfkZPTF/fWNr2Whf9nI+A6lRXr/xLJldXs0WC8xqSykzYrpMTQDrejItZk50azvuGQB
/o90+8kivrX4riD++ieTZw3GQyN2wQyM9W9Ja70zmvvK/QmBHRrSUbFkMO5QDnLqlPg7xI19DHSK
pkhK7ZcEViTS+qsNOXsQl9lWho/kXCFqi6Hk+Lkf/V1Fqy+XmsOCC41jPdCLh9Fber6/ymRglCEm
l+i5YVuDctgbTchugMDHqxtQBTCIlmJiJD01tvGRkSj0qXDyRkAR0aSQMlwoUmk6dqK4jebGfZ1X
2zPyTQnOY12M+Pc0ZX1156koXP778fyyVoS3xR4mkBkuaxneMRcwH7cggut3ZUQaMFYm7iH7H53K
ukHT6S8tF5UMjZHxrI0+CNxKJA+7sVWOzzCpqly04aqzO5aKLgU5wIUlHJ1yRmwIDXSQlaIqhNZD
5yGjH0wlDcwSEpN7X+H7rXxhBJ3vxjhnuKlbk+EQVo5RsGUYgTIdInOL5LlZLGtCw35uXOLqsROL
Rmr09ciZpy/l9htFQHniDMuJc7wwXcoNDXsPyfZrczDkwSpyLx/qsB4K4BL0oVAgeCcBFurv+MBj
CNKdeFvd8Kb6sIjQrpy3BblpY4WFpcECiFUXAICqQVTNdR91L3iE5b/OyTgUEEw0Jt1QGYJjjmcQ
3iQdBa17YAIDNYaM0enpb+6INt/hW0DssYfut9RVYzwMgPOlyVIUBD5BpSDiTWeatrsTpVtazF/2
lwdgIDE9mBQOAU1SS9v0CeJNSAO0xX0hSHy5C4a2Rd/CVDNuQ0x8I51KHV6RkHkv8Miv5Jl6ej6b
/MdnwXvHADEOyJPrCqutJB2tu4iqbqqZrE/lkWx1WKKyYXX7KhqL/UvY+2iOj0rZj65j7ZM8Qi9T
6gnSauuhmbQZQ20cXIzriq+utOsEKIlYOGXbbPPl0hkFoIQQLPzZNfj7oTdPmaKmHd1qz7VxmntJ
wPX4k4hnHPsHYY/4acYHs2nr+GXPDwqGqruBpLhZN0umVHBTDyIlN825ZJaQA+3RXXru87SaKWuZ
ZzvXyV7PiKLe1Q6o0k0izqR7nMZWpOV4JprmV1zYM43sW62yq1IWuGjtMENgDDNyFvxNGshZBBEr
0E33g0IAJ0VxfmrILfZMCRq7zRiwyqQG9y+03JgBbxmW8m6YvaZ232RCPt1q0bNCPwMNAVOgm9Vl
cn+PZ5rYVH9nRdJAgnGqUkyXckggzyvRln9EOy8lNi4DVDyQl+mXXmBxVojRo6PGgtf6xrSW6Oaa
wkupgAeZSvN/qvrOoLfeJCSbCnbIOaDPy/mX+RqoQN3pGMaWsSINcMMv46dYgSHNdy27lZs28Pj1
zO8vav1tX6Aqp5wMuBqJfwYK/zPOuqMHgEkVz/ogaoBK+GD4Apb6UX9eXu1BO1CCa3dwdT3T4Ixm
aU2wKp/fyxdWtoHuMSdXdFMa8xfQXkzgnk8E8IXPboAugMpLzjEYwDPBamxs7/AeSqX+BlqWAKWW
wG7PS6FYbR2tDRqe55G0O+g3jL832E01wtBSN1k7t/RdNFr2fdvOSgGHxEJOwbB6WjSetGOkcZIg
FfZfZGzYAciNzydKjWSzVmWUSKQRgPuBWgUlhx+IfhQfMDW2lx8pEhgKrU7iZzuha/DEjGEY2CaP
owxcgoscgqaeDv+gFcKmyjf85zF3Vzv93XNVA9Jl86nrG3ogDCLp5OSOW/3OlwQnHaJE5j1BfgNV
lYKxvkBbGY5eQmWynCiNDCtuUYmBfAPLalmFpEfk5Fqo1lJIQa5jUp2AHE8pxjQeWQgmhSFJ383Y
WhM5K8+CT5iQjuhOqdffYCEyCXDkjHY0DwZSxuqRwikyZCsbJHx1sAtT8vBpoJ2fqH2NK8CqIDKb
r8tuM8lMmcXCzYoT6WKyS3NT5pK783YJJuRYWgtKPdr+a9GVeKn2VHsb19s6X8ou9u4KeOt2t90R
y6orxKQ2n2QB/lb5XrHJMPDprku4f4xdxSWU8jGls8q1TIkpYsOORCoF4Eifyfvl+GMLcwQ3EiLP
Vpj3KM+00WYqIDzodMs3YOdJ9z5LX5Ra7gbKLBKpCIntXWv9d99+8fbehQQi3biUrdJWl6znzCDx
quiRk/kUKdkgCFNDov5qxIwNq0L6BUK73lRpSuR9YWiqTwx2qVa5FCoaebrU9qzc0UnPoo4Xw2Xl
5dBPQMjjXwiIao7AH6UTgr9WdYvrVK+m8OYbmHxI16kCK1+Fn04/S3xuNwj9Y/g6OsRT/8LK71ea
A1Xiza5AxJAt2F2swUuBrMLvW8vel9j2I0UqlITi0GkV4+lOyJ0eTstVBg9uoPpe7uYQg5Hmawgf
45vRbc/dmOrQk7bA8Epq7qPTqEMVEDGGbnv99reCkRxHfkdhTiZkMeOhMcxu5Iw1CyoN4bKo3AKI
WohUfGYcu9GhnbiZmklmSpXefZlKNF/LK0RaXimxIUH8EL4fdHJ6roe5J7Aw8Y5oY9j2qLKzkdlv
RyWMvlJMK2IzdJhRZzcRBfm+JqoPTrdXzTmMiq9VUIP6cKH+OsxIap5apDSRz+JHOOqTHxeq3Lqa
e34bLveQQAk721j8B7i9ZVOgPOoc96+g+Xg8voQ7NrSyBptICSPK8hXsDXcZQ0S2tPEAbz1SbeTD
8xh1UM6GNSvYZXTgeuzRI/uTSVAIlOigFTjTwlObjkH3zvxMLuDVsVH5SycR1QQny4xg2S471vDH
ixPwY2C3kcndQ5r+RVSur5QjLHPjCo8d04hbWwmZVE4+Sd1NPUY2r2zmj/3wKPq/j38U1/n/2fcL
ZCnhQBVRNp7ugKKb6DlBH8hjLOh31VPn0i2ayr91HMGEkiHICioIxQyss+RWRvbYZn14Hbm9ub0/
y1HEE3k3gZahfkUzBo6QRBaZ+ddYEZ+cdWl+fGJUSe8sSTXzdBWQJHtXd/f5gOM7JP/wAHJohzNH
RI+qZ6v2GOlwfYJd6Gef7VeD4oqPbo2fqhBFdwIUJ0CTu7EWHJEUzdS51DaPRhdzQE7Qg2FsF/Sg
D3eiJ4IpE0nfP+FAoGT7cEmj1B3fIi3k0nFkEyTMFbTNxBMxKuglLdMnGwcyDexSAnk3I1qhReUq
ffhwvgoFe1ZOJKgCuX0ns38VlQL1GAwH9cLZ1lkWb/y/2YvUwmr8mOhthHjL9BD1U+RIiiJ5jmKz
uwxtaywVZlhdauygKNUOt5ZTmPgqViAvrdU1TE0bzkHpBUwEYB0iMJmUa7L2S+qk3PrS8ydkeakU
CJWT03MAjoTTdPcDpzht1QH4WZ3aDGm+a1qieOrsxq6Ju/z3bTKdHkrZHHjcjT2++N6FCzscmu4f
O8hrzaU35lM9SOuVO3/Osr3scnobjI9lVtU+sWyiOyukxYwSFtYEbAXIZNY5nC0brkarCwY1Qk0q
fXDON+kKdwZaPeKd1yMMYaR0Lou6lxc62i8NobZJ1AndW3qt4SPAEpwygvVG9woa0I9NBSMSzaqE
i9rYvx4Uv/Td8wMkgPKKG+PsfHzjGbyn4hp07xLZjA1OLr6WLtbjOj6pICPq9hLuLrMm3ocz3Avu
EJxVP0P5IReFivyfZZgCeJLaFxkOZIcTkk+I4aqJG9eQmBbIc/TcJ07ej8/7CvFhLZP04WmDgGD2
nsgE47Xhgy2QWPfpKY1Yd3VVdp6fvf0huQ90HnJmDq+lA8y5IfI/VLKEcuZhlyEGAeZd/+HbTwl2
x+Ykmlo9IxV2njnk0ziWhJ+NgVdpj4W0F6Udj0FNGDBb8ytxil2j3EBupR9gMTo1vRbtrjQdseiz
EmiPtUVCsLzPAjKemDxgiCjcZSHMgsdgUO2SmrU/1r18dGiN9/qEcsL/4durIQ9MigeDABkJu579
vN5iBtONM49FCpm4BEJw4FZ15ObNXId2eW/yXY9bYAIyv7IV3rkuzZitHAnP9Lo5egfdKSp6TeW+
dFyWe0UUAI2VK3x4btcQi+d2XiELmF0KJWBlQi17MbcYmVwOs/aiFTZeSoY4ChbDiF7A7YdbGbBb
/H3AoKkuVHBIxGqBJiGyVXVQwQ1NA6Kiq8rbgIo3B8dRrqqfDXBlC4GriEbmyC+CdSomNLJfGbQY
1OMbI8ovUGQStKqq4yx3pb0QSRqcu6ArA0v7BOU7ke58If9TtMQFUBOqUab4nMyk326WbWxA+X9a
dlXTsR1qkrzG5p5JSjLRRhAFczb8EAlGEXPMBXnjGfZH8XjpzNeMNBaVxgFX/0TmuaH+bRVCioTE
7GmLXAiYERm8jOlwVY2RiVFWh82m684m0IRi/9hRlNHBQjp7POxyLLDGB04JIL7Vp5B9oy0D0qLi
otmY2rXSHKQ2ASOdxKHGTU1XPIQsOcSG9zIXzgLa0RX8K8KuobAhUbcRUntfY2Fj6AuVhKgiB+6S
R555afKJIB/EeU+T9WR1QtW//9paz4NXz5CV45mOFQnJ0WrBfTq27IK8KQwi8djXu25dw5+3PbHa
3RGqmOuFoKpB5ebxu52tZ2VCZfxqOq7iSWFN691tByIjliJ2nWwfIZLEXhyl6zblkzwNwyaVMXXF
XNIYqyW6Um9VzEVk6PG0G3EdejyRJmuZXM7Om8WDAC553XTXRD8+qQprGU5GB6Z+CMGJhOhHvIq8
SKEEMVDckosD7FDfG8G9YCX7+7pgP50m+cTE+6Gcg6Z8slIDdkExoOSvtCnY993ysrYxJYBCW/eH
EooeEJBcxYyDMT/LIO86FSWRxsfRdmIEkNv82Ns8geAhzdJ8gi27B7JK54GnE5bJ9RuNLQuuxfO/
yz4VXgM+rZF8nLI5UZ/rfXVpUc/kCv8UXaBfEPLv7+Tcx2Zv6XcFjmixfbDULZch+ZL0FuCee2hq
r2xfWg0ZwCkJ7N3G1Dbr7AVOF4iT8FXPkHEh8ek/BbhbK82TpB75T0liVIrA7iQ2kq2GxQVgNicB
J7qFxXwIetudCtkmFGsd+NxGncEiZRZuiXNjK9F6/lfAD8pTO1NCtXNgfh93Q/YA/HUmikiaeKFO
Wi6iM1TjUmM47+ld6mBbY7recBrAkZPkptcRCQTwNkNSPZC03/xBqnCCMZMP0uBH2M9Kmrjr7J1Q
P0Zo99paReU2W1KMnSlrKPu7Lpi4/dSQhGNSR1PPs0GzHJLZ8uoT+YMUFq5omvX0RtL0wU1VDP1Q
2K0NAXYMHQbhcuPn9wUQyTH7eFUDukJ71uWH/ia6JioDuhpj/ZYMhotS6MmVbQzcTRLwYoPNgroW
V6WahUTrbSuclTz5VoJEBelJxz+p5hnuiXeUmNKp5lNT7AKoObN5cEIxUrvoCLX6BMJ+4EmMITbt
sf7ozcUXdlu1xI5epwJ63XuAYyPHFJ2aejySjdo5BOA++JG9Ajq5s5nYQ8mUjT+Fd947xtLP7jj6
Kdn1whWM05+ncBOWQICcTj9evmh7KlrHs8rlJmpGPXOYlYZ0u/sCE7wtCVKUeRRzNOEQvK3RG8VH
5EQ+wWtFdmZ4LeqKREOc/RG79p9UFtVsRutICUATyYjHVN9U/ez0ELrlFUNltCWLTvowlh97pDEX
PHrfuAkVE/rcPeDIqKxLkf9TZMLaWJgGtI/NinmAEwjVoBGPoTQZcnHnCtb7+GhLKCuKycdSYlZX
amwcf1C99cIw2LpAhuZqZS62eb7iCqsZxiL0azXb2LV7wOldtmz1BJxLznbBvPsZyRt0jELiglM6
mjsA/SvQp1wP91IbkJzmVxl0NbU9zuJH9zNJXSJOJC4ilGJtYnqc66VkFz6OX2nJ8xm66DzHe48g
UzL4/hP3O6wPIMo12iCzwPKS4tkGILcHCDOMKFO+AqzxvGmr+Doc6wbXMUOEtAt1yCSIV0KQIvAx
UT7It96VloIOzlIexl0r8CCHDH6wGS9yv06ATMCu6VciZ/nz49L7gg54jkCrKUr/LbQvrthABLps
UkVLzCqeDbSlh+6LD4RzH7GlrMSUkGnMLLQ5UQ+HpcjT9HCvzSMMGR8nk93xD6tn9zoecN5RyoMJ
noi8cmSiPSq9m/01G5ntI8/U+bASkjgegsvrlbb1s6KPbIV+M/dHWMxQeYWavuwZoP5dTwSIZ1KT
OWauPKH3BeHfshfv8iozj7kXkYojm+El5RIlMeU9GRaBdRDXqa0vBeNRuqPXN4UDpwrH30GHEOmO
h2sjpUMPYKqsDy5CtCBw1Gdly22vzqn1vm4ABFEXO32/eE66Tpb0nnAE5+10Rgu4QQR/LA7s8TlQ
IN9CRkNnrgFse6N9sOMGjgrQ/Xi92VhvMtKv7CvaZGGurMY0Vv6wSScd9kHkcQq1KTDLn1KyQEPA
/U4eDnmU+Z2JC+k9xKzZFqcAOzEcQxUIgxDoI9prSGgRCoVp93BcE75rMGcytFQZKN78ku6OPO+Y
E0ZRALViF60oa9KLA/JTFUwvYfSHxjtu8d04VW73JlyquT8EIAtEHQDuJgQNyrRmujtx0SAttZKi
HooREOmkFsRGB1Qx8hJAMXE6S7s1SubyTCQ67esWoiAiKCsevT159O8zoUb5xIYSVdbWdc5XNhnm
5cTk41gcagXw/lzVPKejGHk8F3UE2OnePKTzrtHx8F3Xvm22hnmAgokbdDg9aEpN0ztTZaikklSx
XtgP74qPfqKs85hw4atgUDXHZQom5+JZ7qjjJbEms7tTugGWktJsEGn5qUvZvPgNr7bziYG+kIss
vbV6qYvT8+fpGktHigVFaPnjBuyLD0a4lZVWUU0le8Yd8FA/lnQ9/Dl+vgSkSTMi8YGXH9SADO5l
5q+UU9ByGvwX3OiI/BUY0fCuKET91EoDdg+ooXM9vPjo/kGiKvTtevnSwiZB6wdpAS7yrXFhg3fy
lT+oBpNfQSSvMPLVpL5eOtxXRijx1w4PsBGsRFQFdjN2022MtbHCQn4wUnzk96K4L0K0aEOBCxEx
s+E9/NHWnA9slTdu4mrwCb5r/Dxpuf7B12QrLwDZW4vF1g3E81J8YxdwzJi1gcyrflAJGPZtFLB9
UPcGzCwOyrvVd9x+u3dJr7ULkr7kR7PNArLFSGkc4MrDOACwlTckM1rc3DR9Y5ZNJXlwoc5X18Rt
y92VbPYeCpHSNiibn0N7G4XmUqcwZVqWQIgZOjrKFBYhg40bltIAXI+D0c4jXz3pA0rAN3AtwKKA
J6riX/qu0rWEfyKfGXKV3cFqSLVghnGerZZ52UIjcbaBOh4+6gQLliow1tf9GUr+U/F44am5j156
MYbqki4kkqyTkVqiDY7Nnhn8mIf996IjMy9Lyp2M8Xe8yjHbYP3Q4mTRaNTfLnOgLOrM+ren6+HY
Qtnd2wxgSHAEC3O+se6cc6/G/H9ncf/eRZWaHhDTlCtfXGna4X6BuHR1ymZS2P4sFjwRytmFMHa9
ToD1SZmvVY5SO6QceGncYKqWqgWSewEowQR9UNGlmgdkmOwPB1tp2J2fT+er3bNQ/Hw1UbuNe/NY
xLHqnkbgREKIF60eNSJSHElmnBgHlfU0c4AyYyivDOaWxIk+oonXyC3ubpPYx3UwzK58PdbC4uaz
uJBdG38EGsHwfh39MphZkqTI6bV7PMGxEt9Xiw0NR/Bd5cCZwrJJenDI8kaF9wDqVpqv641tktlC
ajN33ozn7fNmPWXf1K8K+KC2ku1kGLERN6D3PiSBLLqgcGPA9KS5iXYOEMx66AVha8eK2+sUZhDm
44YdD1yeUTg5kdS/aKFt2PM6gpUt1rB6GICRy4D37YkJenwa4oSgVkHe08R+4H1uiACg0IHRzEMJ
yHmRj4stSw+Vlk4F2FEiPYtb2rGWkmlocCMGeOkDzZ8rDas5dH8L538Dwd8xNRuwErOSk0GlUC97
EaIcY8sHeP9tnziKR+4a+Bv75hGR5QxJXesvn7JXZvlo234vRCgzvzHug3S7/FHRghAEd/5fYvbJ
EaXdiofcxt3idzE4nlKIftBXehD1tGmyUbFiqbE2tShXVWn5JS2eKAJsa9N4Bjqp068hKGPlpntF
mWt+hzW2F008rReU5/knxr6Kp4PVs7r0Kw9Y/AOVF+dAb+apMDjUxpA+UBy2KTOQRzXgKSfx3Jkx
OM9optdIWxa8xgyRK46ngo2fHnrGFqGkpwniHsg6hOQAiKBz4yYYzzqNRxRLNJ0i3GQVTgFLRwqk
a2wXriZGTyEr71rtVPpjBkPhHGUm7+gmAya0VtpPb7lpAyeQqT1QONKsdskbOz/N8r48nxuIuZXp
9Z/FRchYEwxIKuwmYQhoLXM6qo/31CJ9VP6MKA+P0ic629qgbf7315TTrNCImRpAzVmy2miCPMKk
MWUexmH1z5BtM7sckT1p2AuYROKRytIpiX4BsLeOh2QK0Dx3ozqaiDUoydRk9gbp2HYiwA7MSdY5
RQ9UZXj7KWCkNFpKQCeY4M6ZrjNyE1lxjNCXEYggk063CRDmwJ0z7Ai5o39GkJzgMggo7dWHJF/O
m108dC1TElPr1aOsDP9Y6fpoH/FEBsnbN6dsLVCyaz+u1OXbtVDtGXmPFEMKX30itzk7bpx5Za02
cuWC5yFgcIGyxkCO2ceo6iIVa4r7XyiLIJbJt7dJcWoAvbZQbbe+IPrxGNjK/Ie2NGE7Oe1dxRbn
6QK0sln5XqgU8P57H2W4oRGUN4GheOh0yJV0k2ULyC2DYA4/DwC4sDkjjWgoFWp7slJEOFESeZ/r
QltZudTWpmbPgIfSHbRqc/Hh0qd/iR4SFMVci4CPUiW7b1of1PBZXv1mH01yD28JPNAuNKSUqBXM
7DvxKWlHXgOICi9yxQij8LHA7TaMPKFnrVXwpJqI5vbvLYCAIVNVU+eJHa2dAwzJiebbXuHZK3EM
Yq4gHJKMTe6Y3M4nzQvhWg2An8n49Tu9JPLyFnHQXv2hNV6L3qvriFif2yNRvJ/qVUzSFMfEMytD
+mOwKsGiUkuDe6W6McTrxlGxVjIy4776qfP8cjJssY30t5ir6iLm3suK3yXgnKeFX+XxyredxaWm
tGFPyAaC+D65W8Q1DLuhpFyassXU4g0/0jmzKd1QGtQubM6Hg7upmw3eP2wZrEBAyAzJdFpskP/O
FZADU+Bl3W1ec8SXEEJ/2vIOnsWPc1Pf2bhklXhnSn+Pj4kq7IPD0u0voqrZ5ahcADv3H6iEIiWX
zlUUYX696b4KOCJ+E4EOBvg02Yww5vFSRexZ2HNIM7rRYxqnCfxDL+wqV5A56wq9ze6W0wycBfeB
H5x27z8EK5CDnQcB90frMM6qtRx+Yd80ExqGVRCZzaXnnmmb3YdJ4KbepjIq+EOPUrBJb+eeYlOJ
hXw6nWSHmrAKpvFfkLsGAtp1rm3gis10C7uy9uaynLINUhiGRMfgCVLTHVRxQa0lba1ZzrZWz9dE
C87ipWMDrOJv6P5oH9OFjZXm9FBXxN/FNCsTaRZoWeRuRf8qAt9KM8foi05AvNq+JUINml8BEIjV
9mAwvycGazuXsCU0ojSndIXQBOXDkveioMvhdZHpI3wNu2BycATo7/BjTcBz3nKSDuh6/1tU5biC
hWqyYoAhrbHpp/cr4yBrUhx7Sq0P96JzSQzkScm7L5VCNTmLVfJ6Yg/82ki0V/NlHGoJks2nlIub
AlDEOMJvmtIwmyln3o6hdVkEt544fw5WLK5EkctED/rY5XrRLXau8So7dCiSno+tv4U+VE1Ec6Jh
QI53nlNqRoNkoBqI3qatD2sK4I9Buvs0E0DJqAO3pN3FvQMNWaDpIndH4tMrmeb0Ozd8rQl91ZDj
OZxUJiDOJm8EodrwtL2VzfAbbz5rjOEQqAJX/3+hZHr1/mS/fpiEz30axzmm14Lg2EK6mXtB4zGg
8bxY555VvzKLA7MQkImK/G/x1T1MFMT/07r/7nhf70WHWfWJx06dci/MgAj5jjHzT5bKPSyq66Q4
XeeMmh3i6tv6KHIRJHGnjnsrABIkk5bvGZeU/sFV7pepTxBvvjNMPBTNTANY9tu42jQ4uskFhlGT
6quQtEMyP4uW/0nr6O9r/zdnUyT9adX1D7Cl11gDauRkSRFzwB1Vlv9rKOR4rlaznQYurytUCIZw
WEzKDhTfUBoxRe7eXgBJx3WflknyCYo1Wo2yIgeawC559AVq6z0/cxXsp4/2I36qICSLY1ZpqVFe
RNjUep00x3TX3e8GGqEvlVs44eltj6bqEi+CPxWP0dib4PubRvvXAot5tQqtMceOmMujQmD8DQEU
3Nsn85op9zTFBWHojaJV94w7qjpzaISTGdcgGZNMYs9uDIbYVmIZfRAb4bPorvLSi0qfBMAEwR3k
YrcULpfwEktRkqLAUytvBJqgXPRqti82ynrR51BO2DmbMb2R+3iExJTtEmyehkX2IAWMVmBkIqg+
+oRVfSJKDp2SsLx46lw1a4zKeb9L/qn4k2wd7CyabCNhxu5WL9JraTNqjjEkj3xj9yAfeDyxn4dg
0gFP+CIPwVtM/4KoP4UQa3S2VoRVaH3zYKls5i41H/NONIrJhnNWagdCWLi8Sy1VUMKXsXDJZGc+
akw30q1R/mlEwlwGBo1VVk+JwKrpipVqB56LKkcoGu1ejksW8Hwu2+u7QNyiwljfoTd3qV2mS26B
c12DYkiEmUxdLbWfwrqVfW5VCZOTDKGYtGjPLEFA9pCSY9+nWayhKkS4/IOcNYUCkDvQ7F0a/KKP
CdhGCIKC00X8Oxlb9rfepnUCsWq3eWV5MSSV5TG24q0w04oocwzQ4t0yVjHJOGNnzsP489TXECYq
TwhZNB2CRC6kNcWAgve7DCjpYH8MwvhTLyK5W4ZoTW2i8denNyZT48KAaILt1I+qb5nkEM/9UGG1
ALjVwYw/A5fUn9hR99HB9kHIiSaGLsZ9GVI54ceAXXU6wipG8rnDRw1mcnQQ42qk8Xcydxka93xJ
Gf3kOvxm51FxN+XETIev42p5SrouMoTIqJHjUbq5cmzBrCZn5omaRu0pXeB5LudXzYnnUhxLEnWV
aUWCJbPmeEitco0fwucRnpgzpFRiRg2oJVm3iikWHVLYGLW6YJ76uu9/l/ItCKaqUIM0IQVm7D+I
0LNbBmJNj4ZjxtjMmG00S3fOllTb8IfpxumYepb+WAUdgs9dd8ImP4J1NrkDfn8UlIzP3AWv2Jdx
Xj/UZAhjuPDDsSjjU8GQMhHkHT38vty57z7Oqr8qOeTIp+XYHowPGIIv6YnU4PQwQxj3wyj/0JAL
LH/1GImhaiXRkHln0zHisyISixY9UgHOdiyhCPZNvtBVgiodeoP4zeDczmDBcT2g5JQeT6EudNyW
T9JAMQqCi3IJQCxqfKPDnrKYhtXxHqr/oSqiYTRieBn/alDPUEHs8hZ9dPPaNiEhkvEtn149HVEh
9uiw9LsTR0diZ5GOgb9jpDfUrabaa+8JtjgrSJnaSiO/L4Ci0W+MY0qEsYNeeKTgorTNueacVfmW
viszxKtBwA5ZZbeTEN2aWUJt7nuHFhESmfMFseEgHlAd2/skS4ZTShPDdiH27TqUtybD5Fak+4oh
RYreEdfdixxwfZpnbhyRpbC3veJhXplMhLru1teSKhjBQ21HRk99XVI3KCugnUHUoJ34papuDDPJ
AANV+C1Lc3RZJuD7HlHNL2fqSIhxfMBPOZtpn5QCarQjML0+allOdBr7NTy2aohlPNh9oV7Vbxxl
L4QA79TerScDn2FJodqMf+GrSOKlbQzhp6jk2XOIB+1S7lImjzo+5BWi3EUZOQRchmPyCIHMI9PI
BJd4RXCZhdqW/GRWyFImA3nQpPuk4O8YWB1Xj7TMk8doUuQE8m6BdhHH3rYL+GLh6pLDi8ob9uPY
2YotUgTYptRGF6clmQDp2nFAU4Z+mhm9KYGjplsR3nboV+ky6T+qvNt230eYfMKQBYV4LyiXQ7sb
Lp0cQqxT2TK9QXb5VLMsT9BAD06VHFjpj3KbvLdt8V7zwLRfPDd8rueP75+k/pOFO9eRjDejDHws
t/tLKdP/MCRH+MIR76QE0q5pmmwgjbMctuSXWm+qCQZKtSZqZNDIC0m4OebkFs/YhnAvsfx0whLB
fTUiNR6KDA6cROrW1EjuVHgSDCJB+QdWYxrXRdrk7Fy06pme5F+2kkUmLtzXVF28MiIr+zpp87pV
S3PoADH8QODm82wd6yjf5MjnIUySn4R7SGXts0GZsOsgshEw82rocvlnZ9V2qcfVU2CXussSWMFA
nQXuKKRpHJSPldGJodVyPSyaJS6hCoVsnnPuwqdtb/mE9lDx4B/Vxz/XgQrdSygvmxph9ycqWFix
vqQ6MxwSzxY8KTq0cSRAJ6U2o7JIsQP5phzMDjBfg+eK3LNRHwmn0fb9mvzNBZcLeCwUTMbA+GPC
avlgstkf1Z0Q7pqF/9BzBUAk3xjQa0F6siVlx8wcSukCJUR/E5Xa0LetK8GhXCMHPPZDMT0s19Rc
zhhSetF+BxEVyOeMBsouXxFVGIxB6uO1yKEDM8dAMbDfaRtG0X7EhQwBYLy30Z4i2um+HV0bukau
sxEAmQhzRBvhaqgJ2Ou+O2TQ21CfQ+537XkmUtA78paBYjeIIQFX9wrQ5EPoK1gf4oNmK2DJ/HO8
wTwNwoU5UchqB+2SWwKrOfWno7+OI+wv3BlSjjuHyV88qOEoX2EOGvR6IeEr6dsEqfW48fRCmEC8
u7hRIlT44jYxxic8IXS/xJ9hLmnhD+NCq7x2R6Yj33tDXDaPp3jnGWJF6vK9kXRKN9NrzvR6hICL
NSF2hYB3hUXqY9OcxWRnPPxB6XPvX4FD6PJLoot82snWURfgPLvCFcZMAprEwqI9WBh6pL3B4iMT
C+v96pWU/Bk706rQ02tIx+59AkdS9fiu0iRHvAVoxhY4QFz5b+3JDwhU61zGGbR852vxJE6G1CAl
AiRf/oQA38FdCfdcRoWayWlr6p15BM0JQYAtEiIJ0FodJhHrTDOR8Sy/w+gPbkSQsLTzeZx9GPX+
ErSF1lBIX1dlZqsf4+ZmbbNfnoFfMuXCGzf/5OTqR0QaUqHdxLyEKdMQwHN3htWpkz7hrjFokDvH
kUnFtD4aoDDGOIg6O+tHg9fYSwdAkQdLnAnOzaQ4nXMZeZVi5EVF8BMjB2z5cykvC4BNjjDZEC+d
Vaa1fIeoC45WLAfu2AVPRde+syXJ1KkUZuB9UjqKI4ShqxAkK4+NzUw0hbMafpq4zZSx4B16cdAV
zrk1lUZg66hW0wya3RRit6iYUN8s+I9tZ5UhVBEimXLgUdgxGUN066X/511lh4pqIrk102+5zkD1
iaRXhWiDybOfjbU2vk1elpddC+qUNYmjM73B5Ikf+ejR/dudc57U6MdneZVDvDWXnPcdVA77O//O
iT2j4VTa8/KA4xhY1Y1mrOXSFajS3nhR564C0THlohWM1bt26a1bBu5KAndACQK7Kc7V0cwkFoWQ
yyJKUZpBOE/4OObYfQvqNmNlgJBm/DPlMzmqLgyhCtzSClJQUJ/eNXrIbTtu83dXkbxq1+Wc0GYH
i1sk0ouon7EoxO/o1vGMSNnCc9SDRsjITciZDRa4app+C6fuEIvmEHbdaefLvBGY+oYCApu/kwnz
cBI1gkZtcyFgfmnzoqfImx1lZjjrMIx4u5eDyewhIYiv7ZfBkDR4Hy19CRuTyqm7cMyij5pLuhKl
LS/fwlbqY/BleKCpnBpXlGC2vKfO0Uo3Jx3XO3s24htP0GPdp8F7XSqlyONY1jdZZCQTN/kaGoow
qmBz+tsJXdmM06w6U6tAsoIQ/8bZnxUAjRdM6LhW+BUlXTIDHRC2PVut+XnU2lWf/Bm3K0T2NCxc
5xAyT6/T4pqQUIDjUCOhEVH6plX0/ApC/p/xG6FPtZ6vq7xQxq2IbBvyRGXZPRzS+9ZPKB4Du1ir
i5+4DzrcIKK3gq2cvF0X8sYaQsk6uBnsriHBpEBIiO8qMIw7qlcUZb/SGcG6dxYp96kq8YZvVY7n
i6LBSHYOr931iTb4foNyEYKZ3pbk6fHz8mW3ioL0sEV8vpYRE2J1ucVP856asvN1r/SxY63syZxN
kxlZkPUoYiNq0rqOt+P7y7qL9+QnKBR3b3AFNt0dWPB1ZiaJtUQXABttRGwJwgtIVkMg3CtALMCd
hY15A6uj0oK8C10+FEwtFeyRY0ZqeloN7SIqEsAXHtyc4ZJ79zuuSvy1QRaLX6JApIUg2t/bGH4A
P21V0fEOAdTi/LqZBt56hWlaed0ZmAMf509NnFidmLQoFTnwjatxK5bw3hvKlkYX/ZckkjoRztE3
oQZWrwytbaEcf++xGXb4v+EdBVDs0o/lfIpF5GS0UJlp4g9KRdXQInCCP1i1GZbzb/ctxejDZBZw
s2IFYqghCgIZKTCCEmVaHhhLgXOQkqNK9+npbxSaWGDB9WfE03QfMqy80UfSNBIVJf8iYppIFmyc
T1bOObtWDVoTZdzeu8A/5D32RUinuFq9L2QKUBRt8yLjXFXPLGcTSKfHOFG69JuQMbbddGs0Gd+J
w/TrDJbe2AlMkmKYLnbAPSga4oNP3GvmVA5q6LdNRu/vKgVYQJrx9FkrBupaJ2Xdg9RB2VkqM88E
/IYEbyMof0a/eVgkRliB8KaoeGP02XWO7eg7OYcsFqrb2vHgLb3Kvcg//itRmo8sbpUFcm5k8tKl
Z1FLvLr2wsWyfZ0BF73fWM7UG0wrUPeT7GMggjpbrnSGy/zyZRlRgQb48k9vPe1lTX3wzvDs7tLh
XosNLt/Q3Bwzs0YEgv2awOId87tAiB0jepz4Tm2pI3F+eOnEIKvA2cdD3CICKihKdnJRCkySnug3
JYuIJD7LA8Z/cme+IdXQ0mRBsdziSAe6zQnNQBdPsEtU/plkN6w2/3M87G2Ms9M6bmV4Sz6mfP5g
cRLHu7nGgKfjXDhYUl7PmbFrOlOtyMZnBDYrq6kT6nIaw1Pdhvj29a5wrZ+gJJ5IwcGHniWzM2j8
Wy5VeaYqYmpA+V/wLPoo8R1iTdhoHDGz8hiI5cMFQfW/9ivAJi4Wty1/yd/U/1ES7XzJLsdZkbfK
SsUUstGzujtbUgCS0l4uuDx5UKTGKMCbiOyROwuxOu/brF3i7kMgApbbVhW5TLMLQu7OYCWoP8zE
Bizw1wgI3s76JIsTWW10vgZRwtv5ramWwTRJuTP4sya5jI7mUKnyee2JQyfydlNIISWJAC6KoOq/
tHcAPEjLupUrp/E1dRoEKx/2b96NkUajTkM4oS80RJDJHrVK9eoYXU1ewFXsdxrmZuc4vT3TkLvw
dMuoop5sqIxqKeDoGjPeRAyz+mXNcmwzzdf3LQ//X2ObCZ++6ECEo7h08lBfMkKtbZoyer6gudUG
a/nU0SvkhbLmLzMpAo9rO/DCNbDDUuhl+tFz4lW5lFt8COM/wT63LZ/O9rwK6RB0B24kcbUl1rIP
FFubmccPWMtA2LL3C0j/zO0aBTs32wteOYqOpMbEcvbsf7219AO95KN9gh01aS/BFJJXprR+FGND
K/8IVAIYV7249RoBUXLod1NGc/t3cSxLhlXmBZeObc20CwKnpDjqXZCP+82XcIbXd95H6jfBTPh5
wG+i4lV3XAl5VptbXz9oiZ5z3F8kk+5dKQjsJjPAOLNt3I2YWO0sNxZPVkdJil4knLDgyEQSD4hT
3CHevbOmcX/3LwO1o32KZzPoyDowDB1teBrdfdMTo/VUerCPUK/kUP7RVZbsJbxeYv+4Tz/bqOWn
0z6Uu+oz7yrvk0UAJQWqq4Tz5dKTQ1AjeUoSdeN7DyrKy6OogN+yRpaXQaRix011iF0IQnFd3z7H
j6mhnxJM5mTcnjWlb5eZBZ11YZTz3u/bJ8frCAu1GrhoqvyfbDLZpYHo+nkvh2f8jtQ9HRq1iu9/
fVCK2FaDBFlh8Aq9AYrcZCin0uT2GCKvuUATlLjZkeZGTWU+JUgfztR+7D/zXU9fi6fDlfxCskAN
RCU0zVkYUyMvJEtQykbtwXoCO/u7NLx8/bJ4CPwvo20ULfu/ttOsF4r9vksMsKaTXmNA3X35QLDD
UEQ3FEQ6ATnI+drjGY62YMpxes79Aym93XsB4HB8o1qXAco6+u4BmZn4KaH/wN8t+t8MhBW4i39w
b2YwQqeVLjg4PAYHZfFOTrK2RCyVzPQK618k+McS0yZXuGZ5XPCARMk7VhJp+CV8QyBrLy1UuCI3
3LiLsWAcvViQQuxwEq7bfEmRYZ3/reuhNh2/z1II/YLvKpTn+98XVi23BGKuHHk2mKvxOEad9jc+
gB727PWboz29/7qJ2nqIJmTt4gouE6mHzpm/gerioIHqxo6cckWkMfi1vm/stHVY7PmpzGXiD5JD
/sQQ5sL0C0bCbci5io3Q1YwUMy1YdMuAPfYmoTpiFWFTHvL5HItFuPzZAttQwjEn+oojxo/PYV/c
YHnL5BnrN69RAEhficKbA6/0veF+yK1KDxj8y29HtPHxMsQKbFBGCyA+I3LP5/MNcu6qs/swshi0
/9mfxfXZOd1sjEin+o3pej5woKX4tJyo4vI3rAU6ROdf+lkBoX6ZzdB9Rk5D8hxMhsw+jQzYGAZZ
GDy8s6L5nDFuJp0kmTY9brGjJOxiT55HeHJOX4YsNPlsZkEhF4XEhSiKT8yIX7vVXkHluCtJjR8m
stmQOsyPNUKZcHW1sX0+xsNdvIr4cvXVNXcRGgmjrSZRtflgxEy7c/c27+LoVo6SvJE/XmArxbJh
oCt2yP93USVHlZlBSyIsOmyompLMya/PROFzqiOe59eYGTsWZWmXQ5LN74Si7IeFJ8Mq671e043O
emZlOUUc2buasF5NXDy81EMpcAi8CVxkSLNE+45ykTvOWa/pIctQYUJkib0kFxTVGUPSM7e0PIGX
IvElQ8XAUywDBK5OeP5zJ9twY1h5rHly7XfSFixeUc+4xkgnBO4sacOhWgJyFfjlQmEA4YV25Fzz
0fDPkaPmTAE7609m9l9yfHhZ9sUH5x3c/A5hFNXHINgQI5FQzGU8INJAOyr5IlASpYQqYXkYPBsF
VQ7oZBjTGWli3l0ckwOcbAzpsWiuXge4KF/mjZc3lBjSXXf90OtwLxSav6ebXxSBoGaDdu8cS6NQ
eLrWLwaHzPuL8mv4svJIZodsQ+lQulpoYCs3Fh7FxwbMHbnNbN6lmy+hUYnX0aM3aPHDuyDNA3dU
JtCLx98aT3FQhIw+j0kGhXWkPMKbzxxW/5o2uMYEuhsghqVP42fszHzJenNa6IWeyqoMRZ+OJzVi
P2vhkOpXY7FfWujC+UNNE2vYqm/303WO4pH4/AA78XR0GIosjK9NbljTEOhRC+v1MoX0LD2P4oKX
VZQRGLGeRdk89F4gAgvjMESSueaUtZfIEJ6fJTGerakiUZlSsbzmzNVQgfrZ5I9k51PPT2q/bXav
nD/1bSTJajWxUc7rYXRnj7Sd99106VIBHkx3Oxd//roDRocF/QPVP8433SMbkGJdaX0YZQp2ziV3
MJWJNQIvYzaMK2ZgAeHehmrrFXwzdsnVj7jMmAtI/OzjZOn6INc4PcMeVMbfx45muZG9zEzElXtG
DrkI+7b9XUMgSs0roZB99GvsEYRpZbVFn29nBESK7LztT8pkHggpGE/sL9lBwHH57UQwuFOa2Iue
BaurTfF5P+fBblFJg4Z/pUgzVnZRz1+zEuD6Gimm63TVtY5aimsiRWMNdv9CpAfZXBuDYtL7p+1n
MPL1oud71MbadNEyY0UsAm0Gyin+HB8ENNDQsNko40nyilNIGHOLzWp15X/yasfqkXerh+87P1io
WsNxhW6i5gP8LcxnOi6OEZlZBIm/zZ7tAyS3NE+J3tXW8A8/Jr6Ls8V8Li3JwckTUgPd8TOVtKol
rsxgt8+dGUB5vsPTrhpECk+QGft36cQshFPOUXZ2CE2UsjiTbTkbhTdDqIN+jPINRxyixTjUvRv5
ZZhkbEWtv8UY9Yq5HRPenZCaVKaywhhBPLjvV8G2aEfQnjPsUl1WxEeiUJmwQFtQsm0ZZG9XIX+e
NvwOU+g5N1/xg8fOKM/3IEp516P7J6IXZy3OmpBxTOS6KPKr3bFsiOCd5ma2MFfAyFdA5AwNu9Ju
qD7eDgw8wJyy20hJu+0uHWcciV5QhRRmhaJFqpFdV9ALXO/qWnvy6AUTrBLXGuh73zu7Hk+CtMg9
SoqCYbldnxdlWYJFGFbUY1OC+Y6NTGlhtQhutzdy6h4E/VX3yZ/nLzXcY+rvGVNRyjT1jusIfv/M
dg5E5d57dfqJtqbuInSWhAmQqgvaxaOO+UFI9YyA9BbQkSlmlA4tTzoZarYuSflbNzfK40FyP6Y/
DVa5vrWvsziMRM7HsUdYkmhLKuDB5dDCyMyTW/AG8lXNzGmR4wA/Nao12cs45DqnfKVHYP0/ui9n
2BPpU9iuwxpF4riaUBz9KlY1Eps4jhASTzjC0wTOYnZEvemIJDcTGSWpgTynYppgDYv0UGQm9jNT
v0F2cX9+IzsPIv5scaPO8/WqroTj6ZBod7MBj1Ef9+G5mTlUziL9/GaXeVHDJ5AsIVBxzc0VGvpu
bpvn4Q07hW5z+fwhmqefluN7VcNZcSL47hFZ7vrvDjXR7klMURYqJBV6Dye9YNyvpWWL8eVfvYw/
6xEVa0jzam6xv3l/l2DMh385CUmhjRljnAC/Mwv7iGkifM8NtGHYeuJ2r5Ui17oDQSLwxcnJRmZF
bmcJy5FT3SVe1SRx5Lk64erNfgoGlxi3DmtNqqV8fdI+po2Co+imOloI/aQIPqORDXWhF/5a5kX2
jpf0mNh3sqXB37OMc3ZsKx4El5wTJD8jjrVOHmtW0Re7D3xQK+o3+TlkmZQUsizeq+Zpiem00pTB
GRLVSOvlpmLKnw6MCD3/ATyuNZ0LD2HCSEBAE/rb11wshC2jZTgY6CrAScRoMjbNgWw6mJpJv8y6
epxp5JvK9TKq/VsX9Eo6EO5ICKQvDsOrkDyuS2HNMkkRCVI18uS3HJsxKHRkA2OzkUfEsG8UonUS
NTCOtbrCjirQWmMKVWgYpKAfXDWbzjSD0ZRn47/3MqjLgv3oQ5k5eA3TIJGzNqfCn4MFoqp/4H16
mzk+ec979gOQwFZygLqGy8SElq3nVBqdL45XPwV8/GzOnhj2pe14rIi+yjeYJI6Ilkpl7wzfXYMP
GChB8ePvPaY/R7/Qfz9rRs6Ks7hS0p7Z7SuGWFB2ITqbu0vUkdcaNDJZCh/rZKarvPAGiImBZZ3a
M2rTcX7O03lEipwXbyCt7TldGMFrRfqKKSr2Esz8xq2MlWkvTF8B3JAXQC9Jk2OfPqh17w6RwFFh
TfxpD62gmCbNXCbuTZeRz6iFBNpXdDtTaerL7mswzKk3iaH7N6d8xvcrJkTpCnETEoCiF6twhFpg
25+VGcOzG2PqehNiimZ3mgkLOW5uof3qXZEuPHDWBv2ZXUKUzEzgvJ4CBOurmS/myVSalQBuWbCE
Iqw6cB+ewIIQZZ+n4hOTslL2cQ7YEf9DOmOZxSY2z16RotvIaluVklQ6qNBs50OIXkUY4fT8seCt
h9xzG7wBbnnn9arDhZV1+DS5yOTW2luDxr0VLgikQKj/YS7qzp1nyB9GCtQL84lRf3y/69mEM63H
bXQGNbpR/tHEIMhKSvIxIz3sTPddEx0bbiNohpI1ymWGOLp+NrvPtUa3OLXOZnRDA9pYMqQPzE2e
jvRU4qODOp3EipzcqrNWXDhq93wA+AT2cOKKJ4fszHwqBqJtNWoQUmcZoVhWtWJclaulz/m9ef9J
iHsS7hF9gGUkeCYJs81gYy2ytpqzECWyy2cY8KFo9NbiKr5lZbQ3u4OscuzJSTsClCQP1+qu0+Xq
AkD7Iqa9813G0JI92RfgfEqQjrfSvdbgZG+1RRa4EecTmz4crd5p9XfLIeZga9EBwn/m0eNzrutU
eGvaTE5dMmwq2SM+5aLI04ayXRKrJsqCG4tslGdg/OAnDUrjYT7r0Zc41eqT9Ee8CkwrBowX+H4d
U/f1PpKQPVryIMKkGjgmiyys7aIg59D2D3h5qAKNO+DhfH3/xa7X0Ay1O1YKkYea2hZV232Np0DS
wpSLVwKz7BtGW53SSa9Su1n//DxCurdHFnWh2jPlg/U5FBqXO7VvgY+SSDvmCc5VQTYPRvssqCnC
4a7472hHJ6gYDOtpvbRn/m1Nuyd2vsPivK7EUcsmM5G9SJnevsGwSK6K0vSO1e2+6V+AuEM+BL02
nlOswqSaKzGpA8Axf84/9IvSFNrAM5NPTZi+loPRfSPLvzsirQZnVhw4ZIksqf1EXBmAci0lip6G
uznqp0XWDm+V6O3qOmUKmN0ertWRxd/qfXFR2A8D90xXm1Dhvxr9T7O2BL+AIEW4zF054HisDoKY
GkEjIVYGvz4wwgjJVTf65DmhxoQRK1vtSfIByE5miiyc8EDZovm98QIs/DGVCieNJ7mcf6Mebn78
GjsqbWORFuGmjmxoj09j2NpQdQETVUouCsuL6eVwuSpWIijSBk/H32vQm8yFnipPBnF1daTcuwiv
ZXk9qdArrc6uE1PXS2gAE+M5dowP4IOZTbvIRumbZ5ZuNkewdtRWVslmJb3HujVBt3Y55n6wlzkm
MuOwAoQ72RInaIPfPKRvYhfi+W1sfnCpf28CEOWZvhl372WkxPf9dzLOG02+d2PoXnOn8jCWyjU4
J90PmxmxxZCJoJA5W/sPzQYqFAWMWFjI+Bsxl8zZb5GiWdd0/X+7bOaaPv3W68d5pRygqftDWDCl
KEzTbAZmA3zsN0pNXVgjAQJqb5muUZUWu9on/Pv0OqdcDcj1Ky+1ZNKn7KmE/Rc7jqIsz7nVDSPk
zxT7szhGdgSY7f8IfROsruO31S7F24igo44EeOtKT8HV4Sf2fs4eE5Y5XLAhdHN1MDbhkS/rcGab
GNcA/t6sWUw75zSkk7g8ygaivkKko+AWberikbJxz+BQtIppy7A8C6U/IpBfIKM1piYa7wuY9Rep
7F3zz0ViL24Cwb+RvMsGnuLJ3O0eWIOT+o8Ma+A6eqZ6IPGr8i07mXa54XDylA4XSGlG38DyP146
I6LalRtfkiz7BWOVEdEkMlB/t47lbi+ykGEmzZ6ba2eXSVBH9oNaMl+pNoC5HIX3NWSHobmCOkCd
CNm3LaX6WQ1aImnPd6Nsz6hcFCiCdXAeoWzfNvkLY41CjfzU4xn1zHOFBwSwxrLz6Ej7H1feXVtY
KeVAhQD4pzuc6fRs50i6WniudTLoLAMMYWNDMXFzNC46Kjjnu/e19o3pZzEMvrmyYLmSNExbrbo1
QCLHttidzxJDsuYT8ylla0rrLDdRR1J8f3mdQEMqyQRDLdKwNIzvGcZ+daPqV82NHFKgxpHQebTq
g330hrWWS7O3Zf2mUJbYCBnmVuLaytd9MzqNoGqErK56lMG8qrJWnLThHag2AUxFtuEMxm2HHftF
VtDNN92UCGAORhFz0k0cTgJpy88uR5OAc+LgIXnURfWydp+OsWg0FcKhA+3Zih86cWpP+CdaboWn
i/0V5pboHzZknkPrcd/ZevVERWcsrwRXZRwhYP3UPgHmjo8JI/zqY2eZ2PO/zFOdpKI+DIXhv+hx
0kTGJ4aIxJZfDIjVmxUEoCg7eWbymjS76w+wWdJ33TiHQjyNWUx6gU0aN0ZDn2A8ovIAnCwtHg9P
WY6HNz2iUuRdhB/0UbcEg60/kqUjMcjnHAJ2Prf/ELfuyRIrOFuFBofUPN6E8CNTQqYx4V27vH+V
wi0lJP39E6B/pKAwqA5CvjjUCL4FGT9HUhDVgbxmxvQZU5ECgXwpN6oPvIf+/f9d2HmGj3i9BhEG
aATBLNC0UtaxXuFeyb2lr2t6ourf2N669CjsRTK/GKl+NTm4xehmDkiQPnc3y4LevfuV3cntu/rz
GlNVwJleDsdW8hxn1KCr23O20FFJw6rxwaP0lY1X4jRTzHEDUGt4EfJAtcPB0kQC9v9inJa5U7v0
p4PgoyDLa31Fgn4BxdDIxtjim7sJklsDUHEAAqpfx6xEb/RHNwcmr7NKr156ksQdN7LRxDwXDwb+
ZciLXi8x0mNYNatWBJLNagSeR9VySdbMoACmHKDa8LuQglKvguL6tsbi0+VSuQqQcme0e4i+uPYH
09erYmANNh7hk8TcV1/zl+zXEGbfm9aBt7GrmGTXSLjby3WiK6lPdap/MSEnXKyc+/8rJ4XBRnkZ
nRKz3Ne5eKnCzhzI4/ZsTONHr+nyWk0aMEND3PAVuJa1gaoHEa2XGCC95g0FlYgZ8jnpagVceWi7
L84HlC3ws5CUS/O3TASI59uGhpWrnQufj/4cvpyIC4rMvurZIvCARJwxixIW6b08oAT5lBIF/X5N
tRKMdGhOtnatRu3RRrzatVNEBe7+SrJY1IqLANgXcrwXsnxJ+VnFVQ2fRsn0AZKLZU2qvUAGjYGs
fXnHKlsAOASijI09TN6BLk2hlPXREgjGwcwTtns0d2Ewlg1I4IPBEAUa1VND7zkHlEw2/mPPN/W2
omXvc02Ejcij65atN89oJsk8ZC8HW53tNRToLzwPap+om5LxMh4Rkuq8aC3pe5nglBfYiHPXHkKu
bYGq8CTkkGfb2hRKmjDPxIBDZCw3ntgLD0dNapbYWf07+FLblczEg36mJXmvnrfHvYdkL/WfdJLh
9tofS/D4Y07UXOIFbD41rYsJyfqeEb32SjbBAhiK4vBnMthmomnDj1/+yMwtZLfMf82+RTQcpDQy
k5wY0rzi+A9NX0PbDpVBZN9JTu+eIkKuNS6ZM13tmGxEuYdDFh8qCRHuCrQKFjyDUGce8esYTN8E
ZkdkmGP8nTW8jiV2+HCrgf9UwNOvl/AJ26X6FsKG6EOPxhk81u6Fad0EKvhbhe59Z693JWKFkM36
RZMDc+pD3tUFJBe3WfX9SJPNMtx4jktRVoXOLSte8/1LO1X9TvT8rWdKc3VGVju6LoCCgyaCxuKx
jOUUVepctlrlQZFtH7Zh4T2EDeeE6zNQCcyAJuInEawd7PTIK+f2I0/MGkICgw5eYQ07gM+hAR6r
zMyHglzt7rAXHYgZi9niu2ejC3I8C649ZguhqCwU4Xvzt7TQgqwKRwHRHA72/eYu7zPnbUxga0hc
x6toAo0TEJzPWpy3zxS9e2i9/dVRW+Y0ZrkTeSS9xBu8R8vOdp6EZS1OVz7k+wDfEtaLUlXGN7dP
MNwHQtsPaHc6GKC7zQZFVECnt+bky+uJgllJSkpRSCbUppws40wHlFwkcbTZJajCn7yhbGejx9v/
kDrIOWyWHoIIfWKkGRH4esv5ykkJuyxdZcopQZhQX648C7MQR/Z3LZCMitZk3BvMfbu5wqQf82Dt
wGGMrvV0BD10+6GIESbNKvBgaf/AAOzYYVlCQV1PWt47zyXnB7F5hlaxj9wTdBgRPZ3MZLH8Er9J
ii9CljHdC45o2tGFCjKoxOyJi4II7ez4gv/9yOabRIYN1rDZQ9u8wJBdYzhyhkasce+ofm9Qpmdk
3iOm6hjUAgoKMhTFPBJrWGuluQRYDqHDdzhbTcUdVrxFKNtqmPinZ05x3kDa69p3Y91JkXqm9oOP
SUFPxarcoKUx8k+xtVtR+/LvivRe4zNvZbEgNLP1KdW+jZc8q5pWdN6D7IbuaEZ+1nyAe/yVms5F
N7yeP5hLcuu5ZC/OSgquWA0RQNfxqAuWcc3dbDUkmoSeHAQCKtu3dbL0awqPb8cFKp8FsBuD+w7p
RWUED9hoNiXs0j0kI9S3SfATQa1rhqyajg7kXcxtFqx//D5WQXMTnfd4Oyk53lwOSFpHAf0kIn2/
JXsc8w4IJg3BmmUyi3n0R+1gDSyoWoPVHHJppsE/2Ej0Dz8v2pX9Wv5Porgta/bVkTF7/UHTAHYD
heRvbgH7WDSyDP72hQuwd9QPJjI4HVpOAUtfRpmI84Fsq91eeuRsgz9LrQo4Nj8sWGo1idMbZoy0
BwJsI3IY37Z8qXqkAciy4e4/y6avX55yYQgjhwBlRoaoTv2AnXcjDI8IsY2IyLCLCGvoYJEsqGmE
TNAsbqCfBTubmWH23FZ0yRGkwLsGlujZa0dB8E0eQFRaYCTGczxJ2xq16xB62nw5FE7X08+bSFDi
vaj6OJTLbEk6rI/eIg6GOYhy2WOFwZ0VKeBINhRh/5xMKjejLMIi1yc3z7TeU2oNWH7Xq7FbzrA3
enefRaDxRX+YQJVEIScGMXrb+eeOIUY/fQhV/3F7L1DfMyAZ8BZr0vDf1CxXZWEjGJ7iavIR2siD
effq3l+IsDuEiHgnKxRE33U2BFZaPKuB2123vq8lHCvQO8H8vRE0mJb6dN28COLDi88I3AufQuXX
f+5vwBPpAI2F2uvMelNck8sxFXr3a/e4c5YZ4wO3OrthKCkgVdaDMn5r8Jab9MG1KjefYJjOABxF
OfpwLrd7WtxyAutau3XCFVLjFMO3czJGRzxI0E7csE/nVSPH4EOD7vY+K4v0Ap/Fp97pdJhusQWt
l5mazjxtuBVWbjVtkqcjEtHABOLn4Wv8rC+t/Hw7Ha7tuT9IMlN9BmixflTQNofH7y6QY/KSZ7Kg
TqHL6M4IIUVBiQqM/RtH7kcBLGpaFN6/cjD2KvY/SVoN2pGDVbCNNjiLgQ1xpZ7Anvss1b9u4S1k
MIXYxXwKwGHCd5vpDp/Kh5wWqCM7EX84bHxDaEC6UJORVpQ/Vkn8AdMcaiTBFlmUIxXs8S43HLfc
dfWrURdLsLEpIqmG5FK5uYsAFjDGugVR4IFgOd+vYLNsZojFV3G93CNrAODd0Tn+JOrjjRKJr+MU
xUdpLG3PsqvIvvD7Q/rrnJc7I0f6EdnOEsB70k0Vpd0XMw9HuHGACgoOeuxwdwtyQe7iivKArtrX
m5eggSSchansyImIXJxrXKynmIw3X0Vm9qmGEUZ7CE31F0b9ptHHH33yjMv/tv/B3OwnQGLDtVif
LXoo0roBea29dvW3Yl/G5YKkzceYpAztk2I+xqa4c+ULeIHON7dprGHqj3buEiIqd4K14N/LlQr3
lu8YgIjUOrWa9fQEfCqIkrFJE1mi0+kBkP5KcNncAU5nGUgltXL17FNDyDHLG9yfP3YInODLuhvz
F0+fgeIjugmnxa19TuBCKFdAiKn3ZpPBEf0/7jVbuhY4owFJchjjeu3ZxopBpkfu4YLsnyGnWFTk
KEfk7hUdURHz4fhyr2YHQFQs888a/jspnnCua9oHCpdxZZmDH2Ki2JGdCADbvbzC6NOw6ldCTfBn
wxOrGBiVTi+uF3Z5eVTrfzPgiRq1OQN5v86d5Wqhmq7miLNZn/239//qB23Gl2fuJUoMslt6KA0g
wPvacO0rpxdHUJnfAeXJ59w1GEb08VH4NvLocx0e6Ts8TlVEugaAx9BGv375UgEpZ0rvWQ6Vgj63
psNIHaLsZK4SAkBD5M7KTjkIDF43kjqtqY0SJMRPKL4VYqMFciiyezhsqoPLe7CMOpkUOdkHkJ6v
N3c29gf5L26n20uKvdY/PSeYOMw0JA/16hxC6663lZfvZ8ZlAOHBZK2Kili1j43WdJQxgX5uQX2p
y/KAAAdkLZ+k66uHNtugbrr7M07fQdbE6vEsjYH1L6lZlD7bYHpETqGWYhQZcdIDomdI03eInpK8
Y9UC6ZZMnvoc/Q6D48rSQpRF28u/SY2aCC2aPYro19XHrFgwfnn1t/zLSUUScnS+zZmI8lrKXjHh
B8zv2afgQisg1QD12alIa3iGt0EZRIbTJQk5IDYQDMRmmN2uEWSAEdC7j++/mgA4/9Bl2r5mD6/k
SmoX5hHwUkoKfQVpTVobe/vzSkjJBq0DLaO/Q6XZHecNhOhvYnPUHJEWpq75ng7cxx3ZSxSzCkHU
27paRTMJnIALNRrmNi2JurFHb2N9HD64ejH8h5vsDCIqx+n3nJZiqjzTJTIFMhHNVi9+LZ//WDcK
3ZPfi1VJSTE15rezJHRvdGghq3s+jTShklCEfZ3LDqWd48aEDMfaeSccPbnuwg4iYvgQFcZDf9xq
udoptW2fG+w7cun415ywmb/EEVADuAitOy60FZV0O+r/RgQxIc5xniI1cS15Ycw8SDY1upFrjA0g
TCsIPFJOKTm0LLCpDMKbgF25k86mE7JwD8w/9Fukc5yWQZVBhEIfKboWB5SMsRL364y6nkmS49c4
enovDl+H3nnhUGXhUICwbBmVUAvqPXj29eGnCD0WjNBC8b0Obk8pm+2pDoSdqL5z6cd4cbKwxCXM
rc9SMXtn2PQATbwvr4nHknGzmMIgtMrEPKZOmp8O6Q7TESLm6E35Xb05z1GS2oRDTnIIbz9Sno8l
pmrqPRPL3su/inuGqgx/5BxXxXlK4MEGWUBhvB8C/ygl7LiXDU8KlKZxUmGwDNWQyJlOmBNEtjSv
Y+hmcAa5FBqJdpZbAZI54007zD84YhNccuXm1OGh3JwxWViEk5LReGP2vRTJj3r2cAc4Juno1naj
izdc4SvgKFf4WLQXtu00E9KxRL9VlcMtJPYci9zIJPpB/lIUDfm0Gp3mZTrDnBy5SKGevKhbu289
6UWuTC0UsYP9rmtJlPdRR9riWbbyrvOk7OFQ4mnhJSatGuojnVjCv2IX9Vg5H7JbNXq80458qmxo
ykdOGu29cvFIeRxLjcl5GY7jQecvhQ13/Km4n05Az5m/YCf3mzvrVMCihZZeOhrxx6N9pRGJskOa
GjvZK/nPtbXYTG1jd3+CnO1r0dYbOpxgcI6fIotzPwlw7LNtenTSZPPSX08E89EvFsb4BVMgq7Mw
VA3xcZP+7+pMB+OOrtoljVIh4/2Ne7Ty75Q6G+SZnj6mdyzC1WB+lOLtq48pGzzIO2IStANQB4tN
ZgPXGSnsPBSvNTxDlGFSaU0rWXzPbY7ZbrFzC6lZCdIEj+4lAKqBgOX4i2Na24nxmWyoFteI1Sda
KUqSBfHTwGGGJkSYsTSEyjClolOy33Yyv+xPdqX+Yv6xJwLTZSPQUXtIqwGdxLuus7gsTfEAHvy9
UUcnzjL12b26ShWM36ppuoQOyzs///etOBr/ArqnkwwVd+uMJDro6/fX/m6QRWQjMHiID0lJqFPe
/gdSKkiKS1tsDE5GORxm8J4r5+vx/BXVx3d4wvVpNyzZc+4G1C3abBdSdLD17PZTsr8W18rOujJ7
GaUl39lHd2B5pOMkRYuKGme9TEUz/NQ8NM6mCeTR7f1cThGIs8GIKfg2T+NQ8SNhHQhIWQpEidrp
VVg/O7pUDmIGx5sQ1wst9JxZRUxlV8rITjzt8kO4Hxhe13t0zppM7xE3KXe8jB3fSqZMJfb+i8sr
llmeEgPY/7z2E7SmsdZzJI4HEbLEwcC+kbvOeUZBvsrpVlNYOatiK5m2WbA28FUNoY6Qfc2zmm+d
4gySx0DTE5nEbG298THMxPGR+nSB50Y50Zdhfs3jHNG9NIYdftobYAtUgaLts1ZOGMItID2sPjZi
g1N/TbWF1UzVvs0mQ5QtCpz5qjCbmrIbYBrkBAH8+AeCRLYunaM/s0Ddu+wwoCI5SNQvfTWI16ya
uoZaBiuZxCfMDcUKPlPkV+MzYe4AB7NjrYXzO4KIcrXGbbZxmsMKA2eGM2AhDPxoaohqZE6hnZ6t
RJ1Hhm03hxHTGfgpFdiNNBS7GSKj5N6lj3N3Tof7Y93bkS6+/+uDHEx5comanWDjoQw6MjtLDDu8
tSJtdvs799P305TRbUnDUqBcYD4cTlQMSyAtxDm11AoyWCBtKPHoGGn3eDNiJB+LfDvNaSa6z/iM
N485tf7gwzYvM/XsPx+imnLc6XA9DbeRTCSWYx517IZiaNO+T2JaUXE2+sSVvTSwrxPRfF9QwZK2
e4BFWNWb7I7kZcQ4U6akLp0PzMyfZVEfABLVg7k+Svla2gkReaD9TISbKnh6rzmkhIdm9aBs1jJP
jrJTIkW/AmVT6Zsr2e2sKaG6ftdlMtsWcRKSXyvhEEEJ4S5QszFMRd69+wDS86svO358J7ynFPoj
TR0rKKy4MvVCW9DoVZ9YCL9QOUSITdG60lrQE8Sn2+SXTG4jA04zfX4uAQJwYU4FthYIlZp+u1z/
Is3sQQJmlgV1MOkPFB7NkmvvNP8dCAcdk+d9vQPycjZFbsOjGLGZiiQuvRvFlrX1re5d9MmjyAhf
GueAcuz9DbPHvyvxLRwNLNQs7uBszFHgBvLg89VZuWf2RwxHB/8q1R4knEDD8uU4CrFWN3JD7nuV
nmsnmPeHp3xrMvJY0Faw1sh2eOkJpGUkb/P7dkvx9hCJCU046aPtX9wHC6KDvUJkfetBMSzDbAq9
zR0t1JqCwtZqn5sNNkv2iyDXy/wazHIRSNLCtBpZ2P/JHNzVxKmDAFg4jPs+ffLpPxHz4sbO3Kon
pZJy8uOcu8H+SxPd9mCLHaFZJnppkrF2YXWtC+vIf39IarxRyzQImptk2OEGYRkzSOcKD44Ii8A+
L7oGlqT5YhiO2now7yT3TT76JtoVxmhp47kLdI1n5GJ9KAfyMMdIJTO2XOBjSUUXzSz6nO0XO/J4
ahJniLlw4H25dpGlEquVO6Zd+0slnqU1KFUrwyzwnzhHzEp0iolZ9i4/81kKVUZyinNpwtE0h5dc
pdQLSOQWEb+YjC3JymrNAmMesknFpwGGdzpQGdKGFmfDVJwldIU9k57SCfTkfqNqol2r9HsFcVR2
WBV98+VmW65Zo/dIBWNvpZCr+sEhowZpSRyprQ6A0nMFuPw2xbx93Q23uYpAJf6GnrueA2I6Ybtl
xmdsXynPuaj9o7i92c+OjExuqWXUASogqs9VubczLR2qHAvmpEFicAqN/aUbNngtuz5RERlxbOj/
zHef0vj7DhFCWBYy5SEpp29yj/8RSstnUv3T2d5Se52McpNID54plaZ9noekRdFiyXbR18jYMs76
qI+JTNud3rGMQSxgpFEDwMTiJ2C1d99lUs6OPqB3zC1ADpLrpAxx2Y8puIQUQD56NSP8PaVFxkNp
Sc9yt4pwTdhBx31+ZwDl6BX49MDpaPBHrLbg83oUBxgbP4gdi7VJHXTfgfd5DCkMON6uATkYJit1
rhmwKt90j7EZJ5l2OAOeKXmbhgtnMaLhmohN91WpEXtKTYI3nFvRxC62pHbJc51aIofwVIxivke1
FT82hIf4o6CLuEVlmndfoa0dvCGaNKaATTL+/4NCaBThA4z6rHFf7j9HAGHLaydlUZYAl0UzazAH
BEjp9oWGULpdREV9Itxwj8CunET3zN7CQeUgViTE2+6iRntSSp6donrHX5fXv+KRdQhSYYVrrdnq
c1FPTHsq4tkPiXNqL8SKCpWJ+qZMKsmZZf1kUuD2nU0HtOVC0JQ6p9loATJctc3Wu+OafhgBUwsM
GXoVeKQMjyUi1b+0IoJG41MuMlG7kMJWzpCPpgn6YJnz5j4wvySdCV6l00jK8Mynj92lzxLsPnT6
P+x4B20LRsKAXqW10Dl3q2NslQpyKPpxjCqzxZlwOpLuRCY1xwfIIqSHIqCJ0hiRHaxMWfDAg87Q
r43sL+u000Jz2itJw1UnB4Xxx6xT8WihGDrMhycUS/kd5dADDWbng8/hqXjcLNn3K8+tof4qe+zv
QfTgNE3oGOZFNwxHNnEM5j6xCIIJYmvMnVVQ2eTjOUeHc2ic2OdzSp7FreL9tRj/QDW6Ol020Mlv
hiuETzY08nVmX7be0tTTsn4n81Z6ul3xMUpJCg+xeoaN1ZptVcjxSTiReN6pYOvOCWz+BSOTsaDr
Cse1R7TrzTs6kbH8cc9W5tjdczwJpSiBC84zlCv3cUbYrkOEMxRwFWgPhsCSn6Dlv1r6hokKmFS9
tN0QU6EdtMwVlLtVHZboIxmdoqNFJzOBtDwMiWa8K9qhMoMHURr55GVa/kBcjvB2C6TzzIm9nYzG
K9OiiKAEJNHFUlBQDb5ub3BZYdGi6fArLHkxnOA1zLdvF/Q/Sadw50aWf3TcpmDdJzE6805NnG1Z
wuGpl1gQsZ684chXfFKbrF8lIgSyteLuNYvwLP3WfG6IZAJYJOlw9I7bkgzwv7py+J0xszmO8UPb
4hU+cIQsBEu5RwVoADzxbSK7oMeD9qaXis8Jqo/fmuId+PLr6GUK3ouHK9krvEYx0TEJiEmSDp41
WcblA1x8gS1XrpmnNG8FNw0d8o1VS0xzDD75fYyv3WERQgWfLojPcfXafeLIS1yqIiR+/o09wbbL
GHLK8vGvWPl8jjMS9W3JHFcasQ/YSz9cHtN+3XEINkNooQvlGIGTm4citcS7NUSBy0LokHWUcCDQ
DbmxrBeYVsF85rOF3tkg/0IZ7muwOc/LvYmV9ZS9AI9NBOz5JbSKyX8aRhoikA9OR4H7MKpHNLDZ
yl5pDxZ7ifxGjbS6yidicIaCyinnsbxaDYUP0zMDqHcpyanR4FkZIfQ1QJtBEWgd6bCsc5NKx/Z+
Swr6HINDKv84gKwNRnSM2O8bQCJVJ3zudGBux0ssrJF3a7ufF6k4zGOlmpXUUy0/8gZdsuF2lC24
ET+omCdtfIDJtIZE2EPoUIbMeNVTbDk+p6g2Am5xFIQLDZCTwATII9bZKcwAno5la8w1wMa8Gna1
chlrM074Xgd0IuI9gqnxMoPhoTZLJPxTZ+lLmqViod7e16524+z/ok1tNAE6Aaw+EKaO0lvGoowf
rwVVzNuA1ktCx3pWXOVaYFaOUyqF4rdEhSumsBvOdnSS+TUimfUKMW4c4TJ9ORTIaefaRQGK+82j
9VZgFFzFTn0hQKG3YtfwX1r7EAqulfZQNWT2qsShDor9Dv1f5QJsH1t8cUId1pd5cLHVtV32AGye
EKV3S5nFUzCgz/teewa640AIq0dR3YO9aBBNirZdmoQqMiBpo1yT19tn5Smaj3hRO7aqyVeiIQ7A
wrtTGX7az/e8lbLNa8XqeauiKMgo4bZQlkwGaV1R0ZX9X6GoqtpI0c88RzZFudiO3wytisdcpIUW
lPLAunWfkDMZgP8mT1l09EFlwB6V+QvY2DmZG4EITQ6og4bDG5uYpt8g9Mq21StnV8QpMq5PL0Yp
sB8IYcudxN0MzZ4EDmi7aLEeCF+8VWsW4uqytE9awxysePCURZnlACwWRNsA/e6QkrvH0Zx/03Cr
EkKIEISzecBOmNWXo4HayyItbYoJgiPMnQrBhQr64ljZL6nmYPtOYThcP+rJdQSEFGy58Mn6SQRT
+vAsCDIqZUieq+BWIxhFbCcE4eeXsOXO8J9HrEOkr+sbous5EJlo+vra0qV4C7O0Q88nR0KDCcUV
CWEJ6d4qIwUNKcujJJZOpqAYFn4MqF+aM5cJQgd0+by/18qnYG5nLZ5/M396SGbAqlg7p3pqjtK6
Jy1AWpCMKTyD1dS31R1wxndh3uZVx1PdnIc+sDyGNEVJYYcZ3WmjImzS1FMH0lB03dLfofw4rXDj
yzPTk/tpE3DLpUag/7zackrBiFGPe9Ltu07Xs+GJy/kOQ9nGU80z4qO8FHeWIBXhjCHZgXWC+LBd
ndt4DATwBUbMUFda2q/HYEo3t7z6OOabrDIDksWFKoFU3npBO5hxBHyT238UYved/vUicspjy0L4
RsfEPT8RdNTmDb4nsBv5/Ck1ramKVXM2l82HU/SFJKGFb4aN94559PysUELZBiknTz1OcZqKu8pF
bo1IuC2ogWKoqNn1Bw7xSSRBjyBxpHhtV74XbI7AyqL3N/ojok3GzxFS1vrM2aNGjgmXvZq+I8pk
rEz07IO55bksi1kTuNizeG/O7OcVbFCfqarwhqQWZXox/Ms6ht6pq9ip2d04xOBwMs8S2baimezk
KprOmobNzP1GxMhOdF/gTrKkDagmfLxbLmjNds+sMAcVOO7mKX8PdpvQNqbZPZWSgUwb1ooAYxvj
rWwFJJVcgXRjpvm6++aWhA6sibSiP8vqOKPaEuKuwp9ntZqiTO1TZ4b+MDFUxv5Lt/c8EGoxVkbe
rPoZavZjuhaQaiUYmGfeUGcN4i8dGly+SoX/MaC37eTVRdbbpKcIEL2IaEHR+UGDHPk+JZn0hTRl
H+K65y0QYXx9ZZ//KeQFeCYKUC3gkctOL8PL/yx4oAP1dctWRGGokGfmr71kwiqM1Hgq797XxMDX
2nEIlx02GkhTPv9E3sFVb6LL7ZqU3wMoygm/fS0PidyQfTP7luJM3sYUny+KwqTtFUFH0raBpAU6
er8+qD6n/+c7hJ/NuxYdcF+hlW+yW6Wq2bdkb2vBAjhl/rrtWbFkrXgn9sE9jcEXMfHR7rZjCysE
Sd7LIwUM0j/FrhfQag1mEvu3PGqDfzgY58bkqZXYrxuS1jzPkyf+8oWAzY+s4lGN/0beMIGDQZLQ
PjeVvOHHEoqVc5sJsD9bAvikXw6P8Xq5pOy438rwweJ3FNNhNDR8aDQ7+Y2Dxww7RFDX8R3vuCc2
wmw51f4bN7UTKwgqqGTpqTezSLM65s13w+jQD36Id/NwCMS3Lgn0uwuk9reF1TSwY56Ml+ga+y8+
9AqvMI+jzEOXfzPTppy1YZVBAmmyA9aIYVCuWX+FKpGbJvzMWRgmfxiwxY4QfcjGx9UnrdbI1uRy
hf6dq7AeFNm/+m5/3Foy/JflY31Xw3h7YPk0QB2qq//37x4xictqg4XuIjE/zGn6x2O+lS00f9N1
OJA9ygIhvkH8W2slUDVJz1yN8JzTs0uXmjHq+k3xBB8dRN8/yUELLqDkgu5/aToBzUeAVoUcOcS3
AeQYWCGEuIjFBCQZLfXsDl07mA8YIsWy9K0+9IYU6QRJCm/fCFISdDYuduSDYtZ/ganr+zFS0D/P
0yjebjUoXfuI4qIaXakDoMbQQ57FzrIjuAej75O/HTpIqbfaZNbEcbuy4CJlfl4Odj0xZAffRik9
nsAMHv0SBcmIYAuvKWzWLL1vrvKEkaPzqTN2Zdn5wrvb4w4Bsd5SfC0PuBtxaw8wE6tbSPc4nGat
Srunnt24CpXh7uiQk5qQH124L0FkFPwa6AL3dRhkytHaPvMvUo47kJ0TOMkeUxYkdG9R0U7kcxqU
2xlEHQvEZ/RLKa+h/9RAaAW+a6XXAnbnBs69aYXjfej4YRm+MiTv6dhjUp1jqxyD3ydGbCx/Y5jc
9Uv7nZaqvdBj8rGp+ntn4mus4R5HhyHfu2yRTB5u7uq29dX1j0kd+PI7+DAarGwoq+Bt80cxynp4
H9HQ7OgGYb+YzBOXqI7wRcSZfaNLxcBwF8QMfEiF9ht4KN3fq6fR2P+6kdaxOoEYmJOS49SkPc+Q
M19lV0vEPa4Ko7yGCvXLiWJnb+rCEpIXj8HN1TmTkQ9mDfWDbxP2G9tU7qzRW33Ot4smpHbu+5Hk
AaH0sNYrwxuRu1BpLe5KVGZG6gHREFBhZq7r6jlmb0gqcGns4LXmP9I2IZz8dbUhV7OInSB7Y8Mh
x9e5BM64sQN09WNa8braaDKLB3cyO2yQK5Nwz9ooolttbenrr6ftORmu44hou8z9lsWsFgKwBHwO
zujKpUgyS8K+J7Fmhzn9O943OPxUbWtmxC/SQwHmKIbZVAtdMVsQ2sI4YU9gjk20eyUH06CXJrOn
11cebRpA5+E8dabbFLWH5UkvUcNf6J5DY3ghT3j9j2mtKvIuESJxpnIFep7P324aFodwanzR/Nzm
Q3pcr0DvIrI4/CvwHkNgpSq5UH5gXqv2+TJia4IUpQuklb4lj3AH9nwTJa0U0GHh2z+XHTO87xSx
e9od4Q88ORnfidHg5VAo5DufbT4Miy2UBb/CGVuPWukGAfDaxeyJhZYdfJSoRRIDfZF4OWzG9v7n
IZGiTl6RYVHPxrn1jZgjcco7FX+Xb3IFzW/x3tBMSsZruaxHPngv+YrcYowXG7j+m0X50pPCG8cK
VFoYU98llXNj4uKBQ7ze/BeLF+xBr5x51vgOtCoqopDXmeF1kGaF3oilt/J0Dl1SVYdhKl7MDiCf
i9iIG23447RKRnTUcLF0BSs7zIVe4w6JAgA6xG9QA8207nY4pGiw56ASlyDr8SwMhP32JVtv/PYZ
3idGWPpqKkzwUqcq3fcQdpHhI8hvmKA5X79zJX+VV7+ZjbTI53hU/2p0HNjRtK7y4BulWtJ6wm5M
jC+BfjdXyDcVPKSAz7heU5xijB6qErAhcmqxBPBcWFOcfWOK8wT+Upi9btNL0zdxTdLtbTkvqdP7
KiHf2GlTumsVu+mip030Txh5kIzyG/zn0Y0a05ZIaBKhQuOL5Ioy9ERl5JjpoKOyzyN/9YDjPcB+
+fk2+WSBJ8rho39dKfyJwy9aVgTe6GR1I75WmBLpaggR3BOwXeik+BacabmwCBUpIiBBjO4J8aSD
7HGc2ENctbLEVEshr+6U+WGmj3wLsu8Oe+y3bM428lT0k0XeaYwCbJ22ty42jH4hg4VsiwjR/+8F
h7njrJAxbCqiMzRqp5og0ycD9NVhFQukfAWj3GTWXrfBbkKB04EkbuA3Prg8FSTt7qO+IcP2t7mx
7n9TOsYiADLX0GOcgrmO16l9j+jaxdBMeVr4KiPC1Fyw2kj0HftXhZLnA6250DY7ZHy6VUHmZWXp
uVf7My84OCe71DY5CrAV6ziX/ZG0hnQ2yYbyD+vZQXB0L6eNCAFSN7GsuAjN3G10OjOIj13oDiRm
aQ+NkH3eX3641KuwFUTFeYnfqa3CkNpICltbYjKs/7ogY4Uy81SpWYG3zS9tTF9uTZdWCPcxvGMr
Ol58sCY/tt6dek11PMDs8HrRl4RK86rsTLG81vYcAKDcsBBindQ4govsfRxbH2LFuvcC/peF7IPJ
3iKEo1Wi/Y5cM6nqgZ3QG38vTJAPwYHMn3EQXTqz+Dxyj985hPtEqCCSPesQrcPlQQbJyP1aO2lj
5OkkFqYuUdVhCIORZhRDz6b2NKZwfDg3xVIcmKwTFJ/evZSS8L3ynwM/dR3954InzldCG7Gimppa
+pRfqJn4oQNyggD5wNnUhuWp2JtMqsIDSCiotTDP/s+l+L8I+32ctQQGsvvqGk6OnD1B1bGTxxQK
lWz7QLYDNWrLtvFObPyov626/FFSFXGzBX4lkbPuIeFP/rR4tq1fkdDJb70XxMBIqCwZ7B9zTULR
k46kwwH0LymhaUYOYv4lZfrHakf4DGp1eEOdWFUhTu1ztwj19tSOpu/YrMQj0BOdc/QSrxzq0xnE
81dXz6IAJk24MiNs43HlAFfMkR5IN8EbvEArpBuiMdNEiCCusnfcWKPQzhKuy+ucLtJNbiUTouUM
HqSXCaMvZKKjl5IqwLzhRvCnLZOSIJ2sW9YD0bXdNhG9qaGabUOqej6itPbrg4G0dbDXcfshWfIl
72tSELBuc5YjyQ6rZm46LxNxXjWqSghtO4ZK+XVYS2OgBFJxGoXUDd8NAhoLUZIBC8pGc84EpG+R
dH74CAiEfydxpd1O/v5a6l8veheR479GZg7FmHTPw/xtes6gdtJxUHu3hKud47ebuCbj2xr41+SH
L9Z7L6AKkjAOXYIoF4yfhWatzNlm1p9YJPI8S6O5Xu6uELhNyVkrK5Yv5ao3/V4bH9xo4BKOTgik
zpRKMwU3Afuk9agOL4UbA5hPWj29OLW6dcot3A+UZX9OLulF8Xx52fb649dLnykHUvkohkqkq0im
Uo3+BXXJsIoy4e2DpE5JraJEQdMyB9K85d9NoQzn3wZrm4cogi8k0dl5v4njp0+a7rqkgV64rxAa
cN8sHYgu/CbFXNRGOWk5sw0tFwOt+SVlV5r+q00LsICfRKT6XF1Xd7HzER3gvUC5dsnMkdGb69IT
I1cb6vXBmq6RfHB1XkYs3cgsRl9YZcGeOil7n9WBjccX6g/2COmIYWkIplfihnQv7sLSnkgvXvho
P/NKfiBc2R60AW07JMCuQuSD3UsC087IMjeePL2sZ8VJKSD84lWxYPKOadMiAdB10/hriJAH+ld1
FJAOEhGVlUnUcLk4XoEjP7usmEa111BNstbw3zGkQtjUVY1HTQKICrpZzjsBrwuRKrDcn4NM71iV
KvIbzyBP/1WW5TKYh0WOJyEoVkW/D14rpjQTpot1PSByVYJUoNdg9c8bhmnfaTdTRPUs/tBZa1tU
xi/qfwOf0JFv7iHEbcqeTeXFYqaxbL9bbOnUR0Q+5soiB+A+sDyZVXTIheAjJ2I13JMFUL3jyImT
tN0ogYqeEkq6miMkRMrAXr0KsRvQk046xPvOTrrdrXWtuTIW7lMTr4tRs0OF8ijvCTx8PXzFKT5H
JX7ujHGd56E20YmSSpuZhqzFHb2qYWICrYR3vueK1DRWAyJOsRwqrM5P4mGm2twS8jB5Iy5kzn1J
UlzvQVn0ln2a4C6pclsvEwLWCAsOZvbfJwGvpOgH/FRoh1QqflqZoJKw8352i/uSPfiTs7/9QsX/
J1B8SsjJb7ds23rEmR36zqhe+SyY+0+i+i6OPe6RCn6MbBrqAJFbD6Aruzk4hqfmxZJznO8jQIKn
3sLhXZUwhcS3hdB2CW3JPFsEhZ1dArkS+0oPldMSq4wtKZf6VrObeXci59cJg1diiT2IeIakhxAg
uGOaL1qIlYaQqT31M+Pp0pnU/V87dQEPnW5KY10MV3k5ivKhfr/AW3BK+EjgFw7lB9UnhHrk+s2X
zdSapfKNbw23yNCVqj+edA1JmHHZSH1Dl9Pt9aFLExNMCcuggbouu0hop5CZ+O2wSmgf4Tv+AZyr
okBnDZrVNEZLUfDC/Jz3WvepBIJlcNQs4RnsZUfFQqEL9wfipWIFTVCpWYJXyuUZfbkmu2gjJ+Ul
vPCxL9+HndhYMMRPqM7tUwTh+err1gHCerswmLu1wwL5dAeYTKF8feC7cODZCF6pTeO+HeTbe/JR
up2wvnmXdjG2oVNzWnOmVZJkG1xfqMdsQUN14Mhywa8QY5994XJm8oKfMQzO7SBOGSUS089olliw
ZmWu9kVSKhUSTF35yrqtBVWOLeC4Q95p7qAYeuMIBl+6bmdxMTHanEHln5bFYP+JO2sDXoDYp0+l
PmbMmiNUgefNEmyRtXqcabmKPP4O2VCwlMlmcKEnze+8z6eK1/upOKGGxkJSBe+Fc4JEmet1nt0X
hKSDlQOXu0dACfcc0h0Uc85Oesw1I0wAu6svbJ/SpcT2mNHcurLvJagvVq7yFkWecg4eSakOYieM
NHKYegv5NZcQrLU6e/AVMy+9TTYOCs01p16B5tXe7Sj5/m4oDW0OTNP2mCqUCi9EDphV6TB6tv4K
1l4EKFXYxWuuTl1feLgFzgS8xH5cMAOK0DSdyC4a6SItXFJNJFs5Ofebt7FZtiZtcBzeNnshBZBj
ytXzyetNGgKOLknhkXISGHIMDl4a+tKWzLygnuSgUs8KujEc3cxvB8JUK/6eNV9rcrXBnT8EnGNh
+UzfAjtcJZs/26DaGrV2myaSdpCBf8s8oXxxrw59WdsePKO/oYgnB4AWYdUaDxpnzMfFI1WDyNAw
zGxddAklqVNlB3tQBkKuIRx+WGgsjdUMtDCQ0AInHucGkEcFox6mHgHPn/4XW+DlgkO7Ty8PN//d
1fs4hb4rWquiNIOGMS7t101kDgnITyJOt5cj8qnvdV1CW1Y7EqTqVc/ChG44QaVRICoKZ6uHQ+O9
GfxvEES9+9nQo8iVDocZeKleTuij6xvgbmWC9ZOMwVsQ32IIfjKJ+SrPP6bauGTNDcf8j9GDBRab
k9YY3kTrtVTSrjA0+6NAQpL58fvZjgX2d+tqRH4hkc+A6sBvd/QFc4h66n0MtzvxFsIUyl8RulV3
yA5TK4cShvThItd7OzpLQrPfbUfwlWEHzQ+PBr8Pf2pYPdzmSj/HBvfRgjt1WZQlxu3mMtdOy6fz
cehkxkQPj928l5iyJtrOdcEJ+lEwMRnXkEmXQgggXWvbOSzNQgeASLYlnUXryJXtyw3X/0Syn8Mv
jlxS3HTKgEFAsIyiNgScVsTUlnCWRBIOny0Yd134mtGVZnvnLD3BbPB1lcaHFfhwajWBixpahhhi
qMsl7R+wBcE1GGwV8owxQO0AJVL+l9nFXpHSZMlt+LR2xMIfbq6gLNG6Jg3ewJ6+hvupxraKliFu
hVRUnOISUKrtxwNiLfsU+7dLVshIW8/yup8c+pvqQ2Mz8LNmI+qfMlRuJLTuDROSUZIwccfuQETI
wLz8T5dxHZdQlAimTnWXmzH2rPQ9Jb5/efjEL/WasXiLmKAJaBNyjPmp0lJi5S0ryRAFI1OuARuu
I2eplKYMQakGESCEoTAQ9WcTQzV5aecf0AOyhrpuA7WSe+qMgwmSG+/WJLOzFjMPoGHD4oeB2yL+
XhnRsT3FZ+NWFiwiP81sTGRIcurbmcd5OvIZkeue/hIYEDH7aUiNRvlv3G9mFry99dhYTix2Jlno
mDFnI87/5H9uMJZtZc5V1BX4HxKJhHX7sVIv2vPPXHLJrXNVkLZ1Lqmuu1J2rRP0QvW8IqxNHVOo
mKW9ltCe/RWTv0WmegGeChAIe8/TNFGfDQni2jDdGkNdsg5KIjM/ywOrUekEfAtUf7l6XQ1tjmW2
TkNFfFiAVrn+tmEMBa482vBA/I2AxiXawkQo8qYjZo/Z/v6BkbGsDhcvlgzo/TU3AFq5Bt6ZjqrB
mmI/5GGWs7Jfboc2KKYCcmKahHntgFejvFJZin9x+uzjJANz+3Yu7o8PpQUgQNBZSI/n7KuCaMA3
vmoLMMZoCJ0muxXuDnS/q3QFCoOs0eXNVDAAcMVsyke5JRKsqBhn3pt16TB3N2X/cgobhHU0t2tf
fNIV8EIhjZ/2yEOr1f42ITkgomDqELGKgqH3rYR+oDwOtGawXkFoGUwmoArZx1VzQWrTItt5n6Lk
1IxGeDNcEumlcjWG2MfHuQQHHgtdxwbszigfX0/tqCLclzPDPf1tzW6V+Z5zZipLwBheOuUAi7vb
NaZ4TwBOz3T93phB2utt4Ov05Ffh1eLaz0Evko3aHDwB0eVtcPwv4ze2myC27AUaUVCLT7S7L3eD
qKbiQCAw22JV4fl1VsIbHf26fkLJIGKc4y2Ol7j+T4xR2AgWX3fUVcWKOQ7CfaElGELZmqZbT8CZ
gmy7h7XCwD50ayfpsKwjmu2+PMnPyjhtCG23TJ5PUSyM4cMSLgYAtX/aXGrdsXytKpE8STboAmFy
f0npgNE9/rUAGbhK7vd2c/H0YJxtWMX1cOs/tTU0eS6Sm8aKD13EtLT1m7Jl5G8vnteitlLWL7Z0
KlJFQFCkr6yUXQntD99vEd6gFaFLQWv5ydMzaBKf98kwo0d74jj4FJ6YiOtvzn4z22jRWeSWRjLR
ngmsFnoE4j7JuUiyFIA6XDhVtzo9j+Q+b+IvApqE09eAw2Pi6VErW1gD3gUglEvhVMzeqq9baqSJ
1UPqdYzMP/u4YEmnthY10oDH1YhzzIaupMAoQlz2REJ7u2Pk8iUExgj24h3wZnD/HBh/KFlJC1IF
rmPSXwcFjk2uqH2593OHG+Bbtwqnd6KVgsxIMemjjnOjnEmQjUhYlALM4CEYB+BLQGdzaufyhC/H
OR+7XhREmStIRHfYntj4b2i75NQpeK0h9q8rt26txoTRTCGHmcDLorw1J27QHfrIuG+SrTK++5V5
p6OCZdfbqZNTJvWvUixOHNKt2BPVgcxebNpVwa0A+xHqxLStuS98miH1awHvS5ekh8FMdwLuJnQ3
fFsDWtTKAQfITp9E4Cq2lSOr5abT+Y0YV7h2QvFi5JDFfuY3o552ZuFovlG4AH5KAZFQOUO6R6rv
waIhN3b+cP/Kpon0fndqDupmhrMkRFEBYdAckCNGJm8ZJlXxgqtZsjpRjAHt2u+JscXR560ylRLG
08GvrJ3t1mho9DC1k5hYXq8L7Bd0Bt3EgkMyR8eqSyR8VbhztsbTdIus5rBH5US/ytlwjcJUTorC
TpzB8s2zUSYe8Dy/GZ8y7jOBoTcChI4Zs6uNC+Nx/9Ij+pJfd8eXYvRrkPA9HayAyzwHNlbc6qaV
Hn1YSMb3pFQj+NUly+6XpkHb1ScaabNVGKs+fKugQ2YbUreHolWA7ofOtgGofOHMABH1MTBdDhzp
BsFceWFhWAkH7qkbsNqKOKcQz49rEBPA4pMAVEK9t3s+2CxhFXKH1F8NgLno6PyxlVjfF+7wQINM
a0Bh7BYckrJcH946gRQDXLu1X37LSVpqNs04yvUw18dAS8dpL1vK27pP0MwdFX7KCCOVvaAAQhDa
/mxGXRklnC5lfR3GGLvOxOE6k+3m2Fmz9GDShDJjVicYdJyb2WM7kBgJc6jHDocQIz0HQS/KGM9+
dPYlr/VDyNe/olCoaHLpoJivYfYuYAgqJTCUDcE7Llu0+JNxPN2Pf63/XGg8q8klQ7iU17KiI0Jt
1T5bTSvBhExfjPDVDZKWEyyTQ8J7v16uOhB3U9yLkG2xpAbiRLvPO4WOxXZngg6B+EeVkv5RzBNu
cdwYsRVvF78saafbcp6g89w7i+7+EFnZbkclVuHL6Unu5/ZyRmYahkX4YhBYsNl2mOcAFr2oq8mN
+ymUklfQkLr/yugw+M7pVVSciZFPutynuUmOtcPlegto1sJfZGX2fYvVJ7q7pYY2ya06g12FNuw8
fDpQU2pWnrjg9Myg/OzWKAaR4mxdxSfXrl/fGw1MCU5a6oVlZY9Yl5wMPfLN314pQxhDAWJ6VZ73
9EMBSRN0qbm8ojjwiXQmxjE3Z6pgqBA+VMRoQ6183ma/2OYpcujtTHLDDCoqfNsBAQHrl5RqZhUy
wjMVGk4ci72ZEmvZx2IeaKkBxGpa1OjFlqjuWFMt0X6R18E84ACcI73Rd0SOUuQIhPZyz+feGQte
OA9y6i0ENSRFPTNk0hxW7rjoThYraapv3xMjueqUfAOONll5XZhMFRKJVpgSa91aqxK+Z7DMUJnA
l13l2QDpz0V10gkx56swLsQDNJ9pXJF3efMcdPkaz8DviCyR7oeFhwTGSkjF6IGskZWQGtseurAY
CIl07Q7+AgLA4I0wVnN2m9gDd7v71F6o6MehktdDKX7/rMA4VY8gAMheX+iZSHGdkKJnjw1++59J
WYzUhftNxlrihJpoDs+K/IKUhtL4zf7DF28ssKNM8ABiGClR1ANDUUKraHfeOqF0llng5F/i9N9o
+pnzgoUqFGnQ5ppJaAZjy1WnSx3L2bjLbCuWV9v8a+p0+q8s52tgVrPC42CI9fcXJZs83vUjN8VY
iA09NaiinG05oZqtoBKm6smOSvAL7mdzLfepOt6Pod1t5DVBryOiY1VSgqIzDTe7aiGFIG9cDjOw
PmcssUEco4JjzqDmn3RRuAhsWYTdT/7gETYW0R+66KUXR266t0QRB3u0U0s7ifjyqVQdxNa76JgM
AsDnjANb/A/maNZwNnhjYyJsmEOl5Wlv57Z5/RkkMvdfY/h+n/WllvBCW1bMkjx3PMVtr/AtonV1
EYRr+t3cXLmfg44axX+SFybSa7dOC1yCGG2CyqE+3f1ovDblw6Jy0R2T9cpPybfoDD1W5vyoptA4
kNoC8oLQYYXMd+uNkycxDaKJ4XmWz5kmJYZ62sOJWpWCIKU9nvZJAhkEQtOc9xtiEXpPmVwhGS3B
64czAlFRKHKyUbkQlJr0z/PIAj1I2bFQb56Vj404Xq1VEMnF08aFDuezaAxSmQEFL2AyEz2IVNq+
/yv9jtboq6NfN+3B8pK32vHRLbr8WsKanrKSZaUC7pKBofKS6UA/MxsJAijrrbYn6KUSi2G7iD6x
M0nyORDKfOWxXzWNBEjP42xzEXyMWCnCUB3oVdd4zJ+vsMvd3usMIcwW8A5htbB+sb79qMdK4zzt
rzTBk+ZaecJ9/wPz75yKzdIf98muPugn+bOdfLTzPWwZBJ7kKqiQ+jRj/RRUin0pJxgDYHPv1rZI
pliTL3dce58gpUhBu6rJbAT4/5m8tgs1r88lyMbBTwO1kJjucRws4Smjeewon48iSXii34eBm7jD
KCdVT9+efHYFNQ1OSrkPyuEoKEMaPyGNYftc2d3Tu6kGP5JbaZ/xLobNzZhIuUn/MXWMKBD0OZhr
W1sjArqrTm7xdNsTchqZQ2iqdbH1TkaspJbaYNGvjerPSW7QGmBlDB8pS9Eo/86MbZDijOiU9NpL
7Bt2pS5P/f0nUq0BSrpbi7cypFbQXAv401CZIf0VrOTvqLQuXSgzEQTH4X0LhTZBkMfcttPjX1SF
pzVmpXcwrxvnjUyI7IyKQT7ng2EngX/j8Rh29U/WWz/ECGHApHS0xUw/eUYN26EXgnk2cNoPC3KY
5rCYm6e+9BpXmzc9JzBrlFAHa0nXam3MBnmOaHuXMywtR4fAq/23fGAvgZIP96B9nQN51ebN4H3s
RpEmyjYkTr9Jeu3CzB/QXDjQSldlPD6UzuGyYhVV1podlt86SZbY4y3oJgotH5A5L4+9cDgCMLkz
vixvv0xuDBx13HaVEA97gI/ZXT8MCZaYiLoyweVkrM2unUA3YnUvGGR3A/YH+w1Ay7od8AUe1qTx
n5lAh/TKdtVqHXnV9JQpHVrMEczL2u+2pI0TZ7yc+uVDA4rqvEB4ni6yQtFM7zI5FSCb2+r2Kkge
r5jzV9cMeaaI+RrsTkYgR2+CEHU9BD30rTEk96oIaM6l12JDCfqlh6rmd6hnmNUEYmUNC2oeE2EX
QEp4LECnxPYc2ayjr+9X2GiYdHSShgdoFMZrRo3WSg0virWgQ4OzL007prBatvnI2hjgdaYixwM3
6TfUcCO2ufzDxFedrAFGA6WND1NhyiXjFMIO91+FNs8cyna+W+ptu9acaTdJ0RvrCCynJdcixzZo
MQ6CQnlJfu6aL3b3PeKcQeZg9rX7zTd9jEN3itNZwaSNTcCOZbpXkzZUa2dIoxfxTOFNCtYhPb9i
voAsDdD5GQdGeeGJ6jQlmB7Mitpm7E/omYGeWoQ662B6QULsuNsrvAPe+uR65X9hUxLLzuDyo2W+
Bnqo33/lwedLwE2/7j+7Z+1Lq3qDMxCOQXEkAQMN6aJpqpO99+n7FUzPujGsAUGcEATFaQqcsmHE
4Xc3HZ3j9LbmOdEt/3necdM92gnGP8cCRiLWza2EXb9Irz4QStB9m4dZ9TtFab9OERvn+L5obDit
+ICqgBH7UCYMi/aQlm/01jN4gCOkjPDGbqe0TaF70cmD+rEoLybczgr7x9C1r2KtFab1ljJyyEvQ
KBuSvugOkZvjKmeNEq+j2Kpwq4IRQhxWSOhivNSUltaSn05Dtd1/V7MAkIEgKxEln1Sjqdue4UGz
p2AgovF+NgIBnKBNMA9ynzj0090f5+GfOb7sAvisUi65ChUWm6X21Y+dRlEOBqRQSgvSXdWrpzAE
uNXhRf1Jm1jx/Znnv40M1zOpigo8tiS2w+zgXBIB1V/Zkt7iUWKjr3C1uGd3wyWeJt1+S0//nKgH
xMBt7bgQPpvaaw/FncODoYuIVxN0rraaruoK/flkgVTSThjkPNIEEQNoT94Yq67RK+ySsRW0oo0w
Ro06OV/Wqorhj2sKzpV04VSJTvGAUjdGJdxahCX1y5GWDeSIEz+pbQRI4pXo5FcciwRpGhYGBzDg
vQOcL0bJ8k5NdaWP2pnZsmiHT9pvDqIg+8FycfWdRinH8bCnYfCCKJnrAqJ+eZ5D3byZzWdxTtcY
yh+kGCrBiw7qNpMrMMND7o1Wec78GxHCimJWJmhPRkEZ0K8APvc0lnSTAe+LDo9UiyazpeUqz2em
U64O0ZWiq0e7fzHtgRpSx5weWHFSNCrrYxADvu+CEl/Mc3iZrMq8pZx9gMTZ9BfZXUOCOKdHkYZw
WA8GTNtotago2jXgKMTG/k98nRgWq9wnlZSV2Qvg4tYHx+bUUIVnsjuR/mZ8qDoKbE+99q/f/Q3i
R0LvUu3/ztp9w4xxlEQOrOH/wb+lRVFBOtMQGSoItXfHvBDg5yYa+A6tdSP3J/9Voto2PiB8P7wQ
qV5LtZmXKRHLboIw0xMpU8ZOwqjAEtXhj+3FqTbXOMR1nyd0vC+1r1moe6vDNHCqore4ZSqGAVwo
t9e7jxUPe+znJPxFPbe03jd6zsA+tzbSu5LzlupR1TPknKuu2pWyHz4leMDWTUVnAfv8C0queTIX
HMQpL7HU3vgjOhXYtNnZgXifmsF0w5rPk6KjVxafAE7x+w+qZnV/xaoV0OLHYdmGD0HQyv5yecMS
doErM4IuktkW0JfifZyiTCPrU9ZiITcPG/p2TaJwUXg8jG8geFR5ZECnmrwLk8qOfx5zABCGDV3v
tC6B4PxW6LVD3DmS/jJDAGREpmoZ9bHdxH7IZbyz1hC/vizUCWhAHLyI1y3QNkg9qjaeb+6frbkz
Er0smqhBo4ify/cGUMWBZKTZzNi9pRX2mtVvGmR5EO6Lh4i+H+K9uQI20jjeKESyF4/AU6VmawfP
9TkR9UTp0thOqU3+nN+VjO/ulUvJzCGjRvh6Z6XT3OmrWpUMsTKE4ITMGuaDw4XRDJcz7GYeVqxQ
s7LSNKCcKsBJFDW+2UA85a7W4Jza6OWJJsDiHvGC8C8zRXFOKuXYqzHYS6UpC1zYM5x0SAGvdrUQ
GqfyydIOZOLOldQwkYo/+4F2RPVqPE7HCIROa5T09AGCX3AgR0qFsSm22Ao5w2r9weFNdFcYSFMI
DtZgEp3PVwr++3PvAtkR64l4mIMPQC6gMjEfe29Av0CSiq1I6tt/wq5L+qFACV3BWP05bqvsJp8o
ymKIJYFxerCglmQ0+VtqoU5yBKh0HYA7VQMXZxq3cZYV2xppBM7Yk7m8gEFaXCJg2UHRf3XtuC7c
f5q0bctziaXLVRHp23bUj9LqqDSv8TuvNiq1JVD17z96y2N7kjHQLivQXaYAN9MxXa9KO+8xtXBD
YcWvImymUztlT8K8qVyJwpDENDXQq4Il+JcxJzq85AaZ0OdxRcetFQOiu96fpKPaGvCW2PegWCf0
kvoC+858m9EwnCzGRURdbLG48bPQqiJ3V4lq/T0iobFYYQcdq4/8C1xT/zEu7XEza6R8/N8tVCXF
iAvzpuIYIulxk3piwBVJEXn0m+qffFrOY44wgn3I5+EFhBdfiofaMh9OGF8XnNzP8GkVvF2yT9tV
RTx/RJ+GbALEikvbRhULamo+8694HDLO8c/y5bcfceXsk03AMdQDw6K0p4V7Ce/1urvwJAOshps0
OqYO9mUL8keDHatYRLUeS2O39oQ0RGrrqoJSWOm6gNw3JjCgwHLjP5t8N26SaKq3+OTT8/3P3p1/
wNClid5a1PUHdbYWqKewIO9KLRe2344W3kwzR1qo/5Qr5hZd0c03eqgNtlgRJcnhXxQ1nwSi4RH+
MHq+GAbEgXl2coAm56v3kcixh+GfYd5JagrCsydsErZAE60V40Bng9vDcQvhkA4Wb6wppuzOd83s
JimCjnIOMejcQz/4R/B+D91yu461M6giMJgkEKR84vdP7c+LoKE+SltjRyd/U7WbYAwi/r5lqGwL
h9gQV1Z/kvKZIU7djQLT7wqamu6EuqqbRvJZbzGPJmonxvVUx8Sveqzqy4+DealnV0jasamhPBHa
PO+lFgXJ292SXMPySGmZjqS+LWDVLaTGVMDczVii3cC0dTfHXgvEwDhilcOUjMXmD+LuUGC4ghco
4AcBza7r4RLIoBsde7fjL1CML6/RNH8IH9LbwC0mpLoDLl4B/eFhEW4kq3+aWfLxe3OV+R6PROP4
E+r+46K+lYIVRlBWMWHIt2ILnVkZODSILwfvbSaafP0gMhqkaS8u6DFO+eaDJxt0o6aDvPGza0dP
RXpagVseGp1QPmYJdHaPUegY47d6oPlZaCss3pInrWoZPlQ1ZmubuQ9E+qrCVaI1sFF99e/S2dT9
F35sRknCj9O15JpVgQYJhbHfK0vv5FlJrUD0ezr/RXy9YXRLgJDsuzzZjUuC75JLK+wtO2wTdQBC
MyFHKzcdb96GNNS7/kXLmWebuZhUYCjZflJw4Grgstnmx9OjBisoN3EVNAeJITeXPtvuxpg2+bnb
gZdG2hP0xwpLIPzyDQVQul+vQA8UOHfVbQ6idUXPnm25FtAEZzFQgKzTsv/gMJlUfJYtuJWuIckX
ay+GBjnZ20TlqJwZ5dpvoVv3IDtqPnAv/IZGTTWB5MT5nA/5viZ6Hsb4mXY8Namh0xWaYf/fEoX3
BI3ci9jNdahSRiRLr6sNOKEKs2qa+927cWy6kZ01/71osHHy2L2WitVH+3qfTgZWrnhn/FY9YRpQ
DK5uudvq4Vrds18tkxJO643ev0SHl3LkojdhI+hMm/HYUVssbRvr2v4BfNDVZ7mJfgnSgi4zSo8M
QXcQz0edaIwkcFiX6QK0PhBnbXEMDgXZOBxREBq0i+hjh+rYpfTfBpbeKxkr32n4q/sLPKGMUqtU
cnu7C2R3cUKGZFEtdufEwj32jUpD5yXdS72Kx7sNqBeTubrWr/ok6xUwm14mTVnHb/26HwL59B4f
ocjJfd446ngDg1hcQTdwmd+Ob6sg4rHCpgfMIAnnGK8UWf8eYPz1r+X5BW5tPUZnFU0fpxIyuQhP
Oh2GCqUME/SOeH+7WnMYhfXevGEBK58RmctZ3oAFE539VSMUanpEyWaCJGns6pZf6ktYgCJnxmRj
XJdBxH3pMLf58bQls0HKbscPV4RSCBRG0OqHP4PbiJdZERC/8muKCJjWakTvY40VAOKwWtyLQcHa
ANhDqz48G9Qmt2cQRApZeSoMRezLsRh6ClIcx5i/zTpVkyU7A31HH8NCjF859Nx6ZPObzx7789Yk
BfXhoOj5t/DkgUiIUzsuu3DZjofwxlQPsESRu34eec0SY4nY1cfWY9SLOodDDQrj+3BrWRzmw5lu
HklyCGXLRnBruhCb32VV/LLa63dArCdUu1xr6xfJA3NfaeGUd6gInMwMVGdgRDbqKl7+nhUm6K7i
f9iATmXVNAiJtMUV3oKirMd7QB1Hw6hkupZP7LntMTU5zGoFo9E1ubcWyPXk6IElLCmpdsn10tIY
Z5aRqqSPcfxA65kHzy+g+rjWle+BtplfxGbffYSPJQEbOBIRBt+nJp21zVmtAe8oOinEHahlY8zM
rT/jPm9l2yLO8omuM717Iv4ryPytnB/puRMpEtOj/rO/H4BxGGh9NprMtoI0sLRVA7SSE84H2opl
Dt+B3YjGgD5EbFxLpMuWNsb7G9LTGF6dLR39ooAeEw9etXONDYyQYyQC/q/6TJknVG9WZGDNjSQB
WJDqnc8F0GgJVHxfOgcrUvwjjdYfzMr1m7syM0KtmdKAUYBXks+pJAb3B0mj+1nyRze8hXIoxUqK
vGj3C153rolfDB2g5l5/VmUGhi5QgExvV+NZi1MyXUb0/85Ji2KEFYW7IVp//Pug4J5EOBe9FkO0
xMQUVge3/efCARr5Ej2UEIFdV/y3dqOIUDykisvznkw/20++NcT3g4uBTguBX2oepYHQbjsfW0JF
FXuxenaXFmV8ErX4vtuR6dv6/Qv/ktAQXL+pQK1mLoUhyEaRfMOEiD60JexKdJgYdIk7muI9cbRf
T++itM3jPTyKqL0dawddyocetfiPj5TX+bvcIKsFwHJ50qYRdQf0KX/dqk9TrYzex6XZfOT1OJzq
sK9Ot+T2LVDxNqc9J+x9aQJ3moM9Cdzk33gk5aDrww0ChWGRBwzylxmlfZzITaEdiE4llcyoVfMd
GXQW+EHPYSZEyPvzYaxXoLV/OB0QdKhIdKSQCn54JEsMvmZIR+WI1lbLKRVcdW/t4MHDFIX8frGY
7AwNHwOARmE1/F1rzZrzXVL6hRay667W6vTiN9+r5ASXoawKIZNYaE2CMqe6NzHSTJzrlVlSXYsB
EZzVR+m0B4oLnRcZBcx7iOThDCbKDSNVLaM7lYfpaAgJcKeZ43P7l1+1YwT3sWN+T6q6LfCFSeX7
WcnBtuAo+4ixHzUllSD93I+ZlUF33zb1NWxE/Zro4VIAZuDcTe26mVSqxmYGG6/6LClS/O+5hHNk
Fgl4QtVeddkN6xLB9NH1ui2Qxz6ieM6QLJIFq4n301YG4DvGCIE41cJmrGqoLlrC0iSOIYshNoV7
oyTspmrvUw53q3ZpcWOPKi3I53XuBfo5Wh77wgyZCaUgm1zyG/yn1ymlhnl1uKcvj0trEy+fcV2S
8No9q7iU4tbfoxvNs4A+70izomkIxSoz0m9tzRhJht7C+YcDGP9Nt37xYpJH+Nrd7i+H1z8hKeHr
+8DeBpKPA4xEDKf/LslOiqpjxizdLm7nFxkuRccYDhJux4/4kPDsCBK8eU/NMG37PdPVGrSXDLIo
wkwGppt4r4synWmcvP4Ed1ewqhYs25TpIXDbWUBMp5q+nSnEjxMOkQ72rjwvw/yPlNcNfAK6w9Bn
RoNNyDb/LsRpn+XUN/jSWKEXs/QZ+viRbJZAn6FpwfxjapCsHfR4X0BXNH7bapSvp63grH6dp+4D
0QCK6pze+RMIdSIz/2H4rJz7tppUD4/kuQumCP7rWE0QyoHdhig7rQXSZD2oasJNUoIFpVB2xNLK
nqfLZWpebq3Hnk58qauqIZp+/TAyFLXY9GO5/jvXsD9kE+jOAUtW0BJodITH2lmsmiDH2P5tn/jS
0QQ2VZVAUUxxB2/0sAjYl2HuMRu1YLpBub8U4rW2mCYZMYC0Ko6SUX2w4nCLZCxpSMyftZ7fvBc2
CaxtMlLy9YQFVSeUndx8RGK4FWOI0tqnB+zBj1dtlhjdxcwEwg+z1+VnaJP+B6pxUE1AOylfocgm
erMcsSrNbdEPH0s7AGwbdFTCa0C6jffFtKY5QApagBctUuvOT9FC3Ld+vUGN9jo7+0Q+Erkwg3B8
WFJQUw5OQKnrQ7w5b3QcAMMtHVVr6gjowfRE+GLZr4Lz0q6HQpqD45FCQ0CtWxdNvezrRZnky9lU
Qr7Bg8x900BeBS8h6gaKSfLuOcgKK3oHMEnA1oqDV0MvDF/wCj8FMdRWWJqQsUYuSd4nkw75iYlv
uNAUr7kBBnPkOxdYdK43gHuUS9wHGSOs+ZIdry+0URpHC9diE2Hf8y0uKAUrUOP9G4pfB2RS1W4X
rLXG8pj4W/xXGV1pW0B9gky4TGDoS8qnTF/RMOZBw/5zZn4Fz1vxr51HI0DQ0wRbFoZnlQztqtL1
m/RFfGfzshvo0hvpXcp17Kfn2Obwo7biXpa18M3tvD8+/GUOGQSRwPReN+lc9nU0HlYf6vMjLdRk
UOwE1lsk//pzyB576S/kLGoeq2FkeszNk64bEo0FxtpcDLtuz3wdvC+YaYJrsuTLbvX1136Q7qEP
5Kle7pVwOSzQv52RUejxBmQomUXLiXIbjXbyeq5BCiidAGWkJrxrkVtzo1X9q0QW8xaDBBJunqSZ
HeR1wAiUevSWTpaZX0LFu5IxmY8NvU5aF94Jf504FIvnIEFqY+ZGfQY0VKYMdtlI9SLW1ot1LSTW
4vi3HI/aUDBMQdHzYGD5dHJq/C75nid0A6MRXQB2j6XkYLSCgp2q799GE0hCQK2qGhi8ndw6WROA
JnCetXHrRoo0JzgkPKlPcKoubT/UVLWngqwO8JvWWjlZXKlC5SHqZvr9l/Z3aMusqOtXMnT7uKoV
Gvmx7nOdeO1S/942xrj20HHfLT06Az/SqyJ4L9ArYFglHjCQFQxUTiX8oQhLRcZfJZOGLlVqNH9s
uk5OowGbVN0p9QAlx2Jo2Mjc1AaDHko1/z3GBbuvtfYZIk+Ci1fT34VJJ8IUIOaWwQepJiUzNhaj
nC1sDylVBP0RBqb5/HKk3aLHF0aE4+1NSocTqeyfhnLJH5XvYzhmZ329HQ3sr5vQWOM7yiEZMlOd
QwVpBElKr3jXh0bh7M8OlX41tou1lntqIUW3oryBRXnqwPcikEaYha5AME3J/0jUSmLrs4BPDxRR
+f3a9w7Km/Mm+eoCXPRb0mwHTSGmmYbQstl/lOS63OC3XAmla7SgqaCyXt+k1du3Zb+BmLG5bW4l
hqs6JCkFgyiK6CwLVGVC1hO4RTebozDOROEQycUMrioPSOcnVzL0Htj4eJbVFlKdmXuJzWxsQULl
k5Iyzf/tPPuwZ5WJ8TIBkL1tliS4DWu5Ogurqytgn1j0YyegmmrOOGnfZkQsIXOXBxrRMq+2b94T
MpN5GcMOII6QgY8yBCEDECbAMcufNMl1slU27Lzb9iB6JPxp+M//PwyNIrEe5kURQCMyeZfNXeow
DkwquwEvS9wgaOt5kx4M0yc+TBTFHXN1uC3QRfSDwU3MQw4ETuzSV6WnuI1gxugFJUYQurLpWuKg
hJJVNPC9QxX2V/naZue9sSJhe+LyRbliYU0uTT5tnZISxfCdulKubbZRxWugkVls2z7Y1mUE73HY
59pfNzDbJ6UtTfbt/wLQrOD2e5PT6P9lDz30HPIdRJMYM6OwelnMTbdHL+YIh6nO91vG949x9cby
fEB/blMymkEeu1Wq/toThXxIuwHd9r+I5aNKofDFXUmKEinqRWsOvyoA3+yf9OYzLCh4vwM/70Mk
PPfSRpCp7xDQRiGHtmFtos06xlwLEhDRI680W0MWV/nX6O4rPjCRdp5CbRGuquCPHy8PakUAma1V
ET3qWx77Depchehw93fbjjZZ1W4pkGTkJyyTW38kEk+MvcrsFoliI4EDXUK4wvKeykKF9LbN/t8l
ceIQ/DWr9J9iPdREyoldexg+VEuMKQIZTOwN5YVl6jj2tqSBstRrgrDC+6B9FL//KakcEJFT6DTm
uZcncTtrgXrhSAQB2f7KilN3YzCjTxT/6KHoAiguATJeJ9enWY3DCvZpLVWJVELRSJLpUPbuohGy
WxS42nUZJ0YKgAfuq4gYgPmbquVaIS6jUCJP5folLCFBOVKRHB3cmlRrMGnyofrfKzoJh5ljAWW+
z0jO6mwJ+p2prxWWbwLBpINqDjzMWI7yXsn78Jg6/g9D1zkUoBJc0CUTMgii7xACNjHxM0MJ4VXf
n7LcmRBSwa6UFjVTahQInvprIio/KFcPpapYj7sSmk7/w5OpBBUZPQrh4gypariSe8Jj/lpVgQDv
vslZ8jqgPCF0apnOlK5/CG3BRQisCYMLhSEZYOqiV+gTTDwAkWMk0SVTYzxD2/V/mxHkf2whdNUF
OI0qG8YQY27yVfmLgOe4ruJPaE6HpYPGKJQsN7aZbN6SFwgKd1x492Fz+YmW9x5dSJxEUMjHfklp
eIggv9eQ9DHobVlJv++izLeZ3IGYfhGWEohG1ln1tJNiStibM2fpR6i+o/0pUmb3g/n6uNCjJ82G
ZaW8qreYpvnQj8LHbPqjbmXiT04QJofx0TWeqisgyhpSzPpHPr4p5xxnKjGm3eIl/vjpD2yyWyfY
KIoE4TwA/dx9IeLipjLG/jiVbcC63j2/Nynq4AZYnmzNjE+Jm7o1wZKeE6yZL07OoKrBaY/b4R8h
BmPq7VUSIhvLSa6IqeILpA5ZagEY8S4oIA63UiAsJBIPslVwJn+52fCoIJOo/zTBBvIPlTRPSYmQ
YWDY/PugVQBHvdwKCjACei1xr5/JU3ag4DlHA/GAuAEnyoBVgKRumZrrhkZ8XQg1RTA0kVmFbplS
lIgwuMY76Or1bAZwNLjhHJUTiYMC19SWTNDCmtaIQ8saGD63vRYr0Wsu80AnKxiTmcEbr/oigEsj
RWbi5tg8+IVtog0O3lANT/RoaRRPYfUimG+kCDiIvA+0nHAu7a967ef1FLURW+/Q7PhsrgpFCUQv
FTg6VuZaRG8SmP8hy+Lgnq7qSUxjpJwZ97E5Vfn9h+n/xLm2A2drM/GRB3rxhxqfbOMxt+vIBCWs
5kM/LYzGF7/YkDhD2eZGZwBD+pUR7FZIgD/vY5b/fde+tRW6Ekmm8tpP0jzbqsbG4UaDDlxQB4nM
srYhYKo0wUD6Hb/TToCal+QuAV+LB9FlpePTCg2CgDm1Il1k+caCIMkQR7ai2PA3alcm7HsRpMVY
Wb0EbRpUKZvy/ukRvWdx2DO1WSE72ftjNUQVB4Yw03+3MLSX737Vff93BaoD3hXDgPDa8TVFCtVV
k3HesSWSRB5iD81I6PKvDsLpBHneWa+VivTARMyMlT7RtV/ZhEPYcTzyUAm3TIXdqnuzZvP7trmz
Q9w0PPD5km6flwvMxb/v3+dWd5EZdvAVfij91Wz4hcCz5cjmJ+0sU/xFYk4qkGJ/O6EGYSTbqjLJ
GuTWx2WJJyc9rYmZuOPbEMQg0w3au95t3uRFh0zIskk8EGpBk8G4d9paW2CmMGleuIarAdYFPnAK
tZTwcR2HWoy8FgER5D8avVT9l0WacRGm/9ipIAyxQy2u+bIlnD9DT/DUbcYA/0wCPhMgLQ8ZuhzH
uApJ/kQos6VjEVQuM+CBIB00EsZenRDv15C3vkkQH6EGNf19VRYbMKQi7O0OuI7M/bHf+92apSD9
8NqyXuUG10FPCKU9yn+G5mJRdh45QRyp0ngfM7L8l3bmRpzNDawkaHAuOYnaOhV05hy+toQGj87Y
yvTZzUQ+xOJNPhWYXzLp5f57heMBuiFDxhy+Mtk82X8PlvQKkX8/8ZdgneS+aHDXbh3Q2k5CTk9y
m9dnzwtQ+eC5efhe12+DK62a1gXjTiM4D+1ROA55wOunSso6E91nZxDhizK0olmvT1uNrgzW1xP1
+hW+mPvjko9Wheg4EzO7O7+VwKtp2ivX3/vsfEyAnFQIzdZaZYQ+O1W4mQ+lPbRmtjUcM/hHlRZF
qE4Xhtcca5wfVxcpOP/ZBCKrGNeTS8UHHjJYymFfG7n8edd1543EbLjlE2E02ueX4bKM87SVuuq2
DE2gloYo38/cfV0+pwEX2M2hLDu35FVw3tqvbg5b6ge+ELwkqKmNejT7QDiDLdStFhFH+i8CH0oo
KVbccSpoUigylQQlcOwcy2AE3FuA4hEhwpLBQQL+cTPGlixe8X0Udc/PzUBH+0+fIki8oiybJ9/s
9WLeaXMtTFC0BRPRzdREyM01sK3Fu0wWcldfdn2/R1bjBvR6ZUrvqZwyDKqKRmi2Y7pQ/4G5xSF5
Ve66MpMC630M523+4sxky43RatL+z5bnwO2+aejUxkf1ReXZPECYKq3fKYIZYQfRPRFlYGUjGRay
z1sIy/KbLJLHiIh7avtJQyOk4/+fDKGUSQnFTPzO1m0QmQiluxjx6Zoz1cuN+hIkyJTeBwUyKXbq
rBsNmlOMRh+CeMZqzH5bL/v7PSbhAuvN74AIQbiLo6Ruh5r1GWyPEV9kTG5pQO7WbER1HFErNO4z
d/2fMP4QVzJN2onJ2qaGzhw5vN8XRArIdKfCCL7GIYq0QOJ2MROG9RI2OobqEUAoQSj9aOU3/k5D
REvEgQr7vk0//vR5kX7nCrAcQeS57rbR/q+2re/NoyfyOfexJx/ZvzXXip862OAUzOW0elk2mio1
t/lsIZ94ytTlEOlHeNDshGN8SqiXF9RVBDuicSt+GB6wEA3IeKcQhec8umO7dS3NvIdQXmwcSIiP
VaDwVx/MBi5NC7smWxwqWws8NoQNTVX1oshQwkJchRR05rj8mfjXICsR1KIEXu4g7ViR0E0zVUN2
fJ4x75BLjoSEAUx/W10o718pgYUeVfhrQrxWB0OHhweQ5eKFuEKJwq0gMNuPm1IdXZOBM6kcTEQZ
qeNM7oUw7bgRJsfKQa9Yhi0z9QFqF49lRJg8HPDFq8JjkUygOJGf5BxR5SJAdNj7Uz3r6fU7GIcZ
XkbkKSeo72p50mWQjq5IOJhSE1IIwcK9Pk3qUsjgFEIsuAJEIv1PV6JlWWCNtxlzuYLXki4g8Wa2
foi/qTixW3lqfgv65wxmrZbwuFojdDLcfJ1sysQlxoLPsGoeeVSWX3NxUm8ZwZLBAsOS4bzymny/
//eytpSkBtRvliAb+vGc4lYUm9HIuPrUUn0VdDVhUY8XyC79t0pKFnZSgMd0ISPP03XAcnYaazUE
devscoI/zxDfs0km1xgsr9Za6yfXyj4iXYqL/U9hq/Q9rCHFIQ7B5xBCVHpRn9chFpDD4FFYnvhq
RZZM55S71lCQjN3yQ1UXURlgyXax0Uum6W9qM7KlN+PlahakiYquP/XbN5jpRSqJSKAM8Nw4QD/r
stiufzKSrE0bt/ibOPKGl8yIHCkJgb0Sa1bM8TuBjBjSz2twS0OPlyjmfkDIQhO0Ee2Egm1H34cc
LOpN/tP5sjz0ZR3MjUr8qTPVjIOzYpzZH9r7CEKB+Ox5OrDDb38740xj+uO9pmYJ5OUOjgOre2dW
XBvV1hLzVJmGzEFqE995m8MhBZ+bEwWC0nSeHg54GeFKZF4X0XYGwQQS3ik5CMlu0dSyuXJW9+Rj
Dk3BYFLnGvntU15DoTXNBhTEcWXRNE4k1g0mhuyZMMs4MgbRmUwCNIoVinknUc7zcYwYRz6LohtZ
O9/Pj005ZnMNa+iyFV1zP3n3h9/7LX6o6f+PuuEn00P1I6DYd4YMU6n1ITwSJS2rS4e/ODQjEEEa
/LlzQYT5AM/qXrJ+tr/xaQXQTZrhyNc5uacsCBFtXd87BpwV9t5aWTjgGGKpCQT5lxlINN4txo7n
dAfpP7BRtEzp1bwV7nIMvRd2c9D396kdwHxo2dxZ5v6XY4WzU3jZN/Uro9dUYYXi0SRekaQCXc07
rv9mOS4XY8yC3TAOxi5CIvbSzbf80tle+VYDjLALipNGJ4IAQ3wOnj1rMWwQuRAOU9Gu5qdBXxG8
rYPpgS6MKCF8s9wfp39NgDovhvKtKtUrIRVENiPPFlhBNO0sfd1Xn+ehIRDkCxi4Lxlqlbm2seMg
xG4ntWI9lki1agwiilyvCcQEIMIULEZWALtfc7QbACUoU1aTc3JhvOGrxeCOYiV6xFDyj5Ny3Lea
pq+0jirmDmRFkx+L4jAVkRNqBjEeqdx3qCVKGoG8IQ3pBxoR7vYomqoYQWM9deVJSodf4PznAOHw
I86lJwWyw2ZLQzqvYQiyV7x8qjczv96kpT628N5QxVpkW0YGMvQrPXvuvg7masQAmELFmNhwg4Vq
/RVaJa1kDIm7twy7YWs/FGXaHOXczp9bGkU0wtBRazGHCrSuPr91UHB5N2DPsQD4EyzpC3ttP7u0
/rOkHgvL2jEsl0XATBA6WMebynB9heAnrA1XPdOvurDpVj+d1dnftt8EdZ1LPghmCfYag2gLiDx3
1Jr2MURd2ANNImqzZR78iiez9BCqCo/+it/BGCQXthB0IiqBdgwZ202KpZyu8I0Yrqc0fox/zbL0
rLB4bwhvDn+1IjUZvp1mLpUXIsz4jB/dC52hOeETZyYytPwmX9NJaxoOoexCmxVjd0BPjJ3u9lso
nNJobe7mDj8VWOkg9nkkoqN2BYNSUhedni0Kyl2f8L9VOSDCJZOuaB0G4nAWNANIAwpvX20x3h56
YPX1bpl8wlZhdB5nQeqb+A20Zz/hLhxskHhb3tfUeHtgOeRusMo+MJKGBseugHWQXh6j+dsXhBbC
nbc9rYDkGb1YwfARboT8wOf6Jcth857Bq4qX/+WB8DrYXqp0lyk4qe4beJ8EXY2zGEgBQHdO2nVn
RCsQ2aR62MIH3NlUKv4YtNnzUtlFu1PveDCs941/lQFr/M0xrob5WOBeD7c1ZOUDVWD7sDVvY6Kc
KcYk06uk09hGAEP72onu64udmt8jaHx75bmNvRLN5pS7s96d1p+x3Tp/30JhLYsI27LZElgdvOQA
BsQ4sfxe3NT2bnSuq2Tu+Yj6rWLiwvAoX/t2GPw/ebTe+a9rkFTktImvvVk2fyZcq+ZXO+ppdUf5
3py+332TF99b2FD9sG/cBG+V7MEcnh5KcOIEVkyeutgEuT339Ow/p4s/7pVb0iN6ggPVdctJoSaN
H7ikggshS47/YrBYoo3sRUMqnMHpTS9mtfzokmmK8tyMUgJDmDnb8Mxkv3ceK0eY/n6Hc8HyxYgz
jysPLjofo09n25bJA+g0SgvvuNXtt/jtrGRuRbkisXmcrwkEvSVlors+nXh32CqZrAuJfC7MHZ4P
c1IM5t/twZQvnGe2+1XqpjyLDC3tFfGf8pi+suDe5YANxtLkpLrQBy9Qi0oTeNhyBxw4a/c0q/i7
xO/R6r8NrQ5eX1dR4mOG12B0hLN6aIm3Z6mWtRdb4O4rRuwBuoUzkJ08sTkQsa2/vkV4KxdZMKJi
2FTPIqnnb2mSvhPSBh84CBjbPFfpWkflUwBnXBQQ0AuahjCdSgbxrFL8akBqRyBZNIwGsjmLxV+J
MQrnOVcncR6mX8ApIo57HLxIAai41I0HoWc/sqrYYez4s4XpmxDXgclXL5NSMvDCk8QXmXrJc/Ei
j7rwooGeyxBNouDn+rj01t8sFjkN5eygt/rTMADc+jM9jh77PBUOcoJt+uKYpetybyhoPtMrfPQG
XdZJIHMVLMlVU+x9+5oAKyupzkGdIa/L1t+aYoC1V733OrfZ7BvC2oGtLgZuTCgardDud6GiR25I
2UC2XerElhpJzeqPJerWTjHNX3MjIfVmtBbTsEPWXR5P/uJgRU0Kjw+IBQH7BZbcjdTaSrPApd/U
+9Eiop+GmLYOtr01h04n/lglTffEoBpIueJLmdtx04LmjViTriFyBu00PAo6Kvj179rwby8KpcNL
SMlWtJFGLnaR2jQPyN+TNZG0bwi9/uS3LwmT5K3RoIFBhiYjIsVQl1ZNOyUdqaViXe96r1c0nbfH
ttJo20V7jxSLdb8XNAhnGyo3j7TtOXY61v+PsrGx8W+A+0FVYggGIdeGL4w1T0H60P1OSBIOXbSc
BoDu3SU0h9qXzzxKoHRbX7X3sgwPKUnH4//2ytiOjA5t51rYRI4OrP4yvuLEs9Ywt5ImOcyvEwUa
h6TCPE5U0Ukh1J3biTvSuQtMuUzxft8pCuGLBREnw/Ija/dS8BwimZIuGwZ/2jsWaPyuRjYIBQy7
0TSQ2dHh15lSQ/FEvwXLGiJ5kUHsFn8YvNNAS1wHLfu7w4pGqR1B/Q5ltT8u/RGujmvReCAM8vMi
/M4IwQ28KKaZloS89kdUN/Si3JnHV9D8SUed5uemgcg3lrlJWRX+4JrVFyWCuNIoEfLJDAAUSX4s
E7uDxZcgjeCb2cWSINRlFrchKAEDmxGoLNO73dj3qNsa85jGYQ49F5mpW9WW/Jh42Mx/YK0MGUQm
8THup9oRey6/7hQ5do0GAJi0WJR9cVcJwX4CagJ45LtgrAJAFHLSXcITEtY15e1LSVmTvB3GzJ4G
wuN+FqtsJ2rCNDn1RiQZKIi5FA3iCkCAqBQXsp/CfYw09xUMXp9nLX3l9BhJPeflKR6WCk7sG+ea
aP+a+qQzslChB+Tz6ZMhq4wxAu/z+fQpkr3U53weEH5Bp9ZBoqCNfb6buwjFaVi7bXYFmqXfA0gu
lvczXECWqVkftOfRk+cNFzI2UxDspaok11x0UGRugO8QROo1z6sBkjU05zkWA+JgYlPXPIiKIiuK
T6LOXUx1mWdwn34flgmzbc5RSC1sxG9a+FC0y8atuHydRruJPu9VU9WoFvMhawqvS+OVaOj/U2j+
SNwOwiIReqYsp8nNQEftJXmNIeXjCGjNp0lfrhdDzQ0PXyNgcTalKILvtyePz+AjmlzM/kxC6d3M
+sCEDsJZ4SEPhkOcwSkU7naXIAdFDFRPyk6bj3xoWbRPIy0NpiW+IBoF7T1HEsE81dgFjwQwnny+
FnQAuuKorzTt/vdHBhLHnJs876Ujp/jt/WVE1chpnRVtUWS6A1ofFtUAUPz8RV+evGtrmfm0ADtw
dqQnC+z9FEKVqIkGbU1INuz2eXMmrCnQWIXoZiy4r8kVcEdWxZoXarfMlmOd58i73Lunp/cpkObw
GQppId/WFXSylWsGnys57PaQ6Z1hSao7KHwFJqZ9ikI9kHaYgFkyAJgElbQDfKkb5Fu+Xkcde2Wl
YPFQeaXa03IeA2l7XSrtAGosnOcortrA2fAfSPVx+cJmR0ojRgJa87CGn6xnBkiwfMkRSv7mcqds
wwQHyQ/tazfEtHZG+Z64mMo+Z4qrDs+sTiwCdl7ARNiuk/1v4siwbHDSC050WfD3pBvbW72ErIvN
DkOFBtihTXyTHhu5YBvwDBM5P5pUiwSf8w4Ys887B/OmKos3ach4O9QWL7hkeS4xTYykjmVLg91h
Wfs5LCQn323YdeNypufaYlqdaBRsETvboiPw68QzlBBhN75baspUG3GsW8qbqUxoI16+MBi4aP9H
cl9IbF/hFuylj2GPdHq/xg3Z34zH8ssnTcFBoXVOhv7Tp+GDbdsXD2SxLmxrvq5JJ4dFWHVmwx3W
P0J/PkLoJg/eolU5gK3fgGhHZubkrSfuFQA0Wqxp/ZkUKhMW8jeSns8nt9db/Q9R/4o7tZc5UIxU
WHeZhX3WK2WLBot7DIhmuI0LQI427rKKJEb1FTJM0CJdGOm+wjZz7YDQky73npwbyGQeWtHxYLH6
4+Qfotlc/CfV9UVdTN+JJuOrLTN4EVSAbQWHllYBx6iQ2FEJEUUbM6Afe6UiAt3XalxHU4epVpIw
9VyqqdyWsNgair+vif2BZvAkwH8NvZv4xyyrLS+ePYqCLNB+rH1tLFf4dstIjLJ7Pm7AI3QvwJiN
nYKp9iMbrUw5ip6kE8xRKR48LgJ2djWUTPDm9gkCCnsTX3UnBco4/US6Fd1zmBx3guLBUG810fWa
sScBe2is5BmEKKcZd2EKYPvpN2Akxw0oy7LOKy4TLhM7291gvW/PQC9r+gVoaVpJ6l7d1FlnUVlX
bLiyQFd9ioqtbFtQLpCkfC/cg32p3k7MSbmrj20TZCnzs0pLS201TAqeExWxUGwfJkkZIOhmB+eW
52tJoBwfBrmPEm7+YpsIDJsqkNoVLRB9oyznFsFfEsJj3KHiQqtulZcOFBP4qXB3UUjrfdeawEbV
RTPAq6szDlq9PqhELjgaiA5yHhhb5Ei1iFk24UgF2lbUXs9f9DAx1JsOAWmgFjFqv0T3nBJU6xbS
XiFL2zDWc2fqH5G1NRlJf2g3+mr/sqhnSXSomHQUxWFK8BcrYAp0qiThbeAyYaiy6u2k79FkcOuv
xEcmCTi/sMyyxOdv5siUS31Gfns6KvBxX23G+eZy8vnWlAYvxN2n2+PREoP3fbn4aVTCy04smiyc
J+LVJ8bj8qptQwxKKs5WN95kwVJA02kmlmI8as1+/b8wSGasIJPMUoDuc0E9WB5uCzPWWhwAtJQq
+4OVik0yFC/wzykKW1YPKfTbIWrMbNDNcyRqv+vGqIYz9zCM+0Hk79eigka/IaoO35qHmgGEI7Rd
xGQ0qsLMcv2fuoeQ8IIKLJrz/P/ZM8D2t2TNH3Q/zw4wcnCqhEQwHK+ej9TrmLWClg8EAsenlYED
YVVGJM2F5tD5k9LnPaYDKPcXDIzNXosZ6RgfX8CpNhw9TvOPpL2QFAcRhM4AkrqSkHDOMBY2pQkN
hV4WDT81SEgh7zmKXS32hLGqijkIgDcttpkBC38j5X+NMbRAO83QLbeK6/Ni8oHdB18XO2h7UH4o
EY5zLbRMaWTC14CIOlEUWILOEF6Kc/zvhwiyQ/t1/HH8sDxxpD0RyM2Mo+msa+Jx8uPY0mJ81Wv7
/ecycg/KMClBgbjHRBmi1wI7RIKS5zYgDRV2pbY48z6sp42Jg4QUhax1JQuhHQFE77eb/dUcvINb
LNRw01+03YUWq73VVAmYlAMgn5mWg0TO2XOG4QpaRFt08hPMRHMyP2T5sq3EjuUDzHE4XJqD1eZ8
t0g4YlzbAYTrVP/LF9/CRE9rMJg3+ClhcKXMRXUFbj0Lird5UC6t7O0mlftbNqflOQoTR76KMnzS
rCpPyLo3AXD0M4XC57S1njcmfRx1Dh8FH2e85/uqxC3pZOyc4Kz1lZ16nuLuweLWh2d0JNG7KxFG
WvfQbMAsRlwFlT24wm9mqGlgrWuOQTcKnmjRom8OBukM9i+MRl9AysVLXuZDfYtvayd/YbkHB9DY
wPvnhaMz9Nn99ru59vvyRznbe8hj3HDByp7niLqlMIAgidVujVH29QBP1Pve2JnjB+QKY3U90ho1
Hy685XDvzPfncag3sDcTwE/e4KAzg1LrmsvhoBkgL1MMor5YIF5fGKaVVsuEr/JbVt/egjaMY68A
nEeb/17sU5tKLU2zMqXgZ5sqtzMr4837OfF+Zb8pAtI5VHDdQZk/ZUdXIzO53Zxs7fXTChLJIIih
cGuDtLl3rBWg0r4kcfiGymKz7i+73S5eg/V5hCZf4HyXO1vjD7JEv/W4Yjyz0OtRDLzDeNJiVF16
+hRANl0zlr38q64N+gyywMOPCaNrytgzklhxtRVeuf3tZA7Z6/7flZlX+0Mb/r2NTRw0O3NNThFs
ugMSo4FmvbYi+69QIQEhkwTkADjuDub1ZowrcMQbxhg66ZxOYOXmhbVclClK7vMTIWQGebXz+mty
LjBjzRX/qDP5Ew2djLzdR0anruTUPy/OZMp2K0VPWQA3C4yahzQU/hBy/PoBJ+FL69Pw6dBnXY8n
617rEFuLecZOkeoxSCKZfcARhWRO2YnJE6Fk2MYGroQcyfJaLVaOWh0SO4eVSKAST6ehEKaE1x4c
x0VlK/H5kD30nMFg6f+ylbj7j8lvTlFTvHEz5Mfq47w3qjcX9+Dn6aEQb1XSCCwnXw5bHN1CBFmf
s3rFu+h1mUBVRSdxJbvCVAlTH5/SkqHYh7wZ80nUBWCDyEJZQ9S+XsOphuT67MBrf1RZwT+HtETd
8GsbbJRA3JL0cdRsDZJsRMgj8/dW0iksvL526aos3gwq7AJkgsROUE4zqk5t5hHVrba30BmxXuD+
jO1LHE03mv1diTbIYu7yZ5a4/uYE0QgJGbq/JbViib/ytStzZye8PJeWfDLwYcnxP9hn54oCs1KI
emFo9x1Ky0lG/um2tXTM5ynyu0rPrIRtK7tiPYyyPzrg9PVJKX5tVQxJodewp+vc7cagVOKK4ijy
91MucG2UzWzBGEllyhdmsb8QIBETaPn11UziZa/5ZNamfgZwzRN8Q+9zmacHV9yWODhkIyhFZ626
trekp6DD7d7zFcZ3iPs57SJvAempXgy4ZkEgunoXDpejczmrjYpSg8h2onUcRnoumqKP1O0xyHBj
8YO7uai4edYE7Yt5OhvtxQxa3qd+Ghn0VBitB06gCoIDN9Skhpw5eP7G7elBHbAYuAMx5xNYH/kL
YuyHxt87uaBxullud4JdF4rkmlh56G/okY7Zf5mfve0u64iaJIUwZdP/YoLeDQGC5ziU6OHQIUp5
L1vz9anFJYRxGYf5r7kuex58NV9511qx8HqWZ7u6dRXZujwXnjKIX9UgmrQ/pMfOvrMrZXg0t2Ty
xZdKB40rztewZMDRzqTh7vD0gn8WJ7AMGDVE0W03QFbhxbVjUeMZzNBbN2d2aHJffMAV13mPFglB
kQbG2vD1oAR5sRmuCWVAstGpMXgU+bYG1UrpMy9nLy6YOL5rXeh0/AmZ0pLk/WENajLoa2yAFxVx
DDySTnKhNglAMJ4hivaptd0PJWPR8AR42GeFEcbdkNyqCv1BqYdmCZawTPfByWPhM9GdLE1atXa+
0i1WpJCJsHI20W3sL/NqD/8o18QzA+s39IO2MYh+J2Ypfd/P1MWVNnsHBAliGjnF58GyFDRl4bKJ
0/5DeX8MyzxGUyQbmY3dAp8MFuDBoBNTas0uumhkMTMm5m2viZ8f2wekNgbetxFjl7ZagT3L4S6g
+ZBdSAyyYB7pjp4j54OXZHYaNYx4+qT/7ysrkjD0bMRD2fDWMIcFk6KPYwQrjpKqjJhQ1xbeJs+H
50ea0Ucki2EM7vA/DNQBj0M+q10zwN6HcgKqjf0SgdRzfKTuzvMlihUPrBG3TiS/LecS6//DY9F4
vhOuwWEZEZwcbzqo4UMVa9F0EVNODJd1gRd0W+GfiYLANGIPSThpcCqyB2vmo7Hj/YF5DkxU3AYM
BBFoj8hqAZhEYX+JYSQe5MBQO6gIXR4ZuBQOuFh7PklP6WtJUHd9ft19L5iVRihntI1IEufldz1o
IVdDvOePPG37AYV2mGPDJ06JRVLs9BvZfX+9csh6IHKuz4w44Y8jm9B0XnXr3KZDlE9KAisnnOv4
feg0UkIcV0tM2tTMsygSDHPVY5Jgwm8JRv+Ww/jWKacr+Zcv1+Qxk4NlwrAKxO4sXxPxNUCl28xn
LOYUQmzd/AG00pGg2KUXM/iImi5uLy/wMZvAexXSQbND9ugozxGz1JnNkcyXB8RHgM2hyyl7HQZ9
YdMbSrfjW2vatEFR3/nH7VSeRRRSwshd+xwDUhVf6/BtWzCfYojDc1KJSXcBxoLna9F/I5P6tTBS
kWcb7eo4BZAnPhtSHQb7Dmsdcr8v2wX74zKQCzHNrjFOLEHHK3zLFgf/MI7bNrJO4VsWSY5jMoSt
cYi4VlvConOVB4A0dS2FBJn7Wl/4UrHeMBFbNmF71ns/h+goJu0Yu7sd2bFxqhAr3OfWp6f3fZrx
/XwC91IkekDdcYMhvI8XzTgKaP6VmHR4nD5jZHaBmz2HTQQ8JqI/WZN4cFl3TObyp84LLzChSE8J
tjZ6tEDo63SA6tuhKnlS5wx4j1wpGADB7FcRCUVMj1OWDuqdF2E3t5wYxusnrxKYUv6JCHriAeos
1OyxMbYoOD9hb8POgV63ZGyo258yrL19tCEkvG2seV3SjmQUCAoRbuoMy4uvL59k/ptL6ZNmYLrX
xDLT3OHnsq2TaqI88JKZgMOBjbFiDizNGk7+iLKmAymvsDAHPF+nLr/3gDBIyvi43NN9qxBsrnYN
mcv/VeJloTGJmBh7EXCa86nRBG/xA5z+vSpwbJcgHIbm2dkXvbzgCfRm1S4QAWtMCEncHBwhmMrk
+fn/7PMOXBKE129+FgzHveqXsBf+gD//142lEBQ7eFrih3w9jIE9+j6Q+noqUjz/c46/CGRIOHJT
xpUOA1Af1Na6t6AxOa7RUEXOkpgHl7u2bdvGvXHeIINC3oKRuazc4vo4lEiHtqnKYHqLUfKKiVV3
v3qxTntNgFPNZVWvSM5hviaUSuhdmM7OIVcNF0yVmO0rtYi3SM8quoHKKezdSdHKOs7epfV9j22F
GXYRO6EyPZutrCpLVSQqrseJmP8FzqXUKuV9TMfmacxqE9qEvZOIR4z4y8H+qa2Aujam3gqKanaI
CBJDtZcCW7KBPV6qIxarsR4b7hwpYg/JCRE+O7ueDXKUfyePPkBEvHxq4txXR9uRsmYjdXczadFc
oydJMbrd0oauQJ9FwNX32PCFsoP/vv6rHfwKLI0iq90ba4PWyyt+iFcCZ4dOqfkyBAGwHcnmevzv
klZhr8QLD9I+1sb/mTaLD935XmwaC6nh2LQx5a9v2wHtEein/q2/OKT0e7L0+PXLScksYMnaBBq2
C7NOrGg1tc8knuY5vuHpIVs6EKkK9R7vxZ2zhbU3Pu1e1YhfIBMkfQa0eMd7tS/xO4RdboyFJsoz
vqnWF9a7GiwcLMMDM4e5VmckuZ5T6NPBxSy42TPb+3myGTO9EGuOQ4beA/tmSjthZNmv/oslTD63
hQBdJFxG57V2ts/LvESzrbpinjzG7OF523nY64F+NLzFApR4rEJFffZG+GGz+7xVBE+eprzbKppC
+Ft5E8TfUXm9spDCL6NZ1W0EGBoKMOyFTmy9IPE6P1AyhwjhKXWqrjP8BTSBLR5Ve8WrRv5xk0ah
kRgjpcECu1IOebwBTatUqzens8pR2WdHl4GCKbJrG+/c4kJQQh0/89YOBRLWjPy6H4vyhQ7ib2Fe
5IWnCndboJxM/V5a/nRulF4T9iL27wvrFjJ8Jtzekj3hIIKfCHaalfIIw4EXs8xrKvxUCFwkBHyz
wEKVXdgfhyfo2jBADDn6wJexnL1jeiwPCVE5S4aw0O2MEUBFL/20kutVmOnP/1vgmZfNkcLvYqPz
TrOhD0gZaUbrr/SrFv19yBPemXNKfmf03PfbyJ2JVA3MCXnRVoY7AwDhUTX2tarrfubZ0WSiOSmw
o6S8USdTY6FokkBDEoFbZFg4b8aA6kho91V6m0rVvhZLWmE+UvIY4KYGHNzowtBODsdUvQazK4mk
pwhazPRX4S0o+OIfTRf2qO1W7zRAAYwF/lSaQQ6KYcw6X9CNJqA9M3PeFeqPMcaHEc7MBaFbH5WM
9DLJb2zx2k9lz+/QhPHcRziq/6XGpv6QmUBfExeIPT6Pa5Cb4rm4fxu9EZ5d11YJ4K97DO84e0xo
IoL2HKdVIzVpSKBDWmXZV/1ZB5VqnhqI0vTu/AuZ8gM0e1iG1H8uDVir+bAxqA4tXZSi/XTWIlNE
wQcLQ8FTt9lLGhywyf47jV5hQrOkfiE2qb+jueejai5JgagYNOVje3LNSl+gGFhEzI2BEumTUCWO
TC3S7qz7o2QF1nnH1Lz5gLRgYNsZz41rrEd/ciGT7aCX/ROigwMSbvvDBDu0MtPF9q5tDSA1Dp0m
0B2/7buDMAqP1NVgvpYn6ymg8c4IBviG2sQpjDLXgsGSw2O7JKQ10ugiSYvBSztx+NWgerHU9aj3
IJajiMCfKXiDllv28lSd08nlUM9XR1SYejj0nyZzkVVT2WzbL5WZcKT9nCTH8XCDUmlZjQqn95Ij
lJjzzLkdoenbZ/K9FqjcxpSuiuPznTTqLnxBjygwc9SgB4/SPFBlqrXZYo8nX44c5OMIvgP15ymQ
tZl6AbcDwvbp3pfGUfCyS2h61EZQYmhvq81nuxlmIRsiWio4C2rm2/TKJI9sqgj7fJ+RgXg03r+T
TySOtqyY7VQpMH3jZj5fE304KlxMbqtlWb0cB5EYVihkdAT1t6HH/XNkS8gkq9tDBCagqxmdGfKR
trp3uWgYy8CQsvkimZ1z1PMRWZx5XY0ya3ZmS6kq1dkzmahA9gp3LdbctLDQX1todMTRpAqRMWwe
mayR2J6/tVHShV0UadGPYnUKkEE+DMn4Z7yYBiBFqOOEG4B0Dml1VuHKKk9aVT2wpGSpV8Q9qNyZ
6w8D5pWYo2FCBe6Ruzdn6B24vjD/rWYyVDzGYrIWkCONGgJjm6Q0myjzcJK2+Mvj58jT/6drNzq9
p6PqqbMQXX51gO++RYZ7S8+qmJnMsRjkUKbcxoDBbnMIxkcK5lPVTeXXHX5LzJ0hBeixY7QauA1Y
PmTwVJIbLqFUoABg48XtM3FgYDj/QExqmYuzoyqM/mnT+qYPeSDni1X2NvjP3kCm/kOGjmBjcGXf
DgrJgL5f2fsPErBdUY5inKlhtjNk2K5+PklhELKT/D3MkJ2fVi/2fXaSrFqwZ7z4TGFr+H8cTeFC
gOJP1qc+c1P2pv5wv+aAYdZOTvCqiyGCoS0WXob+mExkh8MGoNVA2S7OdxT2HDv6yf6TsBzvIGcx
QU+BmhL95tKc75Vqp/NNz15APbSUsILePbVZvc4NmDkDJAA6P/TQGKX+ThQB5YtM+Pan2CgrnN1j
w3MB0QD/ntznZXx4YXJYVIvvkyc6vumP0/zjgIdTMI82dNaYB3PTFQJdtecLeDWw7mouNRoxH7iL
UL2QW6IvymBuv60T9kYTuxzcMzeen8Qf2sT00JS4dq2Xy7eiVZW7wBwx7kAXfsguekuntm1Jas3w
cTIBlk6br10i7dKwU+XDllM4jBy+0l96DG/6Dxt5DqiUa5P3ZO3qx6frXfu5qRQPhy8yRwcY6FI8
ZiBbdEcXsPQwIXUiXbHtEsDvn8pthqf1Oe9aEn7XN46YX3/wr/4MGqLsSFJ44s4SKQlKKmf5cOf8
iNtf5T2n5tz8hPErIcZwC/EKE/Rg2uXjde0hKdYa0lI405QxvFyfhfvOUfK12/OAVUClYLpIoK42
6UCNlTOKQvmQoUACeEto20dTQrwSZ4R2wVLhZD/Y/MaqLAsPOBtYl1bJCo9zUtXWbgSE6/JDWcSO
hSYLKg482tE3b4yEF1zWCvbrQkmahr7Fzw6Tz7tph0kFHb4iiDCM0NidBEiCXXTTymvWLJHjlvTy
RbS5mM4UvuoKBofht/XIu6qtJ5RDqVOYk1deDcFOMRx2lGeA9ocPMDX7I+sbe8Na5bnJhp77qAzC
FSNNIivDy513su07508LS0BYoTl6J7MjyRGB8VezUz8xezhXbx/zre88b0y2Z55WhX3fyh2BcCn4
F3JnCkl1wmJOwGhL5fi/UJ6cgWW8CuxU9GGE7e1kr7E8OidDJ5fPHyetm34kWZ1tW8IemvWMy+ug
mbyJG01x6VUR9lE4UJWHRkC2kESvo+Fep3L6wfeqY4hCk3iDlmemmyqga88sKc7iVMZQdl7pSPMV
AwI2cAzYX6YnM5WVVS926Mv7grLMQYUepmcbJHSl3Jb23EgglihMkBdz8ZjHTGNZR1m/y+V7+qtM
dnivnAZDpYSvL9HXGaDzJlFnTAeSHrg4ERbKfYYNmyDidMtyP1QJGP5GLXMz7OFyd/5oRxfT5aEW
AkNVsG/ERQs16+jt7kG+lS7LJIR/GmetVcx5cNYFOw/c6B4ohScFArhzGWvY7N5jt8cAYn23AwtB
Ds//3Lo7gfo2WfxgyaQ8lPRYrAHNe3CPYSmD7Pglc8KmxbAxsaXN5I5SESW9nSsWiTZH5i7pD107
C6mlldhpd6eimHo0ZyIzYktwok2xHUPGflQkPsYPUaS2nNcKK/4x8OCXCAF9TyI+5EUUHtlM0yud
9moULH0/6cG+u4mblgyGgy5pbnYxm0YVEHexbNvaJ3Jyw7nMSjFL1c8qhqd5DLTfVpGZbKdDGYvj
KqZIaQx/kNircrQpQTzqSbvfHOhREKNA8OaV0WtHlLVhveHlHJbOyU4YXorORTvAVcCBD9XexfQj
Z9Ga4owNoeMPWbiKq06On8QX4WpMFaLV7GIwbsd6dOUbwe8ZAJc8sftwUmkx0j/k+HoRVSKjAzPB
rg3zGiVYMpK5d/uZWO4SfkomzEwOOgzFbcDDduCZMOfvgdiO497jmd8n8iBfSPj7VboF7gE8YCb5
yqYidfXgYD+qRwqstk5GEj6JJDcAnzfEj4sPXd8IKMPVY3x4wpvB/tD78AruBMtmRJituEIbU2zj
vft0Iz0PC+4K5srW3aCQhFf2OpeE12eDRNRnr52wWvRrEAJmv18LAASJFY/FGAvCEJaFsHX3Vv+p
DzsflhZNgFP0kIuQNmzGRN2vUVPaN9Tkh29E/iOvfKraqflmWw/JPh4Sepk+U3+05ivC4fih3Xc4
L108ha4wV2sijb0T3oYrhuRox84tv9L16enTJsveiQOJemPxbnYbQmnpiG8BInU94DKj4lR9TKY3
Uf4QitmjkZKZAnVb3Ow5WFPiRyrQfvTEBr8RKQtTfyDZ7e6aWQZTNDzSjIrjGsfXzzPa9HkjqQY1
3EWZ3jkesJESLJjyW0xOMwaX1HFNWmD4D7d/K47xRZW0AIGI13kN79uWTHF26lhz1zNrG7S3Mqtl
whNTXqQ3MiQRh6wPWbdiffIBb+hNHY+rEFwrO1wl1nbprTUKrGbsaprib1UtXBctcN6x2K5s3CW/
Bu0x51xFMMiEwKCrwRhr8XKyHmuiQhIiPq0X0ZVt40jyKQMjd1U/q5U7sZkcXvdKGhNcuzeFMVUf
c1U8sBF+hNcBkhXvZQ7ROMVexvjOaRLOX4OGBPtM/711L4UuBIKVSx3FPqUSDhqckGrNBgNW/UGC
1mCCdl72HIOfuEdS3/y5G/dLk25ovrzzxZ7frhlKpKO6XQleGZr1JnkQm4C09sgxHLMG00R+0SND
sQJG5DIouVvdRC0Urhf6lHIDgikNRuiknfAlEFW9A+hYidbtJtuSxWFYl1R5t4tH91N7WhCoN6+b
mw5Wx4whYnxyGp0PEfGOcuERzTYxpNLvBFqPtcQ0/AmXi8BI38QnD7cTGr6lCuo34Sqpe5cLSjdJ
0rJgXhlmojzWxk4hvUrRKdH2YIyQ5YNos/xGx1Cf18OVjWT1jTzKz4MndgK5yroGVYO6/4CKmaWP
MnKnQwp37aaSkpooCecaHk2PMjK8yGl5x36BBhJ85V+j5RSqUIXhWM1HA0ovUCqAm1wjYb818bAf
CdlUM9zoKZF9ZN2LqpdYFilJnxfQFJIZIuoYXZUW1U8jc68MFKufia57Grg9zx0Ah7jyTgeF9ky8
iHrpWZvr2vfpDDikwqCstIZBsTMWzYlzn1quGfXxaN6OylZZtvPeri+zYim3pTZxj20Tyu0eC3G5
wIob1ySaY7wEpZiuLi3YGiY2KXXCcPTDqerfsr3hVJDmyZEcWqV/tBjl1ygXTGQbjvnT0g1yDAgf
Br1e3pfnOR/GfAy6sirjkn+lndYGVKKNwCT6Q7fJK0ciTq3kBCv616Rzc4TdNjSGhvIGZOv0XTs8
T++rz4BSu00KZKqgzyX/Oh78zIkdT+mJNmEApBtnBhCDhxta/B3OCk7nlbxc3nG7DhSBypDWS8a7
W946blAsUBCbq1OZr7ctOQiA/jV+U1tWjFcJWlX5Y/RziZ5ezpI5JSB4sNEZ7qe0NOLtHZqgdFjD
lTZYb+S+ZcPUifxI5OPbUBl0nvyro16c9sDkYcucB0zaJdjYABWJmttEApRVXepdC2oHFmf1O0pS
PJTsP4saYog/Q0YOjg6gLLyz2kI23FH/KsIUa7sLCJRGueOQH76e0HpjanJQODfRjvfUdfF2iSEB
De8KzGzqSBVM1n4eSGksYSsEU/U7WLsM8+lDgm+9Tbb2zEjxsM/9doOPweWndrcU/RSHw49JFGVC
/Q98xcUyNvRcIme0F6Tyzv6y7TxY+A0HGAJKnCjEa/otKnnJ5Kn0FdXcH5AYPzW8LkE7/aIdmkk/
pO43PFWjBp7qVbAnqY7PlogT97HTkHFc/iOe03O6WL73gEWF2d6eqmqvfPLZiiqiDtF0jrad+G0S
+ghhGioOx9Q7Vsbm0x2mxQ6x2bC846DeFE6OaqFds5LanstCVRSC4QsSb7qPpB9HrKcsHp9pTQr9
kcNoGzfgZvZO2u7jWroU7IxQvMupHDG8uAvxynD0BTE8vy+1AYfviEp21YGaCG3Und8V6nLtVZxM
dE2rtmToHXoTUAzV4SHep66Z64Cs2d3qf85EVvVfsynDybgyty6GyxQHbEjCOPXVcPAO8WDGee26
tuFwE7DMF+DOuEtrRbM6MpGa1agYnFM0aVobyxNEYWiSg46I1Zz5Qw+7FuVVO2Dtg2cRv+fM5Ueb
e24aVKerwnhVQVQvQhvbIo45QTA8KlSmdmYFxNCIL0UH5n2qyFgRq2ayRLjlPJU/wLCDXpUzsRf6
F9g+rUjD3n3soCJdRukopDfKhUWLt+bRRysbiOH7+X0a+WPWTMTaOeJv7vZIEB8esvZjRcsZO4rd
X74mrepb2kqj5WJkMM8OOVJCf9wAD6Q/UyrPCW6tpz+7YiHicdV7V0EouZbX3dybUZl5IHjN2oAz
fZmtc85jP45azxMlwIuuRy/wL29+H/Anb7XJaK6/8BgJ0yPt4/obKlf3THqK3hQkS4DiNu9VLziw
KaM6DNGtsbNrQ4FpdNSLwq+TDxc4DpHG9Y23C8vJ+iI843O+fWrZ/gCaHEtYvEhDBxaJNf9oB3Mu
RWCGnpfXSNsICVKvwYe9/AS892zzwC4nejQMOpkcNkhiINXdZkNUB79OfSm820uciGVkj264mSNe
14IUGnjCqStIBcaOZt1LhPjdRa8KN84gUFm3Fjd5YO6roNjGLvszBw7AFwhG0EoqEEFVErdq9Xvl
3EAKHjrG6dLpqrOn9B5+bNpflOUMHVa7KAkb2Q380guMAL5DIXdk3dvPEhoPtmfzF+wRqw9s1fvZ
TS0rjKKVMCIu+B4wUvRIsLwfgdsi7aT3ojqs1cIgTOiMie8QQWfGoAqomuO/AdOnD5H9mCHSnncA
I2OcP7eLFgQWtn9gTW81s9gE1tL+inlU+IONkKllxIk29kj0q/VQ3scWJhJs2Tskln4UKEKMiZw7
vnfvo8CPrW9viXwYteayqF2RnregUu48iCsDPPcyv6b7vIJM8XhfTNgN42VVnW7l2UpbzDzEVBmt
dYhK/v6CYrqZCTWzmZmaiHwp4ANA6wT+v6k5GiQ4fKqVKItk4k2Yn36f04LEBsR76Fz2hw0kD7fl
C7rxIU8ExfxSJwMBHU5iPm7K6H/xz10lpyBt4Dt8cgkpJpycLmP0wSodlFJQW+yny2B1QyebYmmd
StVt4vq573Z+TryVKtny7/wuH5A3UTLZnKSEsjJDUUyzitHIummZ84wcuEE0cUED9BvsF1XaeUjF
UY86Gp0FtT3PL5pznLWcftr/7XnxRj76XOc9b6qGmdtc9I+s/q1UkxyVitTf1ve64dc1WrbK13pj
F3mIwzkcdmSXrxUzg/9p7khz/6w3Gsru6BqkfKcbKhOwo951CHLSdX26Zp4oHsS3wUGJigYKTNT+
+tY816206t/0B4ft3vcSptGjqpu5cDsKl4uumRRCgZNAQ6YTAfOsLGSnxoFPOX2ckVFJp9VPZwri
sOMlOGH6RdHAgG4Qz1BGXbm78JT5Hj7HKbXM5cZ3dn2c7e80Tuf3//kjek5VfLyKhb30NBpKluTF
Qf2PbZHVUHl6MdaZv2Kq2MRxu0s73gNGi7Dp6j8Gpn8tbsjbio0lnty/rmM1fxhk8mXPjBg5s39+
UoPtCo8CTgw8Fn6gj3QAHnbvhEjXlm4ms7AFyWYPg8S/v6/0nSzUbSTCaVAjzCWKv3WQhpZYPRm+
hWaWr3II3ECA0Vm5ZAbSpLp99OELlOR3s0nezEq6LLVwrHp30XbmEDXz8oT1QSBnRTdR/jArJAt6
JGyUGa62tkPCXQe+up8ZLMXVJoztl53aygL04vdGQu0of6jZ32yBV+l2efvOdUozhGPZ1pdNaQ8X
TjDK1gyp83tTAGjouxu++ivLsG9WB6ITrmnMOAzq1IWTGu37n+SnQ/LSwkj+aXDXR4Hyt2TL1kdo
TaZEFuVt3dYoR64jywuMY63qVFCCfCy9QG8k/MK/qe3nHO9PvjnNBR04D7WSlS+tgHyMQGUjG/ST
fdoiQJ4DYluv/1vbCAA/Lsi4Sq/k3Lx8mhBJb9mJw+KgbspqJb82Xh54spec10uym1yUtgWN1BP2
zsIO6AXbafeSh8J8ilU6lUJW+n9w4OHWyHl52IjVFgatsDiXJulU/MCB1+PjZHdq6PpTCj7zchc9
+2voq05vhNtafdoNWpc2aubrlaY7iR5yIhpfs3sYrffZY67W9Js8ld53UDdcU0R/yLuvGPU9IVcx
JNcZP71Wbyt7D9JPy3AHkQxg1ISRZFI2u+n39ngCzLNhq3zSi5o220d526rwruslYDeVmcIHg8Fp
bGweL/tai5fBIu+dfkVvA6ArMT/54SjDBBfrKdQmllLZxM7KTDIWLYy5EM+ublGddBqjq9pYrSa1
1IF8uBUbaKG0gx93hcCC5vGGRYJ+lOhFDu70FH1ok3UUxhQjR7gU8SWRHNY6gZ2VwQMkKaLqXxVq
RUuTNFZrpo7rUGojrLkr7MUlRp/hiWGqMxDPmrO31hQXmTq6NHsy6gSPDzymh/kDae7lht2G5BXe
PMcW/AUVqc4TzR71c7CMLgJY7CtSc+mH2dn0oLRT8oZCazRsTEhLKjIciDQ2nBEb9hHtqniafS2x
kZm6vqzhpxmUR4PtxTt944yhEPhS6zPGGJG8fJGDiRfNxE8k1u1//N/oAqHzSNWvcR/QrEKsQhZ0
S9yXwB4nAavnTz+nfTDdTuGKqKGsv5NgUSVXohNMkPXGPQq/oqKD7K5OyVEDTrjKMmiidLFIiCy1
flRbza08fkNF4Wn3jDLHK0rhNZGCvwbefn13PqO2kgyn0lxZ6JM9y/GVh4bredNYzaZVG9ACRrTO
T5RgaSpwm4+XnFnwd77tVWLnabBAIu8RdB7bp7PzJP+Y/+7BdIP8KUFv0+9aS75mEFVm93fC61aU
m3eTB7begG1U+zxaDkzBqCCz6Ge2w5Ojnk8H3/biazjcfMdBaqiP0vLu+BmGgii7KPjAV9CYC+Q5
zjZvESbTvZp5YqKeosVYIhKKqtdR9fIBem6mej3Qs/N+EjnTPVStFQgRK9vQIYdiwwakjJi2MkIw
gXXIubP7S5jsCv/EBUmVUJ8KV3IAteD0ErcSCjYzg6XSdjrDpr8bhNmECWW6EjL9Cx7jGpi6gokH
d6vfKmyL3nVx0uGWFyb3cLxz6J1Aor1yMmjewh6/QQZ/4KjDLTgDaTaGIsCRC0eLnEEYRNkZsdoe
WK7PX0IZqNBlmhtmaJu1d+EHGYbFCNognIf1taI9x2wUkqsGjDxhN9bEWCIa2cAUQ5tQGaVPPFOR
JmEynXgqsOdOWMIpJHa0AVZLJl11WEklFUwGM7i9GF4lynhMriSmwkcsLVSlwq6F/FAfxJ6cDbqI
corvbSQo9e3mtpMvNPWZ35T6TyUmc3HgXv1pZCka7fxF/GU3/tQNnRGobIZ6X7kMHekO0Ehap4ep
69T7cSIkdpolHeM49DPCkLIiN65CB8Xvk6k1rCiHib4p5Jl/qMiPIHF9uFZW+a28wspecXM1CFcb
RIIdGPeSuWlEiNsewacYfSDet90ceDUDdOKX5Pm6p7nCbtOecpfGeSxPGNukInprbAxebxCJ+aEC
mNEciONeu/wUqJYli44fcaaBm+B2R08Nf1uxzY/kmnvGTvqX4HAxwLOlD3iFsN8cCXU6Ug3hVvA4
QcPQTcW7aWA6NIr9CtsX8Eu4SC054nHykRb3HB7KkMO8A4pDqR/5WvmtNaWumPZDl3H2RPWIriQ4
lIXoOFAeUvWZ71ZIfAD7qb3xQrZGVTpoUG17BOwLJ147Q1FyRCsGoYQDZxZ8sWK/tA9cXA6R/ys/
zxdnMLS0tiqtjgul4Aj37V6NDG5jl+ZMmqsjplVqabmWYeNkpPPHi27x6p/IPN2GyXvHTHSwM6w0
AWYFn22C6yhzF2gGHltw3ObSwcVU1kYULRAtxnQUHSY2GPFK0VQuwf/Wt1QDBAGTelA54Sb+U4K+
fSuQoLh4OY6qok2PSaAL9jcKbiHmxjOdKB8ELKcVYauddJ80xg2FOCB2m96idIRQvjqTKp67U4uC
dlJ2r0kz8B1//tjk1avJF4WIykxMBxNQlRCzKMYKTRtBY9r0D3ZZHnu96HC072ODLMqdFcUnQ2K5
XqW1w2/ddH2zNhjCpZ+ib/cTL4V9FjRtYmeTGvHY6yCoOKGHFMEGtoH0H+4qVZ+gfCkADhCJKUWl
PUNsfcyvrXwYGUTT77IlfilBYqvd6jq49I5uqC7CgTZxJ97cfgr0HtruN73f21EUbGg1SskdTN15
q0owD3j/B5BulW6tYFoh9d+JbBodwwje6fKxeAP7F+Prs2mIYOkx+YeaZ3zKXZBFeJc+mkee+uDc
ONbtAcR3xbGhjvVlyXvAxTOd5MnF6eDsb/Agpo/4M/FHVayJEjmPrRdI89t4ofL/waZn3hibio1d
yFPEd3Dx0hLwAuhEQ497iaq0sUig4uODpZP2CBU83VK8af/HTFaygXR7uBSkmPyDTsxLXlCdq5UL
46mlrOg37T6j8mV7nei2rE7XBXVxLSSWYaJS4I5VV/hQbvYVJD7GxGOclFQgYkY6u7oTyuLHX8hO
+6Kv5qPpxtPV9g3K/BcpXP0UAZ/cG48STm6AUE3S4FEXfiKGTgPyd6sDQ9CwBM1Na7IupRzFeg6X
G4hyP4p228wbz+zUWxw5vohjyjZlEkNUZ/8LEkluPUgoLxSPkQf+wQM4Hvq6UHHo4Qr76CiihWBz
nEAChXgt+q79QYfw4O3pJ372nZWHU+8qeEf2ivDmrjAObWElkPqZBMExE48wLc211VkboPCDAPHg
qtkkui6bQ7U4cyJpIwqKTk5grteWi6krBKocxCntju2ocNpPiaXzHs7w+mvLvK92FiEYMmBFyp0z
vtMc46NvV+/gIYW3twBciARgAew1cQrZ0sfH7aHfvsF3rQ+aPgpqrOeuty4m93nXbkv06x0F2aKN
gFz8Lwo1dDFQeBR7Aqzs0x3JYiBTSHjijp/hhG+ekGyhrXnWKfWRdk7BmvWakNYOGKBiUQJpA9If
tZwLAmd3Cy8B8nWVCz7rXrB6wTLeROxMmAWN7MbWit/a06rB3ZSiI8CWSjJgIgZ5qwG0dSOBlsgp
FOFhSYzIIdpoIxrE53wjvB/XC0RKHk0fFPpjryUCLp3nUc50/zJkpv09lCAPSoYOPZlmpXRmbY8D
VeJdkiP5BOZrkoUrgvnm/GTjja3W3CBa7uwrA4KtaGQvAd0z5wfaVsHuL/0ApiniasoXyYwZUCjC
nDGw+i1mE7zRkl81LkhN+nZ+eaaoH+6bsp6c57Bj9dh7hbKw509Nq7AIje5ynQ0dNPLHbbgpXSfW
EW7LOdz6wzDYvNGyNyivU3nUEUhy3ebirkroZ1D6CLzxT3UzKmOrGG9RCYfhbymgBiFMuly7x8dk
eNSnK1FlCkUunFhmzf2+QGTfssDZbgDOPymEs3Sch9tdhz7Ml7hIDgq9GELuvQrdK7z+Amm3MU8d
XX7jwdQjunlq8rFqZyVRLcAvLODqtHlEIONtSQTAMnJNjykwtKGMx7oaByLBUHh+KTNeNaot5Qxn
1QsiODn7er/PfIv+ifOAF1QLH8IwQzssyL6jU91B7+3K5FL/tyQ85AH/5EqrCpeR+v57S/Vf6lnk
VR9+vIXXhsQErBhNy1ImX6P4EChNvMwMIMVJwDbV3zkgwuGJMSAdao0A/5IT5rPlnCNsmD5XxL66
+yW1qVRGPJQPPLECap891Vea8/Ig7bvpZETfglSmhtw2sq1Pas7m/sroOhXlpqFyf7per4Ml+Xj1
H/FMEbal1OTijD2Nzs9OsQPrf3Dcdg0PKUk9Ro1F9iunhLGmL8iFcg9HP0qiUEswXwnOu9dhuq3/
YwZrGUTT+9KhiDcpeYj4a0mAA4ybT8krtWZhxT/Ga1aikJQXoNI1qWGp1cg75WTYrbzkinL3hDA+
9gFwLox7YSkZcmecymiymHVm52hOVji0eST4hPnEXhcnPFWI+yEzBNluSCj2Np4yQ9Nb+C3eGghB
OeGEOp865Pw7aysajleYlGEZ8tjmyTTnsLRnwYclYcfnGqv/PNHVdy3VELna82nV+plFaZnnx3SS
iqCmMIjmOde78WyDaU3A1ZsuB5Xcy6USNXlAiZ/FT+IvcAac1bQFwO63yaFLggp+y6x8AYdTVS04
IpgsHBEiwW1lNqQ0315quDfpTFqFHjQ3nrNZOUC8gF5Z+WfEze95sj1nJGKcU0k45FD4qnTF3pli
/Wh3NYdS0ILe3LdbNQewHeP4ewOOBPeWNqr43g8NVtl78nv9EyDkg3fkrs7khnL3WmJXyxy/yqZy
naAXciO9hmIFRih+RWvYSo1fUMX4QVoKzf3Tq7B+TTHDnaIYRVSFlx6oCl4/Xa3NqC7tGZAnJe5z
b8xPXucUr7tJ2QcPBeAdgOhWI8plzGsq+1x/onBhaiqXjqeWmrORxudy/Q1zoiO6BpLAtLA+FkH/
G1KdiyXRkfhRHAtOcL3ELubHGjykbR5xEkudgDOmwGJSRmraJ1dyDzBN6qHue+wYlBqXo19VYKCO
hQ3S/A+Tkgg6amfKPeP0ogyujsGWYvOuZrONVfONq6HRMZ+7EFEWfLELFbfwm4WsiakcwH6mLnmq
znWuySoL1UGkBhfj8GSANAITqXtxn2nrlyAmhxYXDApLCAoNj8igZvg0GPl3LNafYRFRWNODlf8W
8Y1uQ9ayk5YE0wAsHwW/sXdoNBEXLV4wKRUxuxLdgmq1yFC3sKP6eaaHxQrgUILz+0TLhwDsdWRQ
NjBs/y0G4JpI8wsIKiasBFt1Sw68f+HVI2DR+YHBJzb6CLeDCVVttrSYYsaC1Z02JjdQ1tN2YtpO
AC085uod1wQELX9tub3yUeObVGJ0mCm0fn21KQiF03ZGwMPzZIX20hGkq8CJIoBvQKCIubIorM3c
9ORy0kRvJf/Acli5uExmP8aF6C836TkbxdxQQw1hDREZ2qFJhzqHv33ow3wCjv+9PDJw6syqrIgi
vQ5gN05J5f4iaH661bVqs2LS4S7N+Ncg1v47UudjqhQgf8ygfD+7Bnb8Cl6HqxQeJMapcxl+bu7S
RYhuxOUbRrAr1j3mgBxYOzC1tO7oWvL2KJOJKAF9isMrFMKW6bq08dTgl65qN27ra90K5dSBMIH9
wAv2VZsTD3Lz5a6u5twth0XlIwKrssm7GywtZbaN3wKwp2CttXNGd+DszDYNc1aHmIbrMHJNeZR3
ifuItdj3MUKVXMvLWm8/sXGSdFQwAd0tgdtPyEOh3asw3JepxEh5GE1bIw+qfRmhJ8aLl0HeIXUG
hukceL1gaVM0Mpo3cLgd+DRBzzzpvebZ6JZrrUl6xNkFIydWQdzM5TGleznZRbIl2E5RC5iwa8lV
z5jyFPyzmw/sLDUHrooDvCwkj2C7PBY2NB1oVv72bMd92hG6HIX8AgNYJCczirltmHemHoXH9LyS
S9q7dm6KthCO24KJrMzqm2EO+1ESQ3kWfsB/uFszB1NuEmvLX8fgTpxXzJwXynrstX+WN7HmL2oI
v8WygZtNJsWod9A6zyNWlmt2ZrZHNOPhMFQRZYXsXnuxQsdBz9WEq0tFWgBLUWxoGPYJWOXKFLcK
8gsaaqhogW9TVKpGIukyUTDnlvnvTIimTUVv+cvMdezSncrZNxKCm8GGqO/sWzrh1WBpGoumehd0
JNWMNcP5F4/04XmHWoivlsezmdXe4o6nThbgsnpBrgNdJVt3KkorVP9Oli31vdoJUPe9bEOwwAQn
WiKBdGGT3VUl8T5srVU3p8yXvNCozds9gtVRNGq8LNojZkV7USl1DxL8nu9O4zsTE//+h/OvA7FY
2jrFQTxPlrVvxKtYz5NSONKniGBHEEC9d3WlNy1bUBV6FHVgqgcrz+820TM6U4/qt1xQCfj0pHCB
JowS+y7SP4ZWZbT91evC/WVKg3As8y9rEgP6wGeweGvx/M1tw88CRC0qLkeodI5yyEKzSSFjCQgP
lMtqNXJxQ0NGy5L2ziTpNljlAerkTBySEupwZS16PKINmr6NQjjpl1ZJcddMgqrM6RoOa+0B2ffH
4pshKuKFpWWOArTY46D/AVUBuJ31Vx4oONXfzYJN1JJABVN8B+85+m5VDPjOS6fkz9f0cJVvCPlE
kGx38mSMskX7kE9Pu1OBLGiE5zwCTR3Nrx+OXV7SXfoXd6Pi3+cg9cC2uznTk3KXOzPocpcB5BOB
bcAgnASOhgWoPOQIsQivk8FgS7rKB7QGoSCo7PeyTRlV3ZicrT8kGO5t3hAZpv+lnSq4i8yck85l
v+BFkM1a4r0AflHvdIW81zZzObv/ijVD8ekZhocPq85hDVNeNc7jf8GoqkT56TMjStW1SNcEEG6n
/8RYuBdZPcUNVVqAHNwpzxHWS1OJd7H89bSsgpzYH0PolCNsWnUMpsGJ8vKAXZjG7PTkp334k4II
fVhuCmS40TSxCuHHPsj/PFlwiBhOdRv2sPsjr5L5FX0r3fouG9Bzp5YNFlFXMXiB8suhA/AZho32
E2MDCPODJqk8Ue9xfPmg0CAmGrMJtwfQOmZagL/a2YdQUk1Qzzp1bQx0Hvzt98/juhMQtOIwitz7
b8RMCv0xmFCjWe5yJ26QRWDGprQcbrJNXuFlrhvBT1eBpsR09U6+J7diT8q1tm/Bul1rSUx1X6uL
DF9owVjag81pKhNWrqRTK46wWPGyz38MHWlwikBpVvcqLeTuoz2iHsJPOMTpY/7/v6RO69O8mtke
BwhPcgleML1OBNwGCtNjwapI9nXEzr7qXdcToJvyesQSI3Z6N540JSGlCqWz6HKc84eRxarw9Qj9
HOZrx9i2rzVpWitl4B1H7awmE6Ytp9Zhs90BAf6ylHUxwJhqMp6uRLP3+JIqrvFNwQDX6qASWKd9
8XL5L8kpVHE6oYxUJMeHWJ/kIDcxEhBDAg6vj35R/75cDLZjAJ+GC9YmaDQ53WDOhqPJQFOerGwB
heXEOyHp7gzqay78lot3BlkZ1SuIJcxSWtk+OcCQyYCfDecc0GgfBHZrfyf2xmAfpyzCFgjkY9k9
U+985ubWfj9k8P/NyZ7wNhaYxbIV3EdTlfBpo36O2Zz4YLD2VfmJzVHYnRv2Xd7I2Md0XoHYkOhF
JYHUvl7g7b52ft9xljcPNDTDL3KauuqS2Fx1JSObMHY5T8s8HZ+eEoMlkAt19kRqIVyNcFhS8ftw
Un83+i+g7vfdEdWACqWbmEKTalBPwCHJLMfOcqBa3t8G/tHbkg2uVhRMItmV1mCkPbK/mbex1yP4
aDZnYf1e0GiTTXgTNZFO4wdhwrSYWYqlovJ8Z8OFN3hL+gY5/Nr8Li2OfWl3vT1vuM113i9K+IJF
2AHGvXoJUWeHCpQx/6X8C2+hPvxgoEB/JWhVbAHTwwlKVBrjRKO6j4CF6Aj2CN0RwHLeqvHDEbqf
jtoG/Z1u0SQ7bxC34ZWQkjBDR1WjepXH4axf13ZlYfAjwQs1nNKPsaPiXQIbBmizt/h6nrj3FWFk
QxM1mbrlIrVEYSwEvjBTOel/bR84wLuHlDkmF9+2sxX0v9HWcV5g+uaSjjHTW4a1goxp7Ft79jyv
SRKwSpM3a963BE1ls/ELgVgLkAXXUBV+ed9E3WtZSocE8P7a/2YwmFY4RlfE/VzWRPwSYN0r8ib8
EMGGJ66XXJWpuv/Ao0a4TNOUfu/7OLhP4fKsx7TVJyLRU3iZGSDabPR1lWmCFkCL99HMSPezv9t5
ha9+1xF6eH+dyHbw8HGJzAj/wXeRnsIUyliWX8rAIOxgXiqp71htXys+kxu14dG750G9uRdl8Ab/
WbrXnhd4eoGs8YhbqCuGWdkNcn0xsw6JFIimFsrhVjgbneNZStGV2b3DVKdUKBbgOLek2mWvHhvH
J33rLoHX9xSVw2ARaG0OAL9c/6KD8d4hr68SD9dbpJxRC1QuIsDX6WgMgctxts6FpvMQpE1LvywI
DsSEEtlVSyk5/pQysLdhqKZBKvJdK/G6lgwQ1lOSnXY/anOLhB83iEp/HM8KNERLkKjTj5QLJxA0
Iisef/NvoYn1fsm4Ds9IsldFsOTKW0Uh61tGixB5rlogwpsL1EsjWUGG4+blq/xl13UdyKx5J73O
jGITkKNa19Yp+SeG3AMSHeO92qp58nQUwt0cMKXxb4JSU207iiIgEc/TQWDvBGqhgpoAZhSgQfR9
//hdSwSYEtWrS0R1kRz2K2qH0u3l1R8k94glDMYfa2Xb10xH0nB7BeGIY5gIRXt9lDCKDeEIAC93
AX0vdSVrxeYoHB+xgxRI0MZww9BmDjWz1dPk2ASt+6+F8SVd9IsOQkGNENTXUl3ejizx0G/APdmN
/uCA/pKo4f4bjrtJVZkLdudhKv9uH7pbBQfi7oqMIlqgfVBXl6WGghYP90iLf+WSqHaomE5GHSLh
GQ1iV8f+uB9pw9xQ/YwA3MpdksfsKCQyTMWB/jgw1CRQm2oduzH15H3iq8bPNavB7ZqP4s2kf7Me
wXFZzyuCYgvXZjUw6P7DdhXOvA+0sxsbAVG2jlRvHwFuqpis6aErRDZ/MmcIqgmS0ob7SAIBVDHw
mKBeY7Fu9I+UbSrkEV2ToixBuCBkp4QUqPdNEv/XKlnp+4xTQw537JcRKEE7VdUaJOJB2gRtHauW
JM3m0xu8VfglBrRpK4YE4cNnaPRpDbYjY9inilBUN6ZAuyxulXAu7laaqDSPDCK9dcpGQp2UmK8m
RaiT0M3R62tAwugf4SkoLcJLKrc6FTBHy3bkg+Mqqv6Yf8IZY9Gb+Qg0blplrxAHgDojOODcN3Js
dQjvvLdpzqeygzCiJm6oNLb3Z6moOdBc34ak0zLEre4ErpAx5LKCKUi/cTb9YdgcDBcu0YPC5M0x
wc7+yDATVvM/jtrQsNbJNLkvZAX++qNn06UIV3yNuoGOlw9FRa7u0AGhBMICNbV9vQ3eZD5WFn19
u77mq7GZLY97kmWjD+uCOp0O9RshYCDi9RIx0SrRw9Lgmit4tSQhpXgzk49LP5Eg7fi+wD6UiX1H
xhxxif8qyRnRrowndb11itv8MojrkDS6aiMEvGZ/0Z7rqakbPmb+SBRrwTxKvVyc0ewtnPaEnaTL
2h6iwuGYRl+GdMD7v+AwOqvGR0d2JK86YIp5o1MiUOotpFf0u0/ddEz61XyHO8CoQNoglaHmGKzN
qkUr0wOz9vMGH9dBh4Aj7xrdZgRMN3txhp9M4D3ldCRaAilS2NeuuhF++tETa1r9dvyiYzTTpONe
UuxT3svL9xFcMH8NahC1pxe0L4zp1UvR9SYuS5uQoa44QmgbS1fQKUwiNsc9cp9KB//RUWPFD9xR
tUmMhQNNF+brkiCuMYjaEsZR/xJ5Bi8r54HWCE3slhp/Ha5OCm7r362v86xs3OQKhw+p7Qpic0yH
R7A21IyLmWqw5mozkLb79AHx8efijGUSldV52/w0dFBQupbZ3XAjfwGpFI3HHExqRymOx3vP5a4z
bOKI/miW5otl7/euVlRCzco+FKeV3TRKJ3vjrq2ZCo4mPiAjQvetqS4exDqa8E2fH7H79EV/32Nn
6l+Z29LjD0jNn61VxzlH4s9ehRN0Mujd4J7sJwDdvYZq8oeklGlw1uAcQ18AvC1Q8SUuBIf71+MO
GGyAnRJrYp2ovCMHnuVVLplSxcXAHLg66aj3lLJit0OKD/Kc+TPCmfQ+t4fgfTOuAIUFp39VXu3T
9CgzoTCkgJKkjm4UbotzljTgwoWqX1HmEmf1kBWVEqpKp5G98iKcPGu/Ui+koZpmsFZE380ua0dN
07OPbsr6GS5RGLweUDS0TJ60Zelppx7ch8oj2TKB1DrXG3/4w73+x6WG621POWbX+WAtjldwzriC
lXCo32zlL3j8EZ7K80b53S2njV4/Uhsr6OnivXt1enYwxHVJy6EXno7H8fOXGZViMAO19FnX8Nol
8hScHdW+XdltgEs7/N+JBfczcvwtO8MsrgrINOE7/PxoJbcAgmDpF8hSIR2GjONCM5pHrgNjd6Nx
vGflrk3JoEIEuC9/zQVyilkUHcnwOK8NVsHiNPaWkj8xNreef6Pt/046AjNbk74aL8KX75QSoZqW
3iM177QKu1mv7vDTx3qpZ3S6wAZy/T9oKJLGtUtURzUVUJhcNBCQiEya31MBSRcnmNhQ/Oi4ocjt
J1MrAtCmcWP+olVlgbND8pQf7Xn09CL91Hi/HKQdPzwowEXJEAm4rF3zOXsZ/oKp0aO1scLWyNrh
q6ZbJaFNsB/kSGf82LOKVmbuuQa1oun3fJvqye+hAl7B6dxg/mWwB6S3CyY1pKiF1MN43kY1oheD
I0eeOwvS04b+MUOPFKdh4HwmS0W2DNYwVr12TjUpYqOmcpkdD6RGJbF/NB7hp5Uz5FW1+opXrLWy
YXFF44xvVUEolv1IQ9qCVxPCZob+fuGklADGPhOTdsOX/kVGpfowY397aI0sTKB4j3dwvfRwqhwe
WKRELArzZlKWoV8nXpShessyDqNn+Ch5ZKKHy5wdCazbp6UT+MpyCje04bkddqH1BFHFbGNJU/Qg
z5y+dzxNVol6lSqZLeA5u5NLHABdKVDoN4I3+kgYND8goyXjLhkmsdslPkzvAtQ4XTdJyEkcYZqh
2bE2sR9y9qGdbwtDXi66k/atoyVe/1vQnot5xx1AepPKW/8jDfU+nqeqkRSjoSQpMqtU5HAga38R
I1aAQ+dTcfafdloR9Sn/oN6l+dHlSgrEaCrMq4Afpye9AYVsCO4ZrmHZ19FkzWHGyvLiBpMrlTCo
/+dqbCawhLFhSo+2LZe6PnZ5Z8jB9O9uShzp2cq6+kngZWJXG0hEqzfm0QWzBtlb/5Rr498OtbYF
57j1UB97tu7JEIxfuktOd5qDIc2caXT0sgjARB32Av76arQiiEhdux8msfVHOpqF7IR3WynPU94k
imivLxVRUnlU5lIPSQ8yVPRE5ECtrFyv8SF/Ky0KQ7f0ofXplio4TAOYwd/MhXwyUWmyLf6EcjdT
RTkLEf3AumCyIoaKAWgBDIWrGa7e9rOGY3f767LbKTbGgMKv8AB4XrnZNSQJv7lXEf5ppvnpmd1A
1tLTke9oYaBuXHOE6LcqyVuoSR/NG4vq5Xk73N5TGvuOiuC9VCtiWGCEYHz9UD1N4RVjpKCm5cbU
7C3Z+RSc+hScOvEOGPNkl9X0oaI7u0LkL588++dpY+EMRirFNW+RRJZ5x0ftM8Q2sKP8Iw5P7nGT
VVlvQUZn13kbio47Ct/Eo2F+BUsVg9G5aDfzq9aF1tyE9ATVKXVQ303aXWII6KrxINPdWUT5FeVE
4W1eR5QN7HplRjIIO+rQGEK2LU2et9VaEGMfP3Ofe1F5b8CLvDRJnDltGHkt0ibcubhtJ4jWi77B
3UyF5x23Fiovcz6rhY2MvQtDX4mlrRJ2zRvUBwSl52xjikN7Fc+U1UdlZC/JXSD61N94sTbH8DI+
fMCkVdJewQoPQpKcHHt9rlyOwH2dUPJmHt4Zr2mMwezm8r35VAtbda9SEABJTY6KgANow5OHadW0
cq+A5RL+bwi6lbRzmCgi/No2k1aZ7Y1oe/6Go9uOTEApLcJcxUYvkeAajjNJa3QcqykHmY01fvsX
OlVpgD92APi3KYdsXhfF/m5X2Yz677vQwc+LQ6U+pTOfOk7CswkH4ozttx0xoGPyrQq0slmwTUPk
ybILI/GRrDxAjy5Y3nX+CoYhcXkkK5l6nsOVIHXrv3WCsjfsGh/vfHARahFzUOSjMuJEwj3SQwl2
SG1d/jZkavko1qU+aLs13eFSGqCc/rjRhW5XOW64grzAoI80dp0yVw8D/uU83jNMtd9swAgOIR96
jHpAfMYhstHT6kzFx0FOhVt48gcZzwJyJp4crmPqIV4cT5fMymdFZf4bg/olmgHiVG6w7XZhgYrQ
dt09hbTBBIMnh65o4Z9iHGoE+YH7QNuFCrmwMEQHJhp9/RjsXLBUa90t3bOe2daEjIlODcbuCymC
SbZ9PiQCY4QNFTe22WHP/DWgIp401YLGAazODkryvg+UAPg8nzxrCSsTYJsyFbOAiMG8RdWcyDQ4
L3DTqERYJjWdsHazym0AdwBvuyNPhlWu2ah416xTciIU9NAUrJZZgGLfUcpraw7HW+kSEKxy+ew4
rNdt+6ZxFRxu/JBRBa6u7btsN8q2roXwQaWWKfFNG/fhRpQ2PDIvkgkjNiaraLrmQJchxsLjY3h/
WWZTArcPGFxdgJqyflUSp8AqiWCZN9poP+58+Bd6/C+v+zOS8BJcv9fihkFLjOp2MwAFYaKWN2gt
+s8OmpYqWGZeVvyB1/bMS2hZGBvQ5ree0HGJVy5UyP2g+HtM2oDTAw6ofM+H738BHfIDpyZRyJse
SWGNEGhdPtfTGTN8ShU4toGdp2nYseI3JKdJnmbGGnixAgxln/tTGTGrf/5SjaxaQ4l8eJU3NGs8
686H4AmJ8A0qXnfWwdNjSSD05hQJyf4Qi+Go6vQlOITpBhOz6BO5MeN+a7VAlqokFhzzSiWIdqX1
ibQQV0jxu1T7WPj42cU3ONt5lY0F2S8pQI+0Y8PGrEzuEzK7FhI8rsKmMd7bW4jqsuf408egENER
9AWbV+HmjTbfY7xHIwhpgZF81HCGiapw/GDbiMJjwQ1QTfL89etqoGn0GrauYt/nK5k9e3T1aEJN
Iz6FnmoeBarFwX8RAVwzPUQRssYsAxFDI1TZylyE/rEWchVy0sbD17Aysl8bgYSZbF9utMX9HkcN
JHwto9lzviTe4fAxtIGdpoKfWSQsA1JEgRX/vjSBH9IV+Dm9EtgBzCmqeyI523dHTnWPIXwK7ICd
7N5Uu30qXT/I/udFosqcuq51mKAYAlPYdxFj/hLcLxnVZa+WzLpoMHC15vxzjTTJpT6+tjfjC9SS
hoaPqONz/1g1Yq9vYLN1CuRNYVAWHjat6EjAvagIAIjHO3JBcuap45nB3ROsWmOMNHoKijpQIt24
DF9Fp5oLmUxE4iDM/3SSlmtSFNhWct/czXE+kCNK/37jjdiqI+eGA2/oj1lyWdjbn2H29HpvLmfg
iFiJmuJM7a/aWoYkHWDl+tYmcQNpxAHEFKZ1Avsk4/g+fKM6QuTZvAPIbGXiDwgDAaOHgdNIdF7i
ak2cA6UKVX9UGagh1FjLsQCVamQflQonVpy4Lq1kMSBOg7iGJdMfGwOxwcC9EyAe0U7ygQA0wRQk
IDUmuBZ7Z3qGe0joAqP2s9H1YQdQBM7Thp6x7j5MN8c01UXZNjaaQXdydS29SIrL7hGYHcremsRO
OqqxSdWpFhT8RDO/8rStelVF9PTPWBJ/d0FvSGTkOHZEQ3UQCS11l4aJY4fvVcd8vc9S0IemvJcy
eSvcRdTL684lcOr73vdFlVS1Vlz/ZO238Q1RBJsRQ8WS1VPL1ijAluc7N01hrHikm8PhMgk3GlSO
24oU1PImt9wpa1KD5e90Bz3dOwedbLeSYMgDm2HvvuU0Xoty1Qrk+Xn2MotLaygagFA+p56lTIRQ
MDJzXomVxtew8jY3EbMBEuXd1I13GitGeUERJsq9laQRC94cxlPK8vBrwfKnB49v3uez091Y9r5Z
IPVhciFu3yQmPYrHOR82pK8GcuLLINcMP8I6a4QuVIjMAThQ99g/bPsvabVdUAIBaRFk3Oq/CpkE
wL0v5VbQ6W3tN2BTVHrLQ56auad+8twmeitnJGZBOf9f2WJJdGRASObN/xeLawTO2WqPLrXWl//A
SrrxK9OR+SQNH74k9e6RLrCqQ9uwqPQvXMI4A3aKtaHeFkgF0FJoIihzf8ODAYyT1du0ILyc63+V
rBFXWs4Rdui6AbO+Xs8L6o+gdoM1USmQeqo6ddx6pUb9WIQseVG0XQ5CT0TJ5mejrVAhx+dTQ1Bq
YQiPs8qI4kuTgTVW62lkDn7aXqhqvh5C/LStyOOQxn+g5/1WOg7V3qwicvZMTlVTaN4QEZ1Q5wVA
oSez7h6U8HsfSmNzsahCC3bJo8eGtrnX8HidozstW1iefj/IbxcltipK/ZbNdSl+9XVie1/6WkGn
cWgYvExQK6gz9iDILiCXwNmZHRcUawsTOR+3XJcOkvJ3XPR4zWwmQHnjuc8upJ4LpwgGlq+rujuD
aaUqWMTBzQu/vjFtRBI5hixpnfeBcVxwfyDd2TWWdIQF2hFzz69ANF3QIWHEpXUKITnMYEl0vSLO
VUM2hr8/VY9HqogRd7VFa4/QApQQV2yvwYrZg4yQ8v9trEr+pGiBfdKpRIqwgWxZpfsB4KA2LHIm
A2zYRASDyeinySaJG2OIzI8KmVZWVi/JP09xDjo4OOZNNvsNJClu7anwCXe6pa5KpeiMC7Fh2VGz
HXDUN3jMj0Xhxm/Dc1i+nUBsRlVkHkNBDKnooIyyXEQUDzPEAVE0ihXY7mk5tqPWO3WSrMdonf1o
xGnbxlNkbMW0x7n4bjBEKXZB9Yk9eMhGOPxaSLkIkDT97rMD3s+Hdydqp7VLt613SjZINwcZ1OOS
ZIALxsceOIGLk3920cG4aRfPffzuTL/+kZaB8SAkw8ZhU26tOAGruNc7NnMse5BOW8yTUkqR9Q0x
BuUsK4apdETqrLNLFA/AKSVP0iIPUX6YKC/YJuzBn4tv+tXOsFtl4zdmpc/sgf3MvSzE7daYo0EU
/fF4/xslH9CiqGwkhYxrr8QEHupsvCGXbcnCB5UElPdA6UnwpqvFRX7OV6mXGM+OaJFfZ/g5pDK4
i5b359v7blTPJ05pF+4FsoHxej6aVBzfU90bHn51J2bCLKZ8xXrFpuqagAncocZlvClZceSY3PT/
lB0p1LGgcU1iLCgLZooXG4/bZZlvZKUQBV+FOpvU2Kfbu3BKCsyxkcf+ODVqVgtwYsBBXdOsqdNx
d20TWwZYJ1rgfrpKsXETc8LvSKH7cBdroelJzj31m49GpSCb2qZvDoK19s6p0p+r5ecZH93/aCyP
B92CuPS0mTV3hTZpOZ1DNHTpL8GDpoyAgKeAwo8c0B8DUaZZTCbEZXS0MQqclGrfB45I13jtmhSQ
GtZBwo7Vj122Q7Wn3lbCppoNtwaltJOMLz1y/TP6UFKL1HZLbrNw/wCSHsy01HFWdXpDn7xuKayM
RaKMVXuOJbw9ESSSXBJO1eS+qC32S7Dl35dYHJyMX7HKdnxQVcC4ke5+PEBunAN8R82BM3uC9rPj
U/OtC3sNkOAgnnBc6HIu55rw9wFgWkQVv849o4BCbKcqra3YuqKcamG5XKwd3s7SQ37GLJRkn9yn
amWV/gZ/fQPqnkzYr5KGlQxVfxZD1M/Tpgqf5/egitQ29yNdU04v5QC8/s4ENjsrbp65d5ojUsd9
fgaM9HYyJFV4V6olf5sinxojwRrDcPhVPC7ay30/SLIzoMQT27H3D0f4LUhih3nAsSWFGdg6JMpg
tFLPE0aWSFJS0pPhq+cB7PnUBGRgtPIK90hCcPcmU1y2za5aa/SbrfWpUpgfd3olNSbK/itzMCIh
Czf1ZNtK3D0DH3KBnLobUaqr5f/oHLCju5f1a1zD3XJ2wsh84FcnoMqKdxO8AHpBWH0YNMvIAJOZ
i2W0Bj7GxVZwvsBKLLHj5jeGdrrDJpFg4p/8kKybsJE+aoZplmjWjyBVdOqg+mcC/PN9w5sY9n0M
tvy2l7Q059I7aD2/yRERbHcknHYRZYU9qnJoywBU1FR5jPP4Ze/TUaHq3zinO4uyEiBnO/cnKNlz
DFjmbykSLbK645oRA3FRIS00blg5Zg4u+mUg+yOZi8yAO87Lon7VB1gc7XctgDUOTcNezP/MdxWg
lwfBkejGUkSQrqBv8zIOyQhBO0eV22xcA1woYYjQB4CmG3vduZPtGkh5kmnYHWu87zwtLbz6B8BD
ut0BWvtYAO9P1928ApC8GJcdbO3jThYmKbcNNd5QYp+gL3i6Px5CPhgYsbvc2Fv8u/xjDQpRd8eW
Ky2KNGUtiv2KFQYlt7QmWjN7ZVMWVPyxsrEhdP81lf3Nex7zsLt9hSKLKDGc0BEB+Mz3P8iypQsU
ZNtjQHiQcMnf8cM7rOzYMFZuUMuAmBV4UUWtP0H7SwmRGralOobQuVL2fyNcvdgLuds4E8FWngRJ
V6aqHnicIDAWKzdwn7x/QlHN3WM2Dqi7y5DOSPYXOBZngwEP5Magc/IjjbEanIQMtlgKvQgCbqRG
JhIrgCwEPEhLWXBZYs9IhZD9I1Un2v6TfyDE97AEnVVRBTF3faxyE3OxZkPIHE3imBXm1AQmtKql
cL2fPw5Ld6bob0cgRf6leTHuXGHiSoUY2J9W+x2QR9LBNeoaegrqvckIbJ+Q45AWvnBiO2GGpXqH
lVdQaA9CZ1CrrCjtgm9jmm4VLY5VRe/eLad5YvqXgruNkoW+hAGPpXQCc59kMMV7IhpLkIohK5qT
LrO4NgnRwzcxI8F1/UdjRcQdiIgSSsughfJo0vSqu40ksugQywQwu6JwVVimhQ7a7w7sbsX8SfGG
c2rcq8P95y8xXX6e70fR2WpEOSsQepJ5W/by9Dr9mlaf23fwNy2NoVXJwtZzDKZKOG4bcEWeX/Ir
liNpYSpmsCLdh976BuxhYKsP4UwUFsYjPeLxnNu5SYM5dsydo1qi2Y9y5bHDGKQV32zfU+OxW68e
RyvtR68SPJDgxERw5ianIvBxwq8n+6Y0fSIcbrP+J+b+eJWd4z/V8tLPFrSpZ68M0Y9Wj1L0h53P
jhH5WmsmArXiBMI815D+R2ulFyVLjyssk7d/PUZlVovT94UwGG7zg7g3Yf3VCAOqGUPaQQlt6pd/
dJe8iWxXGcIzDGBdaZHewoDHnZKbPfqJK34xPWddUUr3B4ZFJ8tC4q0t646vz4Zh3xx9TJ6MxZQS
zvzHO+6tXNGOHAL/2LbIGbNJtdopKWIjaa4VKEJLyxLjQ1cuS0BQ5d2m8nVvfATtyLdnNBN5vE+9
so2VO4MSr9Fg16bK/BktIam/qodlXfV5Sz5EOzbQUAA2Hdhq9+LDDW2ZRDom8QWT0Woii5wl804o
f+LN7CC+sUqX2RLYDUAFzXwJ3tg9jGM9Q9d8NmdHSa2cslTYG5q8IgUDa6LHTPqzfpsNxBqAOZSe
6FqPxAU2cq2bkYcCct/1D8QwIO+LdLFC1yChe22eKNkWjXhJBtwc8LTnbNfZ5z/MPn/QlRRGSOkk
UpwziyGio2bVWCFRd1+uEZ40kxrDbY3lLAzHCXMErHygB+CxDGbnTusmsYg3zOvw95ES53jI5glG
n4gBDEu8IVb1rZNuL+e7YaJfSjn8fZLzpZBCqYyEuERg0HMONb71mMA0XttlNuoT1EkhZ3u19/OP
DroBSmcGYr20cB9UPVUMfAosWwp40bebvUrQcmT1b42/ZzIq1Bxp+YxgTzJjIyOBy6mZZnG8AR9Z
JvJC1oxvG+7RYEw4V9cTwellavfOA+7spxXK6YTGQ2GdbESysGhpSFbp7Ab6shKKIA18o9x7yHJj
KF/d6qIqYP7XeTBGiCop9mqpRduz48pXFNlV0kyp00lyo8Ix0zmhn2ynUERStanriFIXANk7rEaO
yzIzlPXjAonWGSJvCJUyPiQsw1z2Ium27J+5ocRYwDROAbbzrgUp4/Mj0OYpFiI/LCxmBoEuavNJ
7hMKn1RJVwJabDN5xqr9olIcC/Js7I1cARyWXrZWioJfZ5qT0534T7uHvlxoNxeXPI/4e873vXZh
PYy5VhJlngrgqrxthM1JeJBdCfpmRaHHj/lUgB5tcMI9utF3R32p4Nc2KMdVy2ll8uPE1VxcnWOE
g8h89n6yPh/0+tbqMDO8E0IgG/1MhE0oRFVHjei3TUS6rtK2ic7480qUb5rJc4ga0NbWVSMImVFw
9TAx1nGqCJPEAxTj+YnuSB615rrmxCEkNhqQNlsynqgRHdFYg2oD8/g8J5Quh4ADEQ2VcNN/B/1X
m+Am962Fl6a+ve/XAC8xb4I3crkn+LhX2M70//7ZW1ZsP7wVBNd5e+o/oPFRK+6Y17NlXTaMunpI
9JfAVinOr7+OMXvtLOs3d4H0k8yBvRmdR2C6jvLlSHJlRZJvfkvOqLhdRaYY+1OMo9mFjN9/Fk0F
EMmcXkDMg92W8X+bHF/nWfJMtqKJPIDMFxjWLdjvC4AbO54AGZkaV9/6tR3s4lRiWyBVfAidjRWR
pUJQr+GI0pQ6k5wp9C6cx6/ZtEEwfJsbTk/6fr5FOzpzARdavmehBNAy6gg0vwc5TLbUJ/cj5EUv
GMGlIACzU99X5Z+2k7lKVFAzpYEKP2KR3tl44JpGngQRrLmY+N4jh4PelHT+Jj9gi2EsyESlkeCd
6PnMmXruRSR/+Iw3UhjXwARaR3MVo27oOo4f1HZcjo5BK1z64fxGzOscSKWcuDmIURyKyxAONP0k
oPOLvsC1Nk3Lw63IAamppyRXP+5aYfM/gs1O97yXcjg9FRRDxUuWrZRkzIkV1yDWvMXKAbdS85M2
9RaBF3uA+0Hmh9JptIsoepbyncAHZC0UHlQFmbfZINw6QvSIBXMvH7+LauifzqY3+qmS7mahbY93
K/UcQY2mCFXNAy/5+7j8c3IKfI5IbjDKop1E6K8beRXCNK4cRVj/yJ6EHGOmQUWT+/ARZcEyEd3z
Sj+GLEZhtYc3P2dfxaW8T9E7vnZd3d1ZQEerNGyRpjGZ+2jaB08WzvuN7dDJLZJJXjzArsUc4gUL
Q+Smd75IObIel5/kLKMRI7O3c2UKaTVtDcaIbcrKGNPjHG4QPzIpeURWK8XBPDXltrjvz2hCrPrI
K7mHZ2zPrX1F+epG2NdMd7cArBHKi4eT6Xy30hf8ccMJNBS+VCDJVHKnIfvGXqEbq0kdTyjd3Za9
D3ypqJ3R0mT8mFDF0DPmRrKVRqPOLKHJb1KNsPiCtf7M7/cqaua4YkvK/A57MQHZD/n9db3Cyx/v
ANyIZEKPEmkYgshLqt98GQZ9w0Ln61FZ4kPSgoUsTE2OFPvJGanSmxTxJyQIRI310j2St8rZtn1z
k3MDenhErJQYszGuyPjiXf48O11IZH1G+sC+k4ffkeLB0b9fFMEzvWCurkYL7LM7I9yxHBT6iUrc
zlgWWdRPjExgdTtVQxtGvwaSZBL3X3kF/up8WD/PWzUWqf33BfAbXoOAZ/qVzWw+HSN0aNg454hW
sj/UtWjWU6SKmRhPGqFnjWUmZ0aL7DW6x7gA/LSrwyncUTJ1qtmKyGe936ZjYeyfvqEW9XIOZcb7
ZrPPrRTSERagOSvLYqv1ToBtNB8xQaqH4UdJNI6fmHV9l9Orv9j/PSxLbocXt6kt6uY9NGtrKwdd
ND7dJKOX6sFNCElmWsWOkNwGQZQuj1lL7VfPxOJwgt6SsBKa3uUUZHhInhc9wjCewpAM0KSV2XqQ
srHIIXvmyvQqLyOQ9/wcZ41FD/sbN2L/RdIdbjaDdTFIkYtEt0DMBqFTTGwWBixynuU9283nITmr
ppgUDuzYULCFS7sjxs1usJUTo8bbqRZckO0MRT/qhTs8xnGFE+KtJywZgwLW91AKO8xJ4L8PRNw/
8KO3zEa4PSBImF9+6OYII+DNphUaDcu5NgchB3EuzOa/OHtQw0JSF9YQNTQXaLY1Dl6XMhVc4Vig
7hzxfFncFOr3gbRwY7y+ufOB9jEYRMarASUPnVn7JHG6m4AcWxNx7LkOtL0Gq4AU2m4HpF7iihaX
38z+TCTuZ/FmHHWjPQv7qguTIpOrYG+fnTRiVAII+7Ew0MQ6K/X6LeDQF8AGWtTQcCJU+wcauP7A
XSuQlqGV+cKRF2GulWW0KkQw2NKt1NNnXX6dCq7UKzOMkIBILHUivwUtn/tiNq+Z92aojug6/U5V
mfxq6DVltftWoGZFWsw84zdZFooNLOSBuWSZyLFh4ig9sNsC6eXMlwf13zuWwuHalFEw8xC9JUur
hSIohVe9vGFpC3t3ccB7X8f+HnPksA3UoW1Uzp/CLbqOOfm8F5qWGbxYv/OseEAAJhpnbcNah0ka
AkoevBWiYzp+y2glEXN0vO+ujVj1ZqQUeAuqRxq+5lma1hCiMeP63gdFTwVhwfLVn80OqxJKEna0
o2u0hPVabTY9K5tQ3TWNolegEQc71cv6xrb4tTPZIbYvJs4ly7WvKPDEEb6F+C4xKRWkLTHLCPlp
RgqZS+Cj9PRRaL9vCqfcwFn99M6zDWZh95jqGbKK7SK55DrmQr8appzz0bpEM54tYz2v67+AH0Ij
jXanSfOk+YXJweZeklt/UatYxWbg7Fs0hxdyW8vE7BC4obiCFXwbTLFWt9oTxhv77NzDE7zmQ70p
E/zWC7pURlK7LmLpZbkaWv7xYgdx6vyMS+txyYALlVGLnGqJsQ8EcOpcS94jmxECl38lsHVPGbRQ
wDrRhMLs2I0jsLGyfwCgP957GdcUG1HBbaczgU++4TsmxRo1tMRr+vX+Md2Vn4K7j+wK0hlkR4J5
oYj4/1CMNjCPJ7K0HY4AxpmbrKZkkYrG7m7MBGQsuKjyq8+sUxSanJwNNPBl++33Uw+kBYdzWPOE
fzyoq/hpafcelH8lReSpFNFcIcKma1aAhtoF0OgtOQdU28KBYMoWwfEIUmuOtAyIqQb4CSiq6CCC
+g4EKSQ1So7dfsxXtPaLO8LieYvZHZSmnoBa/A5TyYx4nX2tXxixfmGmltsIPLZYgF/QfMepLEN3
0ovb+KqBSn7uTHNOtqHMfr3IudPJ6YjbUJpk+BTI7iiwFehmyhosMxOwPU3HnJMMV+c+uoMRP+/l
Vt42+JKLY1WzkF4JOOhGrc5K1D76eW61Gjpwk5YUewIwZY354/qo/4LvmW+rfwG9KwL2V0zVY5Ai
NRXy8zY8j1csz6uEPaS6JhP4r45iRZi580YKK8EJeBFgo3/bqs2JQusUQOUX5UQFVr75Xn9OaG7I
0MtIB37e85Yg7RZpyp3iZY5+qD5eoMpNiZKdSDXFzcaG/PfMkyrexeMgPrrw3d/VUZ0TVw377oEj
Rky0xUGUZBdiIfxNJ5XOLorNB3YoiBbrPx8uQxu/qShwQbtrcxWucNH8orsbklIgCnb9B6wZtpL3
jm/w9seV10hAU0mMairLkFwSq+8SngJ2aC526D/quFIIc8psEnuvHOMEEzazWaJzik09L1dE6FQw
IF4QvVdaW5/Q01KF/+R380S7w4asa8GgtPweXlQ4y+4PZVRsaI+5k/INDDQ5wJPV4p7rk7NqJujb
PjwprKepSNpyueh2lLSCy7V3/CMOqQSuct5Ukl19FcnzyHtykchz5GO/zRPEOJBUfhppaPGgiPXc
6FthdILXPS3tMj5cSDYqWPJLZOElnbP/eobxfUFCPwB4hEGjLz7qEWWuMFz0g4tTZ6ybWleQcTpX
QZAjl78HdCI3ZK6J1Dei/NjgdW6pWLieWskQbUxEXVMp5oUIsQL74RaTW/3ToT6uGZpe8OO455RM
8sLWL608farNbTXjBf1eQsh4+21mdozlp+1iAz+0H9ARltpgDEQ29Z4fNTjvWVJPHpgaQsfpXbt3
/ooYoxI/BHuI1WfCrkvFfn1pnhcBlfuyaznwdJqwKmZResR+M9eJVkQR4/yMzJYZjN72zE5vNUOE
7AvdaAjTU5gPPt2VlgywFlzFzF+qUCcl85EliHKXaeBzMvpOp8eUIhLasDP12TdXreN6riH1aT0T
0lkYR90aIhBTsiLQzN2584EAG3cB3MirSYj6KibcST4uW0R1fElsBWGtMCeI3UynZBz69wI+MuQ5
gMyYbFn4Iuyu7ALOMHBrXCcWfWGgDNRWeoihSoqFRBd8+4ywOT6hMeeqPXWSocm3WehCpQYAToeA
nwix9T1To1V0Iez513W89qhuSzMzKD00dpDrVBsar4S0QqLj11/TJwLgCtlObsQihHMcoqc+TovO
JzROlsIWfKqBnjmGgefxPOLqBK2rvR+mZ+WHOpSzw42WiUDcArt0hrVzJcJxSpFwLOEzWn2OjZFk
Zpo4VDAU29RyPsxnh8GfVQCt7VquThahK9MONLD/MDWanYOffo4JFyl+I+PSUG1JjbRqmcrCIx1e
9zVA3a2po1j7cicD+RgVECbxJAqcHaXe8GoEHK6YsMpOE8IRIu0h/BWSZVZcNxyjGxvtIdBavAja
ZkMvUPhEw6HtNOLApti3YKPb1Y67t7sW0q/7ZFmx9VQ0SI74wP5cSmkv0DTRQqnYxNqcS4WoJTni
NNQs9eN9Uc9vnKt6jtI9cxC985iR18fbsl/Rql9cin/OgIu0Rm4M8iNTsRAWsFToSjWHnfNDNpTO
In6r9GrXz8LozkxXcZ02ezbB5+Wf0aSkPrw1ChB0MFN7QlV236/o0IiHh59bBUnxX1dsmbkPDKQB
b1dTa+UIg4O4GXdv+qe2cojMGGLJe8v+i1t8NITGIsbIWWIJAeiF3aDmBMl7z944Q6AuSoORY34C
tr133KsGwGEf9nRObtAPW1vpQetZUBD9+rsLrkr/FLjwJ1f/Vd6PdzHE1w9LFGqA71vPtOZZnhpd
fQ4Xk4HnLQDgiOhl8VvPolNKcPw7hligB1tpRkaKgre4TxSHwVBNN1ewb6eCBhTvDkWpX1cy5zZz
D7I/ldwMt+Nt31s3K7OCx1MA+pN7dmXagKvee/BUBFDEmuWsRBjXfaain0zY3EK/Jgwbu/AOvMJA
L8ucHjqYTYMhFIh53oFaDyZvafAzUqUv9ATF4yHmKIHqAfR0A7SlI8ruIxk9WZLcxSeoFZAEFIMV
n7XOfq0sTn6K0H3sumPIf898G+fjbDHKbRgOG2ZSGmi5yCSsn96l86+lvq+THl0AE1iLTyxRQ/dH
zWLeb+2azV2BMkZgWiIkBunCdWhB4kqkQudrtc9aGNgFyNT3chBcbykC9F63h0QCy/Jao8uMj8KM
LmltPJiUAa888RpkkLe9hlZ4q+L/mBq2YCUSWSGzjhz4O16hPvpio2seRCe5FPEm2x1E5ZAgG+E+
ighX65r021rUDabWrt2bbY7WJkipdowbxgQEQQcu0L14YHO/uEaWuSm0mSLa42tX0dB6xIa8dh8z
fk6u6QWYSUiECulb2xCR8IbpdAWwApuOHeQQRLUen/r1u5GMV8ls9MK83VSe6u7CZPu6kuxgXrdU
PiJyAYmJeUXkEdJ3yoOZlYhlktX/UUKosd08zYyknmlrAYKF/u6DOYOlYLBLY3OploYHoDzX8Ny6
60WBh1SukBP3ojGrdUYGcJGnwUu51Eu5FNzanDA2GoM5Fdvu6yHvYxRDwgKk2XIEdNa9IBYppvpj
dZmneDgRSmJ1rPME7LeXB4aChJLIFCM2dx0sUbvnn4ab4pACv9bBzpUQSX9m+wpCET5BMXhBOuqt
B7YHHsriczCG526s6zTkxE/JMloyKVf0qtVZpTfHCduq1JGP52EFlaNtxQtwGCcLmRhA1H/R4h1w
66AA1xBAhXOSmpFdJJGfG9LHzEEqXDZa9xFIVad4hiNwrqAKbqIBe6dRrDh3zBte4yLI2GNY6oLA
Ga4PZXBf3rn0nGjMtzkiJ3sUh/XApvyZFrl7vcfUweMkKptbelPWuG5ZREyxccyOmLRR1ze/ek93
1xMDSy4q3gnn2ggaaLmahWoqUlDm4BHxLp1Jz9ZDYRPdvGnfPocLdhDG2WVyM8qxSRmPVtFpGpZH
fnoFo97ItoIgX8aclAyJydJuCaBLvcLdgOF07BWBZUF0KdhJ5ZHcVL1560yRTK452XFjUMejdL27
c53NnwWBrIIujRb+vZKRZK55J7y42Po+K5uyzUnlKGFiz2CLaaDPq7gQFgiFDVWns9BMS62qiNAA
24P/vqzY9i9bBgLSXlzlyQzBO2rp3KZd4OsdHF1qtQZI3EgfDv/6qEucvo/FS+Sre88HEQ/nw3q5
+Wz6yPZk6qVLQQi4UpIAQSWzyccJ5ojOsFangwFf1+1dDHKYjR0ao8p7m0Mf5zM5QGq0/uLYkKQf
QLOpVkLnPAYHNWXJisFGDrHE9eqWocf/OiBg8W3kYb3AEi5yl3H1/0rDSexMPFF+RjMcH2auY2KO
AWYW5rVa0IsC4ofSPqL5Ryxny+xssG2FGvtr9GYlGvhi7yf0+xN0IxHBJ77xPfCTuZccGM9lPUyE
O76BeCFS1lopEXdsWh60WT5WyO2dmwNRk3XWQ6xSyqpbBDR9g+YI5IuPC/on+YVNhtX+wrougzqE
fSRZCc3mPjovGFaI/LuDFNsZrptXGghR+K5C857ie1WjOFjK0ce+pLQcZGdflyRsCUuiUTconex2
G4Wu7uJsziuo8LHNur1yLBhLs+Jg3+V7qDXyeXeC+62pgBD8gpEqkx5K/kWHnjhPiHcQDSHbbmXu
Fcbprg3brgQoXD8hzKW7zk6zzbFTKCQPL8lpd+0tXaHO3knRgBjTHg7LkMGHie1v1BLXUPS00Gs4
gonEiPNnMGWELNrm6cP04yG1+6CdO3FHwly03iks/qkoBhwrU10OUeGbsBnt0NEZsH+Y04Ug6MuY
kWYFrA0fCPx7HS1mvS25DvR6Hg3mZ40RtS6muLJqWipTUo55PIh/u3dav2aYpGAykBGHIuxrV8At
9smRiDENKe+YU7Agp7gZ3FCJKKTzDM+Gy06o7OyzdLIrRZAHgLR3E4HPgErR8v9AP7TqTimF4RC3
h6FbxKU8UKRGxXgI0NHOXbWxS6MRbada02tVx8iuNg6KajvFDNTmrbzKOK+qDvMPff9Kim5mVjjS
3A8rQq9suUsbUe6pZQbliK6U+QWReNrm9dpvGKvWM1p6fsQIvZv/exUo0XS8kZFqRdbhCf7jiIUa
fUmmnGFjT5TjbGPtC4Zpz+vJEEZdCA6O7bSYXSU2ul620hS1Yn8VJPjzSbdYsZDn34wt/v4iV2Qs
VkTOOgjrzoIZAj5Jup0k5JnR1wl69exuSTmEtstaKOMLI1yCysW7BCKezer/SAY2/lFK93W/MSRU
IChYsKJK5MvwcBwQmhf7fbnVOlcwQnVYmIYUhtmxeBW42V2kydAvX5Rbcym7CdIQ3eNure/Cjj6F
AmJMIzni0IwEgMk8as5doVHEokPNYV+U7x4zUVBxgn2+joix++bHXkm7KlxmRejOS2sDAAtTX6SM
+GbSFAWylSqSr0U3rfVk6WXHQwxumOjb0a5fNm4YvWrP4SNaAazk3Zn9ef7kKTIAxdq8k0WBfBlo
xs2WG170qBpe314OGDxIBKpVow0L/IDwwCuRtv64xFYqWh3zPUJcDuTs3/63DCrJO0zZIU9xesv4
3++ITUPgvEFVTn8XJZmI6uVAZShyNCkkgP1b5/WCXLY9/4foAdrYmm0jzBVCvGDTmbL9mxeOWMkX
cU6HTkWiJyN1YNG/+EH4+kEd6fQAqRy7xg5Ji6nxz3YpUVsqIpeitbUPVhPV2eNrtwj4P1D57p4A
3KVVFFjzlOd6Us5snvNeO2EFCiAlh2+rtlMUqwVCHk9md8z8RIh6645PMqxt4stkxYw/3s1cXmqT
G8jzDwE3jSF5XE4+xgwExqT+L/5MvkTbvpru0K6f8uy3RQt4sOUaG9PlZQjQKxO4QGyCMeJ15E8P
bTbtE+yGKmXTZ1RDXqvMLxLV6BZePvA9v7wzaxYmNPUkk5osWFjV8uLPmoeVt/HLg2s2VJ5vttzJ
cd/o5+4NmrmXwtKGdKp1BSYjkHWMaVgPSfDRYjUkKi0VRkcwTE0ogO+znomZ/GlRmkAIPJ5ivmxP
epvVHoW0XTCzgzss3YOCafIkdXE+sxX9p6HVlrD1j+E3Di3DixFSBTqtwqLjD2wB9TRduXeGwuOc
AEYtc5kxhyf1qRdjuP6KWBLHHavaZfVd4UXHMgKCzwVKhRnG+VmC9CDixm0xBN+g9NE8kQRq/K3E
/t8DIpR6m/Z2qK8ONYKxT7ErYssiWv3Fz/CUNZnMqfwFkYrEpu9lYzIq/nMMp/iJ+SpleP4ZtcVt
NKptw8wftke9PslAUnzsCbXOOdzkXVFpuhWwkcnDJKnydPjmYkAtvBA+kzxMb6+uKQ3EMaBNNJ62
NfstkD6V6bbFLwd1JPbzgzSE6Cf4OoAUrBzzkfpS/cyKGDxNbJcMWb0MQ4pYSOFl/dj5ILFRmA7Q
QBYBDxtoTEFZ3HqG04Vr+oHv8dHhWn0QK3LadoP0I/5/Vj/UGE+oa6yFDYrpbfQ0gAQ33S6OvgQV
URP3198tQZ5j0RbktxXcINBC4eXhvfAwSCJth+yty85sJ9/wyBep1B0Ks1d2Po1Xhfmt6XgAXl8u
mW2c5m3S6ZgMnm3FyAB4Agteqe5YU4SIh2AlIpLwUJAYDirL03zshf04YjHflK08JCBX1i9ALWRl
zlTcqs4uwnmv9tJQMtJzOLwJAevOG2/Lc4lph9lNCB9hYymxEGY+2dNWHAJgBzFH4rV8kiTX2Eyo
o3NjmbIr7u1IhRS8kpZ1wBtMQBENcJYE6yYIw32MXp456rQ2Kyv/pV3eZ2TyAi41PMD3y0jM+bhE
zgagbPqlQi/adIJptvu1ZRxcdm/Fam+r+Mp5+yZpfCZmMe9z37UJIGJxmLx651kZP4810jvAwGm8
wrH6yOeuK1M25EyPKPLenSc8T5lYhGXzlwSFr1cUEFgyqSEAWdnCkCx5yA6HsmTEZnAUsPmhXvRz
fi5+9wtU3p8pQYvhERngeY+cFtzrhbYwQ5/QH+lULQ+mlTX/oxRcvE7qK0ywsqFZjVGoPm7MJnyx
hFkuv4Qo6WSB6x7ofd+BeykEQC6GUKCEM9h7hLutrnMaXVvUrzXbEkcPSyN71ISsEuNllQnJ3mTy
Xv9DiMa4JXf2s8XsaFZdtzdU77PPWOdW+xUfmowvt790TOyJEXg6q6+lpJGCtmrWByI3Cu9mOzf1
QSwrQ7hTuH/Tt5Cv23g5qsvFk+0xJx4QzZk985weD7M3wzs2QM0EGK1U4ZqmZRErSnQ3KLF8Vcet
DG5/Yu75zUnOTDYM/0K3YrzGSh0pknS4C0RVs6fymClcjYtDN6SkDERkywgXq69fgaRyJNocIKAg
KU2fTgiQ5tKLoqL6G3rg4rgbBrFA2ssXDPjjneIdbLNacFww7Zo/Kx1x8OeGvEhPtNG6+DLv8rMI
UViswLmqYi13rgaqqSs3og3b6BaF4U+m3p2BgyoYHWiCjjTJjXnlG0xwptKbbCWizA+/P3l0w2dg
Jcr58RSU1mIlQCkg4Ea6aXSFbqh4sH8Tpkq3vNj8QV71NlWIcLwypE42m58GABzrWPeMfup6EXXN
ouJRCG4RpLzDh5MoqHcOr7e2ixFFfpoodVI0dVJnFdsfqfRp5jejPt2uRXvGUUQdQJu1sLwkCgoL
empCTy8uepoQPKTTPREx99FaaFYJuWJXK6M1y3xZFAypfdRxsJPntGiE4g/3Xfe25vwglRohwu9V
jWR24Iw/bPKKnLRMJWFAMbeiJ8Qi6QxQwBdbgrulKAPZXBqVPzqONgHW7iqgGYz9IuOAGZf5bMB3
+FABBJzV2IOvinRaWXVADtKY1qV4oM3L64vzhUO7NTKzoh8UB3sW6Wj7i1O8xKdSfp83mTaq0N0Q
HqY79ZK98JLcxnEIp/PjmODjt//HJnCpmqWUwPdHIM+2l+LfvH9KHNRCTxRC9VrBOwgLFILIh/oK
MEk+/SEslcE1gUPROhHAKDGJ9UVxTJj/X5aqKSTW5QuOw8Mqbg0MIIjvE2aKLI6nYHXYleN0CIon
gmLtC1xlrq5GKX+u5Sf1RyxXWnjm0SRYNmVkJioG5icD3+bdyNIlDav6PGXOMkdUiVY2RwNMMrZQ
vevobqetjXK9Y43n6hYgRMtyqeV8g6AIt80I5I6IcMXAZERd9Ni1U8sQEyBLjqRvO+2dtXUJilo0
4NY/v1JVr7K8ts7vNOcxupJdF4W59uyXWw7e1hugatKO7i+ApbsIe8+BF7LylKukcVD5knpAOsOD
qtWWNcLwsDeO3ofKwIkWTuw8GGwzgXvIccp1x/Bu4resK8nR4TwLBCrRat0qNW2R9tb8eqJMzcEV
ej8pN86A3nF9LA8WEVeW8yDTxfINuawf7ZB2Ock1v+9NNAzxB42jR2IdfoOlgCdH4S6aBN8/zcAb
wOnprb3BIZgdPkgTc2rGE4n9wkMtJkwB+F+YwuXnZcAR9hNXgANqIF3vqNIfYuXUcoMlzA0Bvfgn
LPGOAds9AgXrPpv0ZQ2BBN9WzZL/glambff5eLs3KIuK0d5KnvA4PD2HMfsBpLZM4tDGQHo/T5NN
L+uYc+d64gS3ppJpevPmkNM5XVquw1a4aaLcig8BpB0hpl+5qBKiEr6Qq2wOWHCtmnJ23Zir848q
UFsoY/zF8HdW9DAGMqVKcwm7IbjFnESDNLoCs3UR75q7DHAHLb+pEpVu7EpfVxH0w/pc/6ucaRzL
eRq1lDedJlXvCOUhp7sVRh8IzSytm8Yg+7t4X2fMYw8ULGo+8pO36OlzIUScFweZR+tZIfXn9UPZ
92x/vL1O2SAQAl/6PlUF3q9Ab/0+OXEAtVax86wuowQISSGRY7z9DDj1FlZMInDw+bCgf+Vc1LhH
i+Iw/BX60vrppIIQnbq7qLIaq54KPt2d99YgzVuZks+W+ga872ZZ24Mpi8EREaKPNSTDGWMylLbS
MKIIAXHBb2qm8LRM4h+ZTta/ODdkyyh1MHLS/RzqObPwxHTbGeGgdh2CMIAARkiApF8ankoDO6tP
6gENh2Z27CahgyycP8BAFrhaaizWgyM+r1GKmTKrWiT1DMc2LXjVLCM5gjAABfhTT3UEGFLLgj6o
XMiazB77HvOzpRGyFhf6GuBF3q9dsyBCNssnkf1lP6FdohGOs5SxgCHdEIAeDChrmeHezTxq6wEq
2XH+mVjDT+HgJ1neTeboJoHFQQo62f42mI4INpz3RV1G9Xx8mDv6EcxUSY/vmOQwRjbxWQ799Sfd
+BtoggAbM2CbmuYXGWFOL+h8/p52t/YGByxcJPgffBbhEbVB6uILoLw+eqVd1K3gjhXaI0eP5J9H
dClloKVaNQ4FLGs12rgQ1/GPZhsTEwLHKdPnjqLMr7jNVKZYOaOHM0vQJVYHz3oTUCxf9JRnIrVR
pYTgKYPfiqdF57oUJ+3fExohGQg7zYH7yArBq8Des3W2D3wC51ypW7yK5gVdMuShWliv0QCzfEeY
8nUP1hfWXhrI+nuZmrgstOtOJyz3jzFJDAcymt7lV7tv9AFJzcd5n+Hh2mdTDpY137zVjikyPdbt
TrhKeVxgKwxaPQDdBvmtkcxBXVlbon50tpOTWmMBIteY5WmXE8TmykYgobFsw9kkiZS39nnS+LWu
NELqYC7wPJ3pTktJb69EkwZy31vPlczbZLJoT9Mo4wIJRZJW30bOJjir6f1i5kNZ5vsd/Ge4ZY2h
pgN6PhjH0ZUYhzoAtLPS2Yadp39s3GPFr3qvtY0/S7nBsGyC5JsZK/6C+ux1QPbxH5EbwyvdF0oN
jbXyC5cn6fXMekJ4ML3Rfu7q9oP4Oi9T0I9E4fDwTrLjXnOctTXSkDH8zoUVrEQ5IniFQDmVi2K3
M+fCPndCnp1ddpbKsfhpaWKpnF1p9d45MqG6TS0TFYyJoI701LVI9kNCwrXFztpc+//RTa/Pz99i
1lxAvLNwgpWLOQzgrTT2vJ56MO0SR7prtOdBYY1kwybq0hVPtyGpinWFpLSQmVfq9yAdeS8dhVWr
maH6ohET9irgczC5JeZP+xhKO5nSVQlTeAcIBaNHE9j0i/rBCZTim9yuZKX5yglQeV1Xp0KGZJM0
KIHFztkVJk33kp5Vqq97rcFKTvevJCskt5N0R1kw8c14AByPdhl04JEnNHYkA34khwC3501Q6G4m
k3CuKyWbc3cWigiwj1YGkcP/okbMZTTXwYjLNDNrXFCqjczc8+KwlW6ytxpMhQCE1S+nUZr9ZQ2i
SYnqrKusKzshCm/esrzHGxhLrLUxK3mtYJlHCNrJvtZpHEjAXF8GkoiP2u2+vBUqzK/hj1j3D8i4
YX7vajfT7NlpJyuf+mnaJfOy4obcLu+Iry/ix1tiXjJjbCJuXxxkY3a+t+K4rNyJP2UB519JBBoF
pD3yHpJYAiF9P5vD9rSDrhuV1mly6LG3ZpWLdO2AzbQf/9pE4I3zMo7KrjWTKcOHtNP2Ypc+hmBj
Xf07kqzLHrieKIkogkHRGoPh7VJUAZMblDHoJyghHPqcvSDVHxtwXTtcAQ71pLw2OPb9V/5bCME3
jtcWrgrb4KPSLaj+KC5QOLcjZM70Y3RKJmiYLZ4BcqLcJDgXmP3CtbO7KQ3HRZrbfByAoSaSnK+F
yDS3KsrZnWzQsXB6ZuhT5YsFxnvDcjp4PULtEtNkSuYsZ4/B2OtMKsxsNYS97V7oJBAL7L2fggCr
YcS0ZoG7mb9hWgRr3I0BHPGr+4kANehJh3fPq0hazlLbKJwL0NZ6onEhkTawmdseruFvOtgfFmiD
c1hzzvzCY/23cUISEzo3h/ffMW1zDzC83crpPgc9TctRXW2YM1Fkz6JJBrUwt4oAZLYHqNJw2cfb
jDu48MNwjwK5+2/8hJTDNrnLvma5ntVYLJPykd/r7xVk+ea5oyr6+MlhaUxKAHGhUGHGN/TQJFRs
5cbXnERnDhgTU2UO5mHXxVpm571zz9oHCLDa+v/hJgiSD+jhBBSdqD4z4LQkfdZ8e1UdYUMccO10
GDKJDMHlfqoNe2owGctUEY5Yr5+NBnaW9x/xWC0joA+SQUmTYmjUg89gb+wos0bJbCsSeT3I3SDh
wUkwBH0+aQ1g916i2uTowAFlGNK2NW4uUxjRB5hV3mN1UZnILEp2dbScwvglinOob0KmaoObrNcF
zmXaAph9YgSFiRWBkt7cLyHko9lycYf6XxNwo17kcrTVwTTbgiVv67ofN6uuVEjISQ701nBXaaV/
1qeWlUx6b/ddAUFl15JQeEkY0kKOx1j915S3zWQ2726XrkGoKWjjs943EAhV0RtM7FEnNo60rHQf
V1vn8+dbn1DdqhiIdQNc3NzJ+2cpje3vIQd2XQUVpUGh4/46rwZnsxqRkyhXf/IyRFdwK+hoDKE7
yRAFXfiDCZGghHGAtAQDpV0Octl4fxXzf2HA1WcdCpQ2aQcjFW+fqk85g0K2kNntzbyIBs6ww1ct
e+Aj/nX3HNpmkMurkJpsYzWj3f7q19CCCrSmwATaoEuAYCwk+1EhbhSBsHm5reJiS1T7quwNMFts
QfAU7MV/mRRV1+y0E6MbVWDyUEVtoInGWFu7/nJbLKcFfMeuZBn+RE9JLHohi6D0g8oElQEMikb3
01noBfu3yPxZGsILRMBdZ0NXtDPsuAjrEluzUKzAXjvMdhq0j3lAEXG1wUEx2+r1mKE/V2njyogJ
9kjwQf1yU6cHJpzsZo1dAaVg/0Fzbi6dzjJYuwMeUCj3TCFlgiAvti1Ed60Ovvh6gKot8BxPZpbQ
qOtzeOimu6NVmEyxHJFESHh4fLcB67vN0KI7QzWfgIdF3WC0aJc75T04fND8iLy+L2BuHfS8/uqe
WC7xXu2RfivF1b/XfehrqmVRZ7RKEW+LlocayBNTuX6ASD6ewk8yrShjS4mMszmVAOc8Yr15QaTm
rRFn8vhM/p9zLRaW9OZQuYZgj3/tEwe6dYeEqbfdank7H6ob4fDoWCq+VwsYaElfvqyTzlXj+Fim
BvxrgkKd9QJsALYx/IE3+3BstplDoI/oQ7di48lUgh+Rdgl43VJTYiq22UBn6AIssH0cu2KZcLJr
tk1HTlPvGedI03I3OQaswfmfEVo4eqTblqLZmjfjFBs7KvvuXAFT6n/wiyi0Z9qAJ/NMuKmm4BgM
6wsQfI84WWmPkNu+SGirXt74uPgRFcr5N04ojnHiwvdFf+XYKJmSdut53wUKBiVNXLIGqsLzwkcS
ljSaJc8NwNa6mE3lsiSsCqqzEIkpHHrG3ys49wf/EvH/wkwTu9ZFEnxhxSZVGXt/Rv+SsfaOLsAo
A6Kb8fK1AHzLvQV7h4NKRXze1ovAzZLnkFbU8BXfhSU5q2hakHeEJuBjQDPXv73jg46h+klrDx5/
5VJ2OUtw0YUDWM58e4f3O223Yj49DYrJIyu/8J2h6HBmM3RFNQKm0WTgiabtC1zU6rZdyOrU0pLk
Dolw4EbW+0aSiP1v95F2hc7Vjh528OvTJO5FVBUGx3DV9PygVEYddzmLV3umincjr5f6B0BbzjU4
/paUkHOqjmDz1Q5KBooXqhaaC/feQya5dP0SZT6djdTchALrPUhR70k7kt7WDmpdZLznvg5659NL
IOTVOo7hoaNiIyWiCwQ05assxeYZxqxE8C/Tf/4rDrcRsIl67lKVqt6wswS0VVrLUcBujioSecoL
ckudahj2KwGODHxnbCUFAHlw7gfSSIgvxLFx/1pC9GC+njxdkxpIBQ4bTIkJDXBODxeT9OGw3cwn
DCvoF54enuTbVCdfzkw1wxzp4sYV5/GJYWs1aWxbodoyW+HvpxlS7q3RAJPuv0FVMBC9VPe180Pj
TJaVlu4n65GOlNMmfce/vifzcH87N81iVhzdPLaFtLG6fx5kFwLByiHTtl0byassxopzfL+OgEl3
NELltLdRJ2NYhX3S1WT9tbKVwFOrxw5AW7HRBobjjkl91luJgfF/Px3nlsOOKKIpzo3l2a0GhjJH
Mwchd7VWd0FzrdAsOuo8NmFcSIPFjxnJvtUYaiKT+5syT84xAlKtny8iNy52dulOPvjbbj4z9PhU
0qwmEWvXNRgr66e39tgJ31MhyHXb3j8vVNPztcvXUikpXNATQ7e3n7GQwkXjEr9t4eKVmbpZP+Mv
N9ODFQNyptx50FcZ5voZxcW7Vcdp8m+JIjJlrBCMJMwwlCD7xxekoxKbHfbbHYOsFWByXSFl9Mr5
dFeBBr7q8RP4X/idXqdUjfVT+V/JUva8AoqJp3QG8BKtZCrEvF7N7T/NDY3ubCSsBjwv43bJxKQx
TbO1isJxE04nM9mXZ/jWgp6GSn6BL91nvYF9x5FHIF+c2mz9ivI0qldBQubMmq5MFTRXLr9NmSd3
JgMlGwbVlaVJzUDK7fVRvDOozxlL2v2DUqumrzk92dUr5v8UnAhAvHT8LVzC4+jCl1ue7uPJABSX
nsPv+JyM0RwS30gwnH9r0iPecl3Boz5zIL3AKuBGYY6FwEQe//MGpJlZ/+SanEBy0f06TcfoCobY
d+oVxzZmbFsRlnrhijMdMOwLAlLdTaccJoa8tkf3ExA5HsBsa/JqzVhghJ+nIS5Ezf+5M8cBXQej
qIuO/W8kXVcwYGbiFXia2N8zvUddIiURNFP2uY3db4w5XeX9RzX+QvS3qTZw8iDtYccff4oSJ70k
VdXLDa00NnSOynYngzRQLZJNr49fhB+RVT/G0ZSx0/dWWV9RRteR/VU10Ivy2Z6A9GdQAc5+CcOh
jHJGICz/3rx22RATleQ6paQRS0HNW8dsVz3LrQEJxgS9bKIvpM+GQZio3cC2JWEmPkrDnOFHXUst
g6GsAfI1iBwr4gOyJ1H77NLJ8RqG62jQzXbtw+p1NR8lenNdB/0xoFgxmnK0GAFh2VCAzjPuAGKd
ffG7WCx1jSUd0NzDNGaQF42Z1iPLWgtcAXs+/Dc4azugYfmxyCMQ8moE3quw3WPbtNDMzOO7joBJ
0Sfj2AoooMV59h1Mqe1W7V9QunNcXbLx5gzkwwO/qpVrUn5yJyDLt1DWOeL+SPHBvgov1p7jBhdt
IXImfSq55o+kl5dqtMKOWYni+PTZUf3ybD11Mc+L9vVhMTiZY4gHlZCoGlx9/AEE45MDjEmFv4BP
7TNRVcElCq1on9FaX7vZkodSeDhPnoJBY3RlLVDA5/ZSUgIadZ3tOLOG8D3b9bOc3f8FZgIhQcEU
qBXJEHO7YSERGNn52b5prsejlHavwRqDBzV1LzFBF669+v2ejow2u3qDkJIPrxy6Gi8O5ibXBGr5
j0BzfQrYgDXbqwUKyS11CnDVqgZywXW7l3/Mtm3/d+tPbsRTKamPjaXUqgnlUlsxw38QV0sVYhLt
oGzmGJuhz0ZB1V0mAwp3VJmhzdrwwlUFdNpeZHq3j+ZXx8nQDvY3sZ5NFrtBkyxqRzgv95TYfNB/
brGYoC1cf95iC3kLaczr0on0aj4iJ8tfZV5WSv2bx61z3VhjL/osZrzbHG3GTrgAeycYBrcv1NwK
owD4czKBGMZKYHJVpk7HoPmZaEBVGpuVnlKqb4aF9EIEtRb91zJ/Crz5yHggDpy2xi3bNi0XdgKp
N2AhUJkK5BBjCrC75VrDofBNSq0l2zjrBf6dKrx3/wZz7hodOQfV0uI29uruxQEx2RomM9khFod9
XX2yoRP9vj3vtVDhufIdhMejjfnk5T6IBeToCGAcyEx5cGaKdyWjujYj5fOw2xm+cZc9mxTX8N5S
Pg/KdUiPfxQ0ZuvnRJtrYRfAJYhB0OzvN1cfg/6gEp5+9iLMiBpr63ykkD4lTO4AyWo/VFwdtkmT
OkgcmkP2znxt3z5Hbr2RkXkXkIvBwc6j2lz1S4ulNA8rHryN2G93H/oUeJUrHYENdsFNnJv/pjP3
Eo9uS6XuOgTj/y0MhNpdppV8DcT3OM4nUyX1srzLhwkbM8DcAYcZ9lFPZYvrY7cL8F3uosj5D/8g
mHKo/B0ZxehQ4yEbYf4w7PbIhvzWToX9rsSkW1I05h3WDJB5Odzh4MZW6EFHosDGIUPuDb1AMdJv
xWIZA73aK0Tjm2GBtNLfvVCJ7gZrQFJ7ToI2bNoRbuO3ag3Q8Lp76gzyCBrvwN8xbrKtHx0zeO7q
Fr+acMvhjVQ8dPsnqY5fAad1tuZHkc85T2Ga1WWZ1tY4GZiutEt7C1R1IzKjnbIli5BVM1mbEyvE
gSDvvaibMGOPGHnBnHTHH+zDFQvWtuODw7O8mo5ClkPcMQs2U7bklcy5Dg0G8eP+H3qBAV5oWuQs
ASL4sS0WF7cuQctiJmqIIG4ynxzLjFbUZPU2jvYGRzxfQf49MJZfhTkwKOHn78x/H+G03WL1ZTlZ
ljOjz5YmwlSdQMRr5i/5GVufITwBnHRJny6+nSI/C6iBzEUnRkg5xNUJgB1Byb5LHodGMNiSXh85
dMG5k0PI9mGsrxUwqxD1AZlGVl8eXA0N8UmgU0LFwG/IPNez1wXFDzGzj+nXQFoz1mSNYGGrKN/G
Nq3EJIQRLBZu/pViJ5pVyQFJtmrAbBvPjuhOVDXcLA/VAuDs8df+38PhqBusipygN/F5ppnazUEo
MdWg5Hb3apIvZu5AzHOaQa0h3lad9kRfx1iiRpBef8L4esAXvrnjc3/waYWqZk6XNd1kn5xJuqdX
wuHhmflOH/xSLvOFySYLFeqpHdH90ZfZ+yFMY90+171VVsGUtrMbwEr/TeVksml0AofoC+7I53W4
ddl8vdZ6HmzaSJgerBhyJTZwedik9nIJGRwwygHGg0Na2HFH2wSn+GuPROYXsrfOoIcJzbJl67HZ
JGYFHrU2y+krQZ4j9B6eGjZvrB4smO/3DONRUPCBwYxIzZMlGJmenCLHkrPds7D9c/8iee8EKTyF
zOLCwjWWTka8pge9pfv+ugWJ53nS3rsu2CikOxiXpnFn1MY6PouxdMvhVXXWKhX5jTw1gVonryt/
vz8uiu6wP0HBBXZfEf+OeIZLhJx00l6ZWKDqje1srDWojdDaF7xvMZzF9BoqRRs5wn6zrqaYnC0T
DJ6xvN39GOtc0uiiWq71Y16lbVuh4TZrAtvVK7OK3VPAvaCCEt2a1jNqJi4EDeZTY8Kmt6hew/G6
mGobIu9qm/zYgL7OQ+6N721WDqvcxCkRbGyhxM5LhrHlV5koShO9FmnMsengnOzhVtJ1jilpsVfo
5HVWzL/R3ZY2RWhcCmWp5mkHylk4cMy6qcTpzvXJIu2QyMnII1KLdLw9hKlY1e51bbNZdqnjsoIQ
vMP6BWBQV5HOumzmZQwxuQtXRELl6Q2mhaaqu6FQpx9GpBZD5bYW+xdIhISae9za0Q3ht6JnF5+Q
RPgx96GSfKo4kOuQXerUKHCrfMiCbkLan9+rvsg8xVr8lF1C3KDhBPh+00zCR+kVoYVjqoEVx7LZ
S1gNVW0t7KjeWFFdJUJLC4yw3Q870lvFfFIuYAy824SE5wJcYmbwWY610NAghvx702c1U6cDuLNS
gPEv8axB1JWK7I0eP9qUzX3xBhHw7OeWLSao5IyslNJn3J9qkSonDSNudWb8bw5psHepIAEe/ze9
+7n+F4aldLJHgEIbPKkbgTWfzKBY9pcR2OIpVuHoCVQ4/Zbdo9nuhsI0fngZHchEFmeW/fUwpF9E
Gwg4NqgGxWyBzhsItip2qm4EVI87xRsHovsbtuAmSf7Age6znLKr+f6bPSIPYk3tGB/tetAdV/lX
Vkkn6OvCNDMq/ZVz5/CLhMd5z5LwyFhP+adw4Z7qIpiD0L9QyHDi2aUjRSMSGQevkKvEsEwNBQG+
1BsJyP8Q4aVDYahFb7oy8SBi8xSRW3Rz3AzW+EFaeuiXWrv1NcXAMaATt2qqzXm76k2sIs4f7exE
HPoEhgR35ZOLiOkGgtk8iSNANWFAlsWpod1h6i88ZEz2bx7QNP0mEifK2G3sjHT2QyBc0Iqt7GZD
5D2B4PfV1uh/hMkfCyPUcUnypTKzPnE6q3yT2a7FG93BR5JbSXgftNY2orM1suKBkeIm712J5db4
2VeEi0nzryFXBK0skiqkpNU1NJZTV8OHwNCJu8UFGOFAOIoKcMApFdrGdjndSgiQvrV7R82UeJ26
xpkfe37hsAtdExmgpDNoQRGxUB2ItK+iGRlbxq/MaqDkZd2czK8pPYBZsRkG3HPCnt3iD+nv9cRh
cVMicbvEJK0WUo8tp7RLpkR+jT/3L2F5phLIXJvTc5WFYFlqODitrkwC+B52YEDsJ98zZ1TRyjmr
7h5ZvwzszHS1mv5+hgDyKqWZfNIBptn9lTc4x8HuILxk9D/6RvGaGB4KENVmDyoPf+X6g4kv2Ks/
uzIDumEJnRHNhG8oydxRaSoGB3KLtlpTtiOXnR/gPRzu1hW8S7bzchQEdktxFP3GSbVTE8yu+l9k
KXoCBDRxPCxmXrQT2yB3/yNqLlOsRh0Lh3dHAKZGbVIQuZonNBkFseJgjhOTzIeYcXZJsTv+ufM9
0XE/tlpZOQwBJFD2WvPeGazj1F6LnWf8+IowcxRIOm4Uy4nmu8hkfH+69qXdjz5wgWhhRkheAqf3
UmutR79mWCLYJQfVn6XOW8H5bsIvhQD4p584PrfHgj4AOPUkGISCC57KIhox2kT7xXsKAbx3N2sx
mlPt6+MitBaIZ2s5EC0BPPXz07OJB+etwsrMFpa3FZ24NfyoEx/8tC7x0zzrZjQchtteTHXd/3GW
foUSw1wkpsZbrW8Ghf/N1wk4PUkajv7xmrMtc9UrNS+Z/UlCukLHQjzxCNj6ozIVrffBmtqlclY4
SIqF8pF+DjruC0Tuw/9QGXbS3YSv1LdyAyigjwN4ufTH8JvbK4fcRR3JLY2/GESC0My0g7p7juHG
aisKPq/QucsgfIFyMTkAEAgmvjH6m6uZi0Omy23X7jOgzu4eBNHDEK3in4KooQW8dC4nG3r1DGmy
6k3Z4Wj8PaWixpRm2zTK9Fzo9b8HUS3Cvi+6U/f220TEJ2zYKK/rM+ZkUdfZpDTaFxAwilGyZutG
kbAC3B1bwIaennYx3fhlHk+B0obMHYNlJO8pLvgOPahXXsVh1KWsbbyEqz91pv4RDRY2VyfHmRoE
VQ7n7bFB7OQqo/Bpgg7qhppgJb/KwMctWE1cs6DbDZRfHXuSuUxDWRS5dsfaU1exRfSqnGrEvvZQ
qR3iPnWovUg1dcajaEp42CUXPwROpnJ54+iUgoAW0+Q+YhdGUs0fT9pHH3QUgSPNleshlNy5aSuN
pc/l6RmxCiZizGeefMC1BiprLnqxTZo2XrE70WMbus0stc2QxhcYRPP+mvnnclIVJ6lWCfO6hZww
bML7FErAuj7yL+CEIDlgkTbuc17kIFxzsc7uAwl3+t8UokysNnKYSw+bt4N5X139/TNRB+xBqx1E
2PEl/7+2jWWWcr6sz+35SccsDeWMnAqRFUoUTlLBDB8kzFKVl6AE9YuLVsHpA0F0VN7rXtvtMuAv
h+cxLvaI2jMynG8EnpwanlgucOAkt4nlHF0dIO5k1VAuMK/eCIpdqMhNQbRjcyAjzaMJAg0txj4/
dnn0x4IpbDaRml38+Byw4sx1Zzcx59Rnw4wQzR+rgNLWFBrI2KHnzAn3D/Em4Q5utVqzq0Acozbx
MfgNeazpZRYhMt5v53kbiWa+L8mD3GTfJz7ycwUQmaqS8pX0WIMCWtJQdigLWS/h0iUK4pj7+IX+
b5VkFC0JqzvWG8llxfPJCBLcQjRPYAbzEN6g4gwLpbKiZReCZs3E7IsEv2GP7A0wYbYVZ0GfGJ8c
j8BiC4/P7GHwF0I+vg9mXCxWRybLABbP9Zzn2B202NdAPy1NTbzD1MoM0DYmI0T3is/l+Q8GUAit
4Odkp33aQxn6t3/nM9Y5jAXmHdqj6j8DIlqmexguI+kgwb0u+paoJ9KLd5NYJ5x67PVRYABZ/P7s
81pxn25fOubLAKN2pvgWZUgFVRKH6k+PQodXUEVNHfraDRwtQXHsmJnmaxRB/VY4lworIsvbmlIg
TS4UVGoAG0xINpxw/KH8n/0Q1O4PH7q1J6AjQPSZkWczAiU5nPuTymYMAExZnzzWDnLXvr+qw0H1
eVR6p2QpDDXaHIer8YsfOWW5apZdiPFZ25A1IK6P0UiI/f1slFHr9t165lsxGYYxpvVktJVD31Vc
4haUw/fIH2Us+fF8xqBGdMXt+Wa1XawCow+POLdOgQzigH+A0MhUGntirGcPq0X2wLQC9ot3v3gS
qdTxaXlZ7Oo6kai2A4Adl9kaW9iRYX0A5RCmJZrEQFqrXyd+YfRo/u0C/NEhgtA6UZRO5/NA9n2+
kqpfWpu9Jp1JPgxsPJmbVaUQvgH7g9wU5wvMbNFjMtX9j9bK4KFHjuAZeHtp5NqNyE4w7r0DjLNa
uTUbg55QvzqrRavnfIoiW6zPATs1X56w7EziqYiPlJJBOnoCimB3Si6c5wnS5OY90/NA2crFXe/O
MQ3azKBq8jHuHFg+nHzO8DtD4NmqP38TGlD5QRuKUk/2OsuBo2QqMXrOpTLFTpR6jrTqIExhIwOn
IUX4xYShe44jS/f2Ij57kNRnE3KCKvRfHTHzU1b+RIyiGPXKXFFHWb2hjXyIhjG63p5I7utjOBNW
y00JEGCcBajiEmiywYbo06eq/TYdt66IK18vzixHEkwB4zblcpCY0I/WDl67ukRV5ZQ/XL1FZ0zQ
2xqd93NMZ93KJR7c10hOFmH/SfoV72pCTOcCEJ72c1CqjNOR6tOut1BT3NF0jqObZFhFO9WGF6ZE
X6B7wCE3gFxnjX3soPHoVlWnmgw6OVXh4SuF+rTuj5vflC6ZFQ9JDWuADoDONNPmQZnREe/G8e07
RhXlAlRrZ1igxmZsGL6l1usTUqqVbj3qxfVVt+cLbdtrqNaCuGFWenuCQInAObSGwpmQO5E6/rct
nbAwKAXVMGHrR+EDC5qjqzIrusUVgbgieE0MFsMtLGRGKLswvn580aHz3d36Tr7hYfE5NOfBykyK
5LQZ9474fihWF+pW6pucpZP8DreQWYy9WBOTp+PMLjtg9qtA19z7CZlxc588BwvnFVTWfwFXT4v5
EjRuC1idHm00ShkkZXhEhLClB0ibsJMRkMyBHooDSCPpdOvrrxIPDOIOFQyH3lDRjupyIvCDrT/1
tTCAEEo1qA4qVZaL/8RaA9eOMnE3IoQ8huSWZeOVehyAh91lbJuU0/PlTsSwCpXkZq03gQjr8Sv2
c19dA03TCr8OWKsBXU0Z49ZOVDq9id6G358yuiLW8vc9entrt2MRQ/jP/UKvYuXN4iELZY7QbFlt
T5CdoW66flF5r7r17znM4uM6+nZ4xC1Mc+Dt/91WyLCP5CyFckVxh9XapwM/CLvFK0pLNAs0C9xS
pVT5I7dI3bqT1bLXZL4ZTuX39O9UsjH6C5fYpGoqs6t6WewrT4QNq92gk2saLUibAq5kSUiqn7OZ
FrGpxA404GWsBwSnfcsKBqc1h84ZvMEz1doq+qcAztPvfdsnmmXa89M33Y4vplQy+OrsRSx6lYOP
JMtoSZgkkHgDAxVNh6rtE3USOilY4SyzjP5ZWiMPCSbbMvHDG7uCTd3T4j3r8uD4mhxG5sFviC1T
P1Jx8hvh6THFRHi0Yw3CiguXkt3l4Hc7JNfqWVoze7UEO7mV3Q8tBQppRTfFIy7ZGBxB674cwMxY
JRJfsU7CJwQoEL5W0jevXHE6W+eSp0sN7jdFANeYpy5gq3boPiNjgr08zJI0nB/XvnZPquAmqjW1
uiN4sbB/86AfN2umBGVN8v3bHdGpY0FP3t7tnu6sRpKtaEzEYKnEdSaWP04NGhSXoE6Xl6+/7dgg
HMAyOhCqoyI239I4NRmUqqftP+qJAmhEukEUdOS+emdzY13spyJs6vz2PludBEcD3yopV7MHKEpq
4NFrPy5OD04AT+W58sC+bjaeV6HFWIqswTIGyCgtuUi+RuW0F32F3UZImdWlcwnG5yh8/oDMsR71
ghLPMYCqrlShmfyXZYhMXZF7OHSN6EjDuprgDBEt5Yy8kkH35/iSNxl7h0PBN+s/MzFNv61g2c95
m0Z0tSfByNDptA6PACc+L3bkX3KMUU/mmm514M1oVzinMwwbUWVnSnrTX/2tlq6ZIPO8eB9r2s23
e1GTu5vNAcZjyzoZMgCJApaVhvcPa0HGRVg73gzjLWR/tyQVSN3wEMKLME0xUQwfjXajp1zivzFd
7wtqqV3x8AtyYaNCKxMvBuwAP/z3ldO1IlpFPwL4FPGv8SHrthHAbXjTh4c3FSkT+S7JNEcjhTks
nXCVizdZPYST81/Y8Juu4BOtxHydtVHgZBAoD3IzMYPmHlD6u/SgugzWHByIe800YhS180JTmeRz
TlLImXL4zJ1HyD6xOOoCZLs2b8RxQxlDCOZWmY6Jmc47uoWaczlCpgUCBM17YT8KceS1OPcHtP4n
uqUsDvv1k2TMK7zHTv8nB8DTu9e32najb1Lxy0wxFXbIvyRcH8/OxoEkOaulBTUoI7QzFOkduRrk
IfDnow+yqPXhDA+YYzaXEzGc7KcPx1rQ3OLM+18sBL36aY01YQ7jT86fZTr5O7/V7p/TXDS2mMMS
YfnISqmrdgLN81ZCQoOOXouj1PQF4bO3AE1rePdnuh2/L8dg35djESRkZ2+SswF3Q+D5V45SAFO0
WVMaZ92wEfnE/ze6Pi/ufNXJaUoqvlDYC5tS5TtMUT4FwNO1xdk/A14olvbKj3ocn4y3Qjqj5MDC
1hRyeoypXThlJRyNILd4RKZpFNvLtH/0bC7QtoptPGwqAqW4t7p+COJ+xBAADEpbvExBPvnC7eM4
Hx883QhC44HLfxBdXfSZlHRVad2EQe1t3/fGhEEhSAJpAaemV8cPV+ODS3c1FSrzUj085KJyzdCz
07oNqtwZJNykW34p9h64ea3hMh56bUewkwvbAkB/4h9X5gW3VFcYTBk9ozSufHl+2AldpEaz8Fy4
bOmfzfgv/CexjsoC7vJX12vSZcJb0fEvsM325MiYHtN3GrakCz41XlSY/KYVKF7yjxbC49HOCdEA
aAvP7i9wmOQXYQSIRpfajqA4ENXN650EEmv6mrsWeSEpTLu4OSJPKv3TwcvQrwbQz5nje/slakNN
nwUbGmDEeSDYoHYhyCGjYYcFIaHv9DgXWYDwXd7Xgvsj7V/8OIO/OeAn+geujKhOgwn2oku5Wvog
Bcqf1CQ4UNhk8ulg42I8dfzU7SfxN9eKAUtbTxHqYVgLHCEpAlhzCfDXvwTOI8gmB1mEiA9vNzwm
eeiIQ+JSLr8F/ffkHJ89HXDbgQDUMef652NA2REnWe447g41jw+QpRUENHJ7fKZLlEpk2t2tX5K6
sr8oPFgtfsyM8kzo3rpuoogv/fPhFel4mu0eeZaQsO0YUnXbCajAc+geA+o2v40l0WJkZH+qzAnT
bqqlJ1I+KSY1JTgd5cli8i36IMuHObvwm7tvbo3HQLcLlKnNhUMFA/iY0rZw7JwKPswEfChN/dGf
Js+HTEVjobkTxXvvYF+S5Dijg+CgJKlz5aKGCPms+VWrNQI+PRw4EGdzKKMGlIeVOERvsDyJzc+S
BQ2nuKd4BHCzYodK2g6kf6JRpx49x0GeTJx3Bpazy0kR6p2y/Fxq11qCi3UaGwKDbam4lMa5gV7b
PJHHIeMbXjQW4mXMOBf8Hss+3VkNo2/lzk7GN52/Qbru1ROkKrkz21nu4AiUx9DtSoaywV2+HRbq
E2heW+hYsZOsrgc8ZHn8TXgMFPjJf64l1AAykd1LSsr5okOqXJORIRLPnomX9saAFMxd1JYmS9Oq
zm04iIBkSwVdkt+NB9yf+PbciUQtyqICDn0p9f2VEzaSvbk4za/pbC1gJ/dD4H7lzdbkGQvMTuYy
885jOFw2qhFClWJ76jIKGY8MUJGWuWnnewGnuEpiQtfDwsg8HoSM9vrbHOI90PxmmruVlyHbJ+09
MMqXM4nXixEajIZL4DEj00DnOZHzMVxjeAuZqEnWdM8JeZVE6f1Q61IuPIgdUnZ2T09xiya9UCFr
cGOmk06AUsQkuLPPELG1XJF4J1DFtFf7311FWDurM6DErZOCrkg8nqc1FA3+uvQ/lbyKCCXM+8tT
Pop1h5HRNRJbim9fUptu0SNxX9Nlg5zGDtOqpQfGbYcuIvrlKsGJIWpOtQoPb+qOLFODDyTWduNP
iWIEFt6139/VeEOi+5IoZfg+nS0ElLPbC01d5WjXAhI56QeiCvBuSX/JcuE+UQL7aB6Q1tleM3Mz
P6+4WMgk7MqlagILOyhj+ILgWD1SjaJNNS4K3MbiYvpp5BE0NRuXxPM8aaKzS/J2QrS0NHWAJCju
FTYwS7AFg3W/3ULl0jVOaOms/jn70SVA70mA3WMPhtwMnEbKIF4X5Re1CW8EuKI/mOcKZaaFuLj5
UldfaS7TbQKRJ4Ob0nizAaLumXNl3crKo3Kc0kzaXD9fflVMMMqaR+fYuzH5wTSId7NK6RCQ8dZl
lWg/3tnYl2dL1PLl2J5aVKPPpb8pV87JOx3r0Hg4cSfXLcAgrusPocfK/4LgQw2+FSbaj6LwjTex
0qSFwRKkvszEmHoadoCDMbQOe6LRvs59P/8KZGchiY9abglW+CwOd4UJ2T3AJHe4xhUQSuJn2zRr
7MKqAOMsIHY8pYhvKavBWulB6N+1GKxHQHUHsvuHwoPoL67eeqNuJT0uue3ICD2gD287TpcZ6tIk
A2++L9UoRulDis4keocK0BEXASO5NecseEyKKMJOusLjUOsghyq0ISzVYFFauR/NOYFemS99JnQA
FiAvY2JOGGkUzcQDtfiJP5EBp5uHv20aUIHjfKWQ54w0EQHplGDRAlaWRfcfdvbfTm0EhbSdjRYd
pYnoAu83aerILOzCtxaC8RzUy36zQpDSN4OxxV5i9XGHS9R3r3wSdulVP3dkKpnIlM0H2OClA6B6
BBFki7FsUJhdm4i3+SZyGgCTyRsoq9XYKeToqwBlr83qoo5sJTsBR5cwnDdxUV08fY9acjIu6MCN
MwI3ZQnf5i2csuqaDJrx4nF9TfUZ7Iyn/xxf6somAe3ZfkX8KFhh4d61MB4dLqdW6Uy8jxBgzcWu
8+gJLTh+36xrAS4M50LOpnrSLTY/4oQLbw5HlvHigjJzKJUQ85e7bY19zb4LCAvHiaPVsnkTN+PT
xMz7TsGzA/7BdxHFkhQf46QQlvB2PxMlIdAwtMy4nnBnJVshT9GThO0/gONkksg307AWNLGIrODW
9x6HHEveKkyIhZ3VTfk1eXKlp3Pq1unOXNNh/a1fn8GF41fD0udUiURbzuCiEaQDkj8cC8UG4Ae/
m8wDEsW9qJLDYLWQFqMl/Im1TF8t1VhqKflQ6rVrmyHL+nuxWttT7oUur0R44almsU6zoCXvi0hE
wvN80oR0TpF03crv10HLZ4QTudce33nrzUbfn7eFhYr/AN2FhEjDb3Xv25Fg9BLosocn/MWaYoO0
qO3sf0BQxmeVSFRUL6zdeUrLzUUUySvRFxSjaZIphHc4ssJboHLG0DZ8FAALYw/5RniL9Y8exUws
WCkD05O2h/TyBqYKKb1HRLnknoyVP84f6QSi8Q78yxgiFOr+pP1jsO1mE5DAWDaFLVj1zkwAP21J
kiRU/PdIt1LMu6PhyG49F9OGtl63qdbY+aMihrT+QazH9b87Yum1ZvKXDR52gMMWjr4V84O8wsIS
FDRbWv1Z/L8xRAleUKE2bYITLPyDUrBmuHwTtzslcoBxr4S4qd6DsLMoigA5C9Rb+XDsrHfuukWE
SBcUZhJsPX5HQ++Ja0wrz8vLiOqRgG+W3caHx6MujJELcU0PUHG3oZYOhBr1DN4e3X0e97GZ2539
h9rcI6tGFzRSw8q1pUsVqNpxydvrbf9WR+buH86Ym5kbJxRLZCVAnMiHk6aK9w2gXxmgVOdSnZN9
bqtuXpAotc700CT50wfLcXSTmlqWLqIcu9AZcmW26QUZVU+rt2B5nbycrNkVt9uduQUt25/xOpnZ
LVM4+OjecPmaDDUWAAAErm8sOm87OSOvOIiNk1k0snMyDPQAlSpCY7eFtyjLGS3/U08jzQsgpq7I
YsIf16yW2OUvkfMD4NYOLFClFwinXaxPfhrW6m4xo6pkKfxFK9pfmdnAZi1c5vN8nqjVNs5dsVRm
yrn68bnO3R6PToUTvbMOWLyPAjTmlFnham/rYtWfEW83v7N97fhlFkRDRHR1lwWlstShywHnxuhm
bvPqoSVS17BWIYn8/7+jqeBJatKJu0LWqu0YzIHUeJ6s5CXjt0+2fS0+G95Rpr+bXmYKifvS2yLb
HmUYA2jz72zbx6eceNNlsES8s5x+Z2YL9wJIfjpssBms/iNlzjzo7Pgud3aAQeDG5ejMXzK7g5mm
gqm8fvuUy9GtIQuFzamKE6mjkPlPNuRQiZS8uST020BKrsB13MmJu+DizDUxAPYc8cgIC2rzmsXY
zu2FgRivkGBxvdWfSzEw3cIfTCF+XB2AWVeqYrmt0JAY2L+Z+pgAu1StR+umnpxXYkQGNOhf6G04
RAZiOeybAHabHhmOSFdYccteEHKswi2TTvCFNVdEzi0MdbwpSGbRURBbHD+HnmoIdfccgTW4BXq9
usEIr312TfjThtmMR8PMwAvIZOTAJGydV9T3/8ftdhzva/fYv0rMCA8SpPeXRCuJ5V74HSFCz0Ab
kvoKNLvRXeCYX4+h0OGpYCZ+in9Xmd7hR6IhXlzwwflyx/+hrNHhJ7Xe6t5vx5hTItSPJaPzjlOo
LGQiYy/gjiuSHzAFYlmKNbaJZXEWsOH2BI2+4p96hSX2IVFVMTX3RrrjM7SxH0T9hrNGam6nFUBK
U1/3A/Wo3X2CSeCP6MUHZtdrCpU1XlNw+mQmFqwMiRpf1Qlv6ZQKXzx50PXBnK1xdMpFO9+W3xIW
RqfPy/NMFNby2ejiY9YHkF5EMGM/eNKArogxFxt2aG1OiNti6PVH+Q6ma8GDF/L+wgGIbJ/mkMWc
E0FZrO4JdmEUzYycauXEHR9C9bHKmeMbANRDr7n6RLMCD9lb4gB3W7atDSSCQr173vZDgdnXTuZf
EiqkupcFpQLRFZ31uLp2PvReqNRAU4/+7RCdM2DxLWQSkvdcBk3p4n/lxP6wHjtvvkCsj98/8MIq
nc4YxvzmVn1wTXmOtR/wsScJ9OIKl8AWZK4poTSOlVd1fB1RTpxFeBTFWam2Gwy9aWe3wO1a7x57
cjafL1hX4XFxlA3iPIYpXvevQKpvF8w1Gd08ahx6/1BmteK834vSei+uPm09hzolrByzLzX1BDp/
SoMoLXwna7bEqbr4H9ZslJW4rXqmuNohz5iJUS75/Ugn7n+UQVuSABmY/N+/JNuL3ucwYNUyTSLM
ZZkI5FY+jJSQyn6aH5DeAsMl+RDLrRW9V4oVC7hIUcfr0iUwBVnP+ySZk7xWAO/qTmiZJ64roDoJ
6+0y8YP1P6Eci6OuMT+LXsX/b4MCmXkkCcBaG79MMdcv/GXkq28AYb4YGFgQ/csKtY9gn+7ugvIN
OsZptuxuBYx/8xVqE1c5jjx9+fUjO/yUmQC8YZtphwgV/SuQ+h7OQCwcIMRUwyyEtw5cSPn/CbtM
p8zqEMI/KX2T8ZkwPIi4E9XUqn4Y3p7iyNjria8mAkd2d1bSunZj123sSE+eVnGoooQo5ZHtnThb
h9APJS+xmlaCVwmDas2/Uawtk4CWa4oRu0rTu9BvgwGunmHuSWlXxXrMEwynvtErXWmLXuPQ97CB
vqcXbEfgGByTTEEzx5tD9tfAudU3yQn3MdjUnIdVorOhHx5yWdnunsGtESWK79iPKmp1tuuUEKA2
4EtJDWVKQuEik+nr1mf9Gqte2SDXkrw3OBhirQA/d1r1Q3aR0tW79zyW1z/oGdGnnS+C/2lE2gFB
lpuvkXiVuhZRiP3p4sMXynwP2Bh5X8Q12aIQDc1AcHnGAcR5XcUXVTUWK/x/0jiMdHLthwkOqY9G
7suZ5PBMxI/E9KUx72Ke6JbD9f7j8H9HTMMjIZjveMiIrAALmaOK+FitFtYht7ZGEzl6xWDS+LO8
gqQBIg/YKFyEnw5YybqJEnjrHXmS2zEUtsxCxBhPWON/dQf/LbEMAVxWPtpGYoaS3YHMcXZ7JCgf
ammFDZczzZQ9zNJWyOH3R6W7k7R1KlJl4ByXEIpWpJxiIgAHEPDLd+91+1PLH1WbjJueM8CrODfX
COATAAwYE1tZdCvCrteaPhhMTtBpsNY3q9DNZyAsTkD4RKZ5Dn4xV0/NI9n1TtGo39bzuvBk6xqm
WxhAy2ESrf8KTfEz+FG7+51TXfhaEjNTKhs4DDyYhScntR060titMmxtAS3lPkM+lftFrQpkAuTA
0X+TrER7qq9SsQV9lrIxEZdMFLhMkd5K9oKmz233+7LPJ0fD1+oRhdfa8oasthUBYSKZ0vRZ/u96
K9CVeb5rMrgQKp1O7kJcr9aKAQLcS2amYfD3thsIz7RghL1ST864Sm80V6behJrOYfTTnwz/kDSw
1JvFtj1xAJRGKXPRocdtRYbMxbp9+vVTKN4PvkLLPUSOSYDGDhFZVKAbLJKGzBa3aTdBUOyUCKXV
q7lIrINOgOGM3VZObXzunH30QysQlHH811iwmrshUEUmCfDykeoCkJh30eQfiL3Rl49+sWosOXxo
hJ6xjV8iXZTnY0XoSOqr5on9cjVDyqJza4fPfBeZynql0xcvL02GEZc9YknjE6nvyq9lvI1u3crF
0W+yeEftLT0FpXp1ahmc06cLPtHOa6Yug8B74CuABwJcSU/nvNsNS+ZU0CzHxL6pcm3N25HkqzG9
Z11nPdwxGyoZZQenA8mEAlXgshThoC2AHMSGkPisehuvz8YgIAHpg7Ro6W20Xcu2oaYOoduT7G5k
D0g4/mQl5MbGlCtc4MYEJzjwOFjhK98vL197vK02uCUoy/4HG29Ih5SKUfWtZ3jSpxCkRhyBkKQW
MVNlxoPDKmKfaibue8sWJlHhYB+jQBnMXI0AJJSYpSETeP920+k8S/rvBUBs0J6dCv8Ju9CR5iGn
On62HjUP3P5sehvgHSkrQ35W+Hg7KXQKwTnlHYn5uZdNAq7nYOuAascJLiHtI80z+7AIB1/xkenT
wIlqi05d3lBDifDh9B81V6GsPm1pb14jhL1xLQRajvS+TQDDYxgLDxrP8RdQN61cJ14lQUktI8aQ
0aLifMMISLwKJgB0mnv2Wo46uiPQmy+DM5okbwJjia8rz4/bOepWaxZgMN/7lZl4nEwEHgIRhYHx
aDNQPceW4hcq2aJQoVsHIkqV0jg/Fn3zpH5Okyz0yje1dfRKZFmELxYsbjDJAst2Dwm2PImTFo2W
UQbUymHGPpROlwwSIr/okFAYySDSHLM/yWgCfj9FsGYq4ssgF61HhjhUyjJiwP5wVTAm3NzKUj7o
RmzlYpi1MTESK+SGfNCXUQneRo6+SYhiMJvkqQIH+23SHWwFXKvrW3tNWEoxoAteT1KgB+V988Ye
3lfL4ScRJH+Bf1m/LvdR/b3dGARX+qwueCrDNtZD7dlcE3J1KzFBI0/tlOfAOOjvr9wAwxNCa0un
Kw3rRwgNMQyLzAxnotCqcvAOFHfXnKwE2Sb7AOhGM5CY+bfjkzLOJqnIRX+lVGqQYPxpQ9s+NaqZ
NZmQZwmwZJXLcHjng7H6KHQsvYTv+LegRtdJvVogG6ebEou99mG2/CQ9TNZQ1J5VLd0nIZ7gA6Cd
iVuTTkK+5sIbqbTBKjPWSwUvr1ff5hmJ/9hSkC75FlMAEWeEnPHhndIuBYgWqVZ2QCiwLEmJt7m5
DoT/azma8HSFqht6M1+fJZS+X2u7/8dpHCxa6vmwRbi4xATHyi4YluViHTdYYPTUeFuDRFA3A+H2
ag30L+M65BdC2RN9OTDxOqYYsolfI9TN0bqRsDiGgNMDW9YWbHF8PodBPHdrzvl4PIaI8zigjCG4
G1UDu1dYUh1pQiK2O47+VBO9o8tmI2VZo//b+NYbbSEG+SSzRdsnwRZq7vUtCiakLipkiOLk6CjJ
R5JOEL5c465IEG3rWpjvQHfwIYkzFCmCbWaRMZwkyOFkkmjbwr+S1RGo0sr2luVwoJPTm8qYiH27
nbIpg94Q9xz5R1kM32lLS1TZDQdDIuZ33jEMnFrV1zwX3SWApUnEZBUL/wQKLgqSGnz738XyrPP2
/g1zppnIBVIUwBrotSbb4acDQkh78XSnHpYuOCTuBxK3khatfdxiKLwOK1vBhfSXuga7EoxtClRG
a4ZOH5pQNxPPTh1TDA3gYBb9EySZLJwKUByF91uQNRs0uaEN2RbsjVOSe1n+iC7xRR59LscHTxUc
91w8ASp95tsBhFqtVce2vJwk4U0oi6OllnN5Xd1qxm1aJNtNwSi21z8C58gPdTQ6jwpm2sOpLIYg
uoxgbzPupljpzcuUitndoKNnt3LTGKxi6yPGuBXuZ43+vr2V1779Ysdhf9Q388N+rN9K/C8UG7Fr
hBbMpPLCMsK5hK0IIZqAbLlwgM0XdMOTPLwXvCj3aHivp+NgNhV5irHltDk/QV2kGxAjWVC58Rv/
4Xn7/NKG2tkPct4om8gUsCMlWQBvbp0S0AOfLIGyvukdNllhbjDpo0zVymCoIMzbDoPy8Gcjq0jm
jqJQWrhs1Ims2/e84r1pi07UhRPJUqxrNK0hyer0O4Mavn7xhOCEqD+tUjybHHZHaSZRFepk5q8/
yQT8l0xVYBOUYEqjiWZnU5qVlF71wBGlyXBXoBdESWjNvEB6Zmpd5046AhogQf3y8pKTapccstgs
UxgAQg+fXjdMxARNvlLOItAol3NviJoh7nNTm37vFi18eM/ZseNTI/vgjBlykQWc9tsM1ZpUkp9y
+Bcw50DoU9LIyysFuUAQu3jPh75cBBPLDrNmIXwuPyXEXlkvwn1/XyvgkcgIfFhC5OREXP+1/xK0
NuzbD5Tk014K/1FSn28D+BvrW0mJ4wc6Lufme5LKsgC5uAr+5qwGjUVXMdmKHmbWkI6KeZ67C0hR
YAyrkB8QHfAdm4+U9N9QHa5ZczQymVfKnXenj1GZoiDlm2xYUKIFn6KHXn5ShAZOsmggSpfWD87L
galbTZM92dWuqx/7KkIwrDV/jqH1JLOl4pc+bhCB8oz1ckJaaO9PVWiVyICrJQ/jfw/jLP9zPL1S
OMCx4bzXtfiVOjwi7jABZ7Khu7WNGiXk2qZA/tQtDXJiuRv+8PVBHlp5MQNoqFT5f2Pnu9I21yvS
hjupQG9UdjKzsjl5l5G9CZcWbpkv0sPlTUhcIfIKzbY1HhACzehh2Vw7Kd/q0cRcoPv6uz+l2xXk
9xgDVW2VR5D5U7HnNKMie+rXEXya3eArkkDUnLiQB/fmV3GjsPO4bvIqrobftNNWbAWKhzYuqPYj
ycGm7QtxGsVHaUBPynP4jc0XjN3wrb1TMcc6JW4w7Vi0A3OkgXDJPhnnrVuhLbOeFrpn0ZnEhTRl
gMb2owQOk6QU8WU0Afu2iYkNtbPY/46RWWNt/ILBWk2iNx9M+v0Wf5kk2n5hunxKfnxiSCWJF7B3
aQVP5VqcFyVhrDk8phXy2ptV92vHnutqjLuSgskzPTGZMkEoF+9kp2Tsma+W+Xnl27XU2eCBlCed
pE7OOrZdMcNOLFHl1COp6/f78wQB/A//pzMBCrl4k/YPWXFm5zzxOz3xK4AfFf6W0imBOXm0H33x
+k04LtyZgUcXDuA37mDXJ8P2IFbhwafnhpYkX45HBoKtdhOJ3kayG2GUEmLJyfr6wYFW+ru1c7fY
1fApLkEOSGK2RNGiuZq0QSlySLUbTm7Y0Y/I5esnQE8wMe4YJ4l1OrZ4uQc9zIaUgQLRCqUtYA1c
VbHkbXi6bd+b5uuDXXGyeLWCNrXGdZ5KWIJuhUnSMzGuPutJIok9X3PKT/0pVsqMFqTuv1w0oF9E
4EjFAGh63VUYrQs1i725VtxXVyznr9pdHSXAVm4cXDtMp7YUmXweohTcgPTY/yr3xQ/okKfk++qT
sdZ87E5DeC2al+7620AmIsL7JeN4dUBSUK1zKF/etU/RfTHILa9LYzQrPPfM2zwzSpEfOCBauoso
OUWrpdtOHsdyeyg8DO2h5DvDLruxHbUX5KXiu7GrPtjlECAbTyK5M8O7MKEpRtd3wbzD2RXC39Z1
nlH10ABuakQbI5+Us1JWXw9Tw8NIHSYm1Bf0pb6v4o+DJFOsh7fX55Zw7eRqd0WMBA5gKnNgF8Cj
i/8X3oKsRDWH7fC9wZQXgo3pOUvneW5kMpbKvdVGBug/a+CEQ22zKISdXihBnGGpgWqu1qG/5wYa
eBVH9ZjxiUUjwvzj99K9pdaHhaDCTdKonO69j+ny43BMyN5oqDvm3mJhjRnOIOYo/t5ss1xiVShU
odxDtHimfh3tDTHqmxtrWEjn+xCvPO3rf3FdreNQs9ifXappWP45KejTRFqR6/+9SL9Jsl9KKCaU
xoN5C0WnVQWDggtEbx/fSAWDD63E1CCtf90+aiCTDlz4Pacur2JFWSXm9+7OaBADK3mMPlkW2joR
FwucXxRMAOTb6e1HV94JkggaoC4AvQli0srx1QycUsMnSWK+j9UAmaQ295nOHOsQ4XHwIiOEIDPu
eTzV/Q1/NKx29F5VpkIybN2m2OTVnnNt4lXA9frh1zht0CBhiEgjbuooahYADtuPR3zVavlzjM3g
68EG5APs4fX7/YfcNO9x5ZCMz5gei0AWL03k0WyTtQnhtQfjSyS1pD2RihA/LL/xcsov2MFyZPvX
xSQCtmbMA9hgRKSG1kpm9sJayljHpJ4Se5K0imwLJTYXTKgq3S+ISobJKo/9/l9Q4nEfYdchsqMO
DN1YVgA/2sUSUxas+4+OSpls+sVH/8y5+BCkPlhrhORfrGUlULKCTDdlXH9dxHFTCapSArkti/f7
5U04cofqCHFpjk6zBK+tX7Ddw9ITKvHZW3HAhGxyNQ6ckDwYwjtFqXrcTKVDLGZ/RMcwi0czlzYK
T4a4XhJMZzAtcCxdk0hxI6V8HFkoSVTL8fCsFUy6K6OaKKmn8AGQYGoEEPmyUqOcqph6Fli9gc0p
lJlv1KH7uAlu1ipp3z9fv+FnmDpt3C+Rosc2Jyv44GBJuix3p3l3NbsXtVDKYiGvfUgsnaB3QHCZ
d0tg0td0ETK2wNZuxOm618nVKbqopmx6t48bd5Lg1DmJKE3RnQiVYm+tmjsWHuWbQFzm5fqe5Dqw
YSwik3UFPEcDefuJGdYV5rmMXYU/DI1qd/r7LAc3hY9Mj992Anz/RgLWzPdiEe9OzdZV14dK13R3
WA7QGURaQZIbBH9Li7bkSMaDLN/0r6P0egVrVGAK9+m8nD9tPqnUw8xcG4H4xHkiSIs8jCEqxMZ0
efGLJfQ15oQlMmk3X4KGAAMTR6UF6RsPNBa02dH7lYXXXZzZaWGPUieCL5Wd6L7NsnnafTyIaIgD
XmYbUz+8dTzBZlSddMNpJOgW2b2NRaFvwtZO8SsH/4uyAwgdSo7oFGno9RDqK32bpMJ8V0ZdYqXZ
gnzqJ1dXoJbD5xuxeKbyHzDH8h1KiPIUvt4UUvUum4Gbyf33QHtCdbjXDOBW0VwK7zAZYMxvIzp3
y/d2S273tVooKOx4faVNEoRWOPmdrDvrh5F1hSLclQ2+F/6hASD9PQ9wic2St7d64nPfrafkRBZp
q8jHOJVlnkJXtfrF5CorbVz1oN08fqQeWJJHILpVKbDzltZOu8CKg+WkIpSNKQl3EXYqPUCuL6xC
hXke8udHwAkjBv01BikV1xIzvFEOSI4nchOEIUfbbmPg5tnJmLNL6HOgfW7/qBTNz9PjUZWfa8JW
xP2mY4b5qYg8RYQY8BWc/eYpLTeCx0KpWPqWnOm7JglVOFp04jji/1YP/UhKCJ/MZWTFtZbnW3Sc
IuwqTknwPKF46o0c4Z/cUlVrjK09I7mChYZUvQJe/GnjyXLPOvnCh247FYcKryZFd7wWtyWQa+Qh
f35niJo6NKRarCYPgsK1rIBCw7rP01lpR5AnHWaD3XRAmBszKIjFXhmzRAGalYD0wDPXXrmbVnmd
KP90AZ/8An3Q+CDvxMNJWSGW1Ab/Q6R043Fr1JKLl9Pfsx+f5MhTkN3lVvBjQzaABM1HRICbzCbS
ka8DiCE9R/foBSLZfnb0CBDnah+fGUzjI8pTCIlxCe4oVylHgAqkBDd+vytZkfXFUCC+40/Y+LRU
GALSHv/5naleuxHCbZ8tlmcR7AXoeYCwS6aD4dgDEdl/8h7Ht2avRvySZOKm6W/tbCC2ykVQOW0+
7sJLBlwTB2BtoD205VMNRJ7xk/qJnQSpHSziC1iampI55AvhNibst6MRFZ9HSFPv/niqAasX80y4
rWYX/p3ftEc7ZKUIxFU7mdtobf76RzYDEztCBTeD6YrDloJI325gai2GxMRW79G1Kl8Zl6iJmW45
k/MDvo+qxpCrDHrV87orL5Q7JPRLftqN8O9+jkLJ1bHOfgJlCxQYPa5CqhA7gYM6hHuLMPWacW4r
lGndoFnYe7rbi8+0KX288K7wE4hQqeQYDPM5dYwhKSbo3/NPSiS/7adaLhDs64362YVVgLosSFmT
KkO+Pbbx/FOFMTq1tBcgFHIlsm6mLPrsovTyCuXQcPECmODafwwPkYUGjxb81VoUuxliefJsKw+I
m0D+J1QGPr5ytQSH18PPjXspedV76lFCFso/Wc9HDgZxmju+IjabevHEuIWcx/WfAUdw/wPj3HSU
yrvRawOICUCWi444YMGf8Eoxf8uP7tFnxSsFP5L+RiZy83FJFwnDtfzAW6gMl6IB1moe8Me4YAuZ
zSz1SB8qDCkF+2wHBSxxL6VEx+OaD0mkactFFMmnWC8o2cJ/WYROxoMKlR0qps31dlE9fFKvPA/t
3cMQjkhPDAi6RbbaMOshcTGm9jfVaZxxe2FYT0sXVMKda8CZviLWkOR8qbtpq6sdVGil9Hr37lsF
hzGiC00U+7f43hHX/7+znUzXRCCQak6iI/RzAL32kf8uT2sIN1ehG9kx77NUeG/MPCUXxysjHdN/
4Nj1MjAosZytOwMdTcr0U2SHpUoGWsi+UjtJ8ST0pMYO1kClPkaJQ8ISgZcEHTa94NiBr5yQhvmx
tlqUWDIuZJX0HNoAS7UzlxXP9YMvNfigDtBnXHr57Xgls2GnD034dDBRgZ9COp9kun+O9sYZECo8
tzRxTx9CkBX30VLkTxs2m013W2K+O53anwP8QrxMdI+VaZjgvBAaHdmmH9cUO3dT1+7qoWpqFcJd
ttf/BOxZ/8Ht6uycP2iWRLX9EUQsGfG6kjvsEhG5dImqH9Mfa6rEu055VFPcLcacZBZ26+oMwnjS
dixt2+MEizpQDQy7U3uBmiHR8kpcizibxnQ8cX+u6c7jrmTV7mdEphumSZcVhEMkNthzzH0De1c4
6BOfm+JN2NDKcwKfhDNgFEu2K1yKHNSWM9TmwpYWdcjNySc9NLUgpV06eKZsWjJ7UBOAnP2GKMv0
5X9SYGbHJxTm9nfH//9N0KEKPnkuBDeznUaXtmmUGYeM2dPrYWXkvO6MPlImmBtkLh3/zEnOU/WH
0qlZtD8DPG103niG1l1QgLFU2QDLYhGuOZlhB6ajq2l6hayrDhzD5jv78SUBO0PjcA/FF/YqTokM
1xIy0/e7HECdvztpwKiGaT+gn2uztjjzTJFjryxGy7K41WFUE6SKglkhiovZXF/D3cUsjNWEoeUf
Xn2YOLaujy4hTAXGdl5FWTmlrBdz5kkOOyiVaSqHSO6K98583Ef0tfObS+QpIIxs04W5Q6PHeFcl
OTrmoyOKDEt4JKWZJ4d9bBDPQGQFwilG5xvPN1EyKQ1QSjakwogVZONQam23mfynWEwIjt0Qncvn
qiWu9b++tMtI526ZVwU0pTEM1M6ze1R5XB6kpfHGmZs5AMU2NTwLd/rms9JX+8FN0VXcRnmvXkdo
3xi7NNVj2N7qAzLvN+fLKrYPhuFX9BApzO6iKHcEa46ntiS9tnYupOgw0e62avBtyNStcIfBPWga
ghUMrdu6peYT1y1+3yCnQhkwrDCXmD3ZF/kVNjsYYv1/XSXfHmLsbd+uBMyJTUfAeL9wSly5fVyY
VcqpEpcv/NiZem7LVUflmweuUvpf+szEQrpdD+RDu851/4aiqwo6njs5JvQoSlHTSpbtxsgGoKm7
d5PkhvgWozD7h+op6sTFy/Y7t7MKEXNb3h5qsdRE/1OW7cT4x/qKmwXyV5UWa88e7jtO9LByUqRG
3tkm4+nmMrT3vCxUTQaY1k8687Ti2OWvUzH19zoFOoFSLq2jCjhE1gvTlULRBXiwP/vRN6ETww1h
B98Mih+Q5eQoqjgjY7dLmFSOuBCUMYD7pSw6HXHS4eBPuCkQAnl7x14tYG21HaZHOVIi+kY3LmLv
LDqdhlvjyOvoJ7xpWKYFdDJZ0pLvTnjlw+pVLyd+xEZ7dpjF93RisIVLj53OnJd8YYgc2tHIexWk
u9ypslt9kZWaOo8nAsaL7sE7UXBNn3frgcypmyResq7JfS4MpEYq6NL+0ySvJWKNpktCZmWm5AtX
KmFL0wTmAVZ7Xp6NCZEc5YM3QSliWcr5J4n5G8sP3bCRejqyXPLGEowcys1NdQoQhvCV7KbZwsZO
6r0Ujwb19b7QB9AqPQ5xN6tF3R3iWhuk+ulKSeQpgw0qVH5zHg2fKnW0ViUuyj9ES9cpZ2dbjEGa
YWli5zBYrfsIflUSklZ2+NQ4b3WDEjx8mw1Y+K13UzWnkV5vDExfuvoN4nLwA5nLAgtUA1JlZVxb
4DyhwETfShli4EUyxK6ZOH9GFj+yUsnrx08uLEJITwmHKtSRAcxMRbcm679EB34oFTkCdDMmz8XW
ed1+ClVoITJAKJ4YtxtC6+mIuiv9Jw3UzTO55KnJoFQANgH+ndNAo/QOztZ+SYE4sS8kAibgnXIK
SqcyNx37Lf2O65DxsBvk3ot46QehcdsbclY3Lx73civ+TOvPgkTV/SEIQ8VTY/l4772G0+4kpvTV
RnClHXTY1MhuHHTAFQ73Oj0gnR2ZceJ95cdMz4tFQqS6k0YGawtpizQ3hC69Ax+r4wUGa+jnNABN
MEUpZdrgUM2EL5cmjUX3xIGOpwrjqlFvJiAN3hV+OYmEyFCEJ64HjOdMI9TAuZLo9rnJsD8wda/X
lAoGLxt4KbP36Yo9VxEhbPBd5Sls7IzgpA805f9EZecA6xgjK4gXDPHfXoSSh7vztBPyYZa4Qu/+
2k5y8+NFUO2gFDV9oR3nUSbr5zNqoEjviTEGU7rct3Bq1F/jx2UZW2LCKnfpJja8sypbeDZPQ9Bw
kpi8VoGShq/HVrm3wf9ETeGZzTIcmYwC11X8AB+mpZx3hqhQQ6ZTgoCAKBWd1JTNW4vM2gZ7mO0v
YIMsuAK0Xd/F/ZVQc4Tl3Tkg00b4QWkOsio945mtgWnAmQZCtp6llrq/numsUfKhQYAuKGJ6qpO2
Ft8LpeYLryDO1awztVB+awgJJfleVADlR48MJghE/PCOwduy3LmBOPYG/XZvyGeY0+CguW6XQ5Ps
mr2fgoY63ub41DWkodrQVPDM5Cx8BZ3SfDs7SsqGKJLa/diKSMC2CVn4rlAEmEscRhK4W28LLtQ1
m1tTq9TMsYklY6IWvOkXfA3mWHeAVL+bJ6i9mbmKoInWsnbCExH8++IMC1vxHV5ziMlMFLj77mGL
PD+oP3ZhPs/K+VdgdQPt5b7c+7V/885yaZFD+QmbrtXK4FhK1u7XMztRzszjR+9EQ5qck04FI4fl
iX/Ai3pJGEpzWflzPrvXOqePK17uQQyGoVNzBaBV9ogt4p4Hn4DeqW0hCkuVE0J+Xzwg3Z2KdJc1
J70bcrFOmb1BaQ/3WIl2m29AX4S0m0Cd2ccQ3jkWggPoTHfQUfMNdw2OvVHV+Az2nU36uK2JBlUg
M6HNVxVTPtAU9INaGFfKLu0Gt9WaiRebJr/TJ73VGlk3/MpdONC2uKzUvmlK9ygfqdnVORS+H1y3
qlIIwEUJOADFZRmjhGJTwdFlBj8twJIsqEEQ4oO7kI8Cf3rGe2PD/leYmh5w+kbAxCkTvHQoyxwA
gad0/VQk4fGEYR6idFRopqrGqg5RPsK3NLF71mfQS2p/sSX7UmIOHF8zH1qi33auxQu5gYMAmXEf
PgwKEdR3LSwu0DavcWeqSqsYl6pOR5fr9VfrF6KyALLoXA+DTLis3pD887lKVTu81XBw5JF5JKaE
9orjZkoRXrYV4Bx7KMxJ6rE4NqqaEs0pSVfS1wNY7eqFqGanXCwivHhYFQX0WMLLP91cSGV6xyiU
E4iwN43ZmMRCmkRmxXEZyBuz4B0WDskohsd1B3PHDT2tFXhiHuYLB3MDC5czYIqlWubaMmP/n1+0
3asK0BgaTTrkWF+zHIuplALQUu901MeM3AF0JAKzoiTCs9UaYdIVAXfw7QF+5sxTDlyCgjprxbTs
jsKXDVR9G41a0VzQR8ebF76UjYIoiWrKHpPnLasJ5A5fmRe0wzheogCULwfLIL/ofoWzVOalUAZ6
kNbl5mm1PnSdhtWwgP83nsmySshBFcklGnvmAqooaiM64+Wxwtj/eSdLF7Ib5UlfCr8bt6HlT8LT
BcYHk/0XpetXp7FzSi35vTjUS6TDUHxTDhb/bM/UTZJK0T2M3cWhrySqxHnKUX6aepDIZnnAThC6
2QMPkExSyM8n4LxUK/10hi0sueNs2GKNEcPDuHqe+0ndZXBjwLeXsXXtBaC7IqiRYmDYYzAA184/
sjPY4G9T6quxPif/LC6IKPtKnllZSyqdWoJCCRor5Q4/mM2Yr9a5Mvvs0TyXYJL/EkNK8WGqwJcW
HbOSRQ0yl5KjgBiyepEdbn/vfsCbDuo7H4AKJ6M8bGJaXdtHo0+RCN7swjxevA6MlhZaN9MiSzQV
Z+CH7/px3PSGnaXCpQeDjm8NuLofwFdvpSU35bN6iL6KdCARnujZm8/sTurxECLG912eYgF1qEUr
ItWOK/HAP2vbCrTf3cnAbqi3Kmj2Du51Urla+V3E22evj4/8rZLeoTzMV3brS3bOZa+2CBadM7D0
XKXCNV7thwg3yoZevdLcpE/ibTQ6UAuDtVI2AEEpICvM7987CfPYfE4KiVxICHWybMAI12Xn8ZJz
Wde9VpLR+VEzqVfwJW/PdEmApb3hzt/CEFl98PCVNPIQVwAEaSaPAZ1ym0lM3p5A74Wye0OSKpmR
zOyrPixkLWvvb9ZXDKSFzZqkB9s+cIGggqFDS9QELhKeVtoe4BGFNEbgmYR2CzBvat/i9nVujAyx
gTmG4kR21arosKZviNBfbO6t39IP7gyN6GOFZ67Vvrl4GUtURs1ylfuY7TjM7ZketUa2U7aPKoMg
fKkzBd197EjcbeCuI00NApXIMvAeOCror3B09AIRkLLf1o7uTjlAJrqPPqsl2KTxse5rNyBJvylC
P5VtFMjrvl7v75MESsAoE0t6DcrnVOgBfCTuKmqjrUnIBj72dyKzE1jVr02RRmTrJSGrimHJOnPI
Ds7h1OZIbVuyrnIS/tG1X50qEiGq+CKgNSOZqonZ+w8FHu0dm8ts2djtRPNviNfQG5F9/fz6wvbn
FQw2svE5S+0cklPAK7cWEEshQDkBkHtQi90+FCiFF5KRz7YSRw0bGwLG/iU/oC9n/h08vStBFkcA
5NCgoDiVMEDHA4yVKjOZiyz1XaMDsp/5l9lC0pShserhwfQS57kE91c5DaBVkyd1eimskX7IyDqo
EGpgvO4Atwnmr7ZwGWMonbCL/jsqm3bT1/hVdsyF9c4tHX8fEhFCaFQfzNF1Jtj+QST3X/RDQe+e
gmy0u2NAjDHRde0Q0v0eKA1sCEWDqECOVu4b5P5vzXxSAta7sQtTYT1HeQpTqQMFbNqDxvFfFkbk
DoQ/eem63tdzSoLcSoZSTKqIF1EQc92i/7oH1t+4ovzJPkrOgK2ISm8/Q1sDMveiKWXJ1e4kdsfM
0W+Cifx27D55AzfsRW1f4YXJWLVzmHEKHVzabls9RhlwgaobYU8Oq/wkFmRVTm45YU/FmBh/eyyi
7NHrurm8daJh9m+Nvk7SuBZUOKypGa77Ep8mWFMW26CnG/bd6e66JkTMYv3MbxRq29xf8sCtXh/i
Imjkrl8uwXMS148W8S/QjTm0Oy/RBHZCWqDE6I7MEvHgV9ukeGJ9xdCrqtSIH6lKahEiRH7pM3cZ
oEC/puqDC9qM6Y+xufjhk6xfHroIsKc8Kn1vyGGDzlWGsVptaJ8D5JR/BU5o0WxEVeeEfqrFSIKD
gChKBMyL6easep71T0ABkghPUC01odAyMbFSMPA6NeKHktwV2o5AgMmCD4LoYfPiVIP0avePXlGi
D5aolJ/MYuxVuAqMyaBZhFc7MXc2pP96+HB6d6ZyYui8ZRu8xzqhIbbhiLHN4GbKlbwPfSTfHbad
OKSolF9kLTOfKLf5y3zHcFqIdTbOvTO/lG5LFdDetrA8ffAia4JRw9+pEzxaUlECRKcN36LR/CfA
7eQsbGcrkLv9i/1NvRD+E4ylrtU2JD5PFhDBRJ0chmjWsHThvwsT4vpYF3pjTUD1+n1hpOP0FL5R
AABLwFAjEuUg1dghfRYaoI74R0euXgWcmZA3wxFlbo3XxYwe/kRrbxT1hwQHgzmZQpUEyKuVSkAB
4xlArphHn6WaVQjDAc5dPntssmpgyLse02Szuu2bLM5qbig7a0kzzQ4aBzVfTMZzUw2AS862wZHr
/8rUbQiodH/TIxoUN7zUnAscB5OZNJS4cYC7fBXbbKyIn8Wt+rh9DGpLmTxdv+hq4UPtkGfSVFBy
oZUc7MhSGGjZfkfJuJmP8AnirquPek+AtovZM/sMEP2P5JOpMMKAbND8/s2XeXC/Dra7j3lSaE2i
dgGWGXDUH2Ar9N77LVoUadMHyor9brX1Q/wUwKoIMRvgbEn9oZw4dO57qbxdkfx6SJQFwUMup+Tt
Rc7OIN4dXBStxXRyZ5eXJ+XZRHn686rN0cQN0eN9ZZfLasQLkeit0qPFA1dZjheNTk9Aykyibqwj
7BpuEhdtDb2gSyo86Gljkmmzp7nBNN/gIUTrYM+zry+Zi2873UMxM9A5+4tANroEkpS0wr/VQWQO
iu/Ek7b46IM15WRFiqkoJweVSbukA580f9sMcbT6rxgqIyDz1JA99FU67sxLMZmY1cEOBBGK8jY9
UhsX0kFvNgh9vpQa2qiCXkOAa8ZsdXdeHuwyoHqeD2Y7nlwlFPEZWUO+peqpK4U2JeBbiTXMklVt
7FIChtbSnBjtYWM9xHB7sB9m7uShbVaeRfSZJJkb0/S0+/wIqlECfey37CC8xsytaSHU4xaQInnt
v3d4WjAvJictl2dvWbecgsTYWBFwgUJtC0/6k1aXNm5C6mWToq2LsGZMjb8FIlr3KHWQoT+QJZb8
6NYke6zxz/AAOymjXkSc2q+dyC3H5j6j8QLVHG8AqTHhHFVaRKf2Xaz6OQx+15iaW7WaXU9/KLfi
+wXm5+ZQXW9ORW1QlwRn989oyhE9YfaEqh/YHMUwDDC9FGm2LPSPRijxS+U2ybpQkVGx6Ys+0XRb
6ZM9E8DNsQLEhEHBAIis+1mJn5tNYG8qz0PcBQ3297/oqqXqRHc/bSYtv7Wj98r0XLEXyy9OoFwv
6XiWylDRHH8T1TXkzxW500diVumMfxvy+6rWHkoLSnHCAqrgZe1yJEiTcDNucQbK2a/QF55LibPh
vkHBj/KgMyIl7DVODfEl5RkHGKAO2sKe8wi2Cp5r1w3uwcb47IS0rML6NKJkZ9RhdoGjnLNZrDPX
NU+DUeoy7YynZEO5QF5CJPu2hrfd1C0jRbhB34cFoWCDGIxoJwjy42IBtr8XueA9n5xu/nEODkr/
7FCOWB1/4jCfVEwU+jvPhm38FoiVV5aI+Cg8vMbtf2V/vFUDSL8+51jZ3Xld6gn0cZ9eaZN1V5+6
BIXspj6P4NURhTwr7YJaKLUpsWaRS3/apHRYLoPHfa8eCASnziK+FGKyr3Rys7r6ExBJOXcmZf5m
JZ/LbHJ9nH/Fw6OX99+QaIo4TIzjRtxUoNW0nhQb9T0AcS1Bv/RYi8vznyecckMRfLUmU5gQX6TZ
flbrBnq3hcZTOveqj+JV0ji25yJH+CFEtLGjb/RMKco2ugEQk+Oqn33NaV6Vk78fwyciURW7Suv2
PSISIJCL6z4mcGv8Rk85u2wyQzTk+Z20X6u8D8MQsrHtgrj79kVCPLbdHzdk2PN0J0Ip8YkBbTOj
Du+6QxUfgCPlyKcU8tZtTO7qb7/aa7kWEaj1wxBCRyJKtKeuCIQf96FJjsesf7cDzRwInDwtPzaU
mFZoXnhTHUzcMxi59B6YjWfMfTuxZWe2eFEW5m6RIJj9UQxVf9zWMgaql+FF835bZYaJYgsp/t0H
O1RGYNALk0d9W2hjmpif2QnFjmCXMp4qKF4LKZLkr01SUlfuT9o73OHig3FrJPS9t+PyFMeAjV+V
I63+ZmgiF1qajn0zdbEuy6OA8OnIb60wROcQH44D3ks03jtqS46vY9q6XZy+RVs2CUUfFwhIyq/X
POk4t5grL36Q8X5A46W/941Xtwfr4sbJDtsO1MleixiyF610gpEW/t3L6dmmt5zg0WGq2BoXgCNb
f9Jbh2p27sgOrxK7oJL7hFHOShO8RWoNd6L+3IDJRYKUZeKYeQbp2Bbg8+45HiLnwE+ScieAExPW
L+pwUS1N0uJYDcmzmX5dI7zp/+w5wHE2CqhfZ41Bn/hB64KvNXBS8fhcYi0AGkewjPQUCXlJWmB4
FH1kTnMCsSibLoY+APqTLCRtGS01OCW42FhOl/HOualVaVBGq8R1uwQYKxY/vWQ+TNOlUnhcCnmK
5O7Lr4JUUOiKr5P5YpSD8m1eKqX0ZRswx6Frfuea0EQFYQqqnA3lbRUJEpCc1udhJoL3ckaHw7r/
2qcgXhnNZ5F7P00qxzfhiBToBWECUooHxvPo44KIrJEBldxd6r79c9dusDcR6R1wq7QsvIcpm+d8
O4X2x1IS3Nx3B776gvx3JFiXvZM7S/OekaVv6FD9r/mZIA8X7ATv/NjWCRqWj69Xp+iPSmcPndQs
tuTKZbimlohBh2aW14F5FYSfoGsdK6zuQ/KUnUSTMuzEzgD4nf6NcJzT4dz8abXDidZjyVCp4NvX
9CCzexFsxEukvFVJm95S6KENqqkiTZ7rY2gy7Sl7B4Vyjr3L/P+FTZGOzQ64b4hNbsiKdEeVQj66
q0UuVIlZ6nGke+RHZXoe3oIYTPleTboa3QBTmnww0Z2Butr9flbskwBHGKL+aPtHoQRlQb/jzv9i
17YSajW5mHvA8G7VvdPzHleOgcYqewftIfyB0vhrfJHoMb33/E+nJwsUhkhamb3wjzsJzVADQSMw
AuqFi0cKI9QMg4vWzbBt2kIyytlV2XqfRiRKnPjz+NoLUPJuSEb/pgAFgUtkbTLC6tig5S/RzBKh
wPB52/O+IPFRwQh34WyfGLSeEwcdZ8R9xLKoC+WJJO1l1SUmlnrjuAYMBKjN78aJQciYiUNytmr4
PrR1yULpzGW4nVdK3rOzZEWn2m/YJkeitKVQhI7k+sXKdKE7cDoAfzQZCchbuS7MQtXc2nyJoY4k
qcAd+e1FawwJ4Q1F17QcjbOSf72IM0AljcE2NyGvnDDeCdMRBHT0VaW92+aNKqno+ZQdjbM7k5cz
B/iLTrwcfmMs7eRmOYzNz2WIFIrk0gYtB9gRJwBaZZkv7WjsYEIIWhd+xkhrWYQNq2GuJQdZAqLo
qMXTmils7ueLK23ZA7kgY/exr5RUw861itVb6xHBQzVNwvTnrBeohWU2+axrx0xCkK2SURqOWzly
idAnHHeex6ZtKwizulhnJq4jpCU7IXuiHkFSclKvkGsDMi+g3qUAuX6Q+pLs1nfe/4YVRcnWlJ+e
HgGZxEXX3pxhgguZFQRfsJ3y39Bsyx/NKg91HYagrw9jsesF1IcCTC9JIxv9V8FhkWphV6urD5eh
1T8KruXSimcwq7TRRlojBfShoQTIve3ZQ6pT4BVg3wS2eqDajT1aAWe5ssDb/xPkz9rGrWpvhzsu
NEsb8uKGUvjQqoj0gR8ahy4LjTc5SDrpKdDKyyqRZzTplPejH0JyQhrOFZymN496THWyIcKUlrJB
svAb/0SazjUWwEJPYtxp9FXJgR3PJgiQqoc/p3e+IHBaChzMwPvIxeDDSFmclHJJ6uWos8ha/IMB
O3qPS14CzThUDWPo+G2FivxJDrds2aHVPvTmiy8sBxLqb+VO9UFGTluew+bRoFEK17iXmAI97MgZ
lYjdcJ+sNjVBlV52OuFoDnlQVCNxlQHSYOBeDl9WlmwjclWbicJqqYs60y1N7uhbTWG6Jaja+jwt
8rVxLNDIkG51f7yEsNtxLuUKHUn06xdj6+3eazXvrkYWGFQMBbjq2zLrypokIo2DbdISrGKD7lBN
JeTA1DIatt5rieZzeZvoYpZBYSdRTolKvxXB19yHBMBO9RwH6u16mGk/AWubeb4cOKiEaLhDaCnf
WUBb98VMlvM1NozygsoOrseCYtS/9dE1kKaXYzqQtUnO5aQtsW9pR0RZYZ2ISukyQ5aOjMlIT4dz
oTMpknwuksZTEvPFZuvz84kOUCJQUPc/gz8exhYMueOimOS4M43kmhDA1KVBfypqf8CeHFAIO3gU
3VTIml7hKlAkTQtJ7uR5u4p0JTZkWqSnHwJjRKhzbCt5sqiwVyWXnAAopzkxKU5tzwoBrCJ4sfhi
D2S/7fyJx3+xzTLq1nh7ECCEasU4+CeLyfpBHh1Jj3eULYxBkdDb0P3W486RAh3e4D9AQxUzjjg1
e+TSO6ZCO7NKPO9/acTOCnqOzlWB5icX/wLT07Fd2hRxMdMOi2vOXNgxOnHnzVlhLsMoEXUJbMxM
fsfmXPtevhdy3OPcjs6/aakKB/vjHYyPzQGgZdIWR6M7ImKQjjZD/x4H963i/KB8wodaqmZGR/y6
ip4flJDHLsx5Oec9S00WMLeBxpMsb9DLSDE6phUeP50FDq6xkLESK/xLmN+Yg/4phohFnl3l6pJ3
1fS5hLB2lUERqg5QENU9Z8XFjbtsmM9lU7oZL4l+hG8xKI0ZjDcWbKATy15N8VfvSwyBkOXR1mlZ
0p7DqaugkY9T+UML4Ncwvop6czxszD7/e0ltUXM1PIYd72XS5ITWugheWodOOxfWSjlmAE4FPy7Y
WyQimIeYXGf3pAyYub1CLYxJ/cXR/wh/Zgsowpb89xRQXVP3z/y/+c2Gbd/OnMn782LTK2IzA/f8
HUyzTQScsHJi4lC/5EEfPFYlAXFDh4HdkmdvuxWIa8KnQ0i8I4nHyoeTkHejsqxVlVPRaxEZAIQ3
ecaN3Cn5faGo5tNn0trVVWSdYwtZPOUTzVlxBB0AjmTIU46JJzjP6V4960W5Pbbca8bEY0eHVJZS
06H2Ragey6xYfxjPjvkCxN4f7ASs0M+a2G+GahoZrS6CNtGMxtD6pBVynUlE73se+SMNCpVchO7A
uay38CQWUFm89kVc8qih3KZ3kXstTx2Tp9ao6fsIvkIeSLYlj1+aC2xAp5poZU5zSM+MJUrD9oOp
1j1ZIRvM6Al8JO19U/nlvztItLV3mDYa1Ui5N7ohbNJoZGfu+NTuMm90WsiZx2USs/JCJ3acNEJs
AbF22cUoHzzrLAr+ACQ6eSo8kw2tqOl4pQ5Jnf4MVRjmnWzRQg+jQlVLi9xyf271JCkYZKzRiugK
qX1fOTQfg1TX2j0j4S6HPKazNJXKypNlza2oVPZmPg2Hl+AUF4IK9KI9ZFAeg6Y2lJdrWtMpY/Eq
+I+cqffPUbkThYxOO7zsRwFuggy2Q02XtpbIpEQlWcTNufbPyqslqRy4XCDwJ0pevnKGTxjizi1j
5UJwQ6UA7A5GGv535a6WiUIbI6QrEvyGMvtHjh5fjQhu4nbohW6GV9+yYegIudi3TVMOoIWTeoOp
QeB1MHh1a01ELd9HZdBryO5Id/aF80ht6swlDHoWNeL/PKjrujmEepAkd+LuBOYTQPcvfCT2ZCKs
3GriTy2d5tJFkJgqmiGtj8KePl1SjebgY3nQ2bvhOz0eQudV0Xfl58+AXOdqLC66mapz13B1EyDb
MylXkUzfZeXnPzRz/PKPT0naz7zIKfMcWr89z/WWTq+zeRzpT3n71Iw0tqe1Zajnysq+Kq1y+bzI
s6upoyMYDG/LGoxK3ZUG/109YKq8PcNpMnfQte8g7S5GX18TipoSQrbVQwHc+mtd4LDqbjcMzvG+
h1pD9TfaACTk825XYutR1qNpu+nSl8ZOyLclG+NscfrQ3Nky266Jv56aGRk6urizRulmTjC/C2ZR
foZOEW3jY2J23zamGgKOJ1X8vESLpkpqaPK0Q5T6D5L7uFS5+zLMkuYLWHJoAcl2g7vCoNez3kbp
wPO/AEf4IgVn/eYVi8c9mvVK2d49IOtgPECJ1GUQMWV9eY/zvj1QPRMThEshpATLYLTR2gfEmkpA
MA7wTGYKtXheN/YASZTGgP7KIZrqIOq89IJyzJhEktrWjj6Epp4yUmhzqsIpKB4YqO4UbL6UFIXZ
FGJ01tjV/6csk59LFjjKArQ8G+ABlxGyao9Co/JqrSrTbmAKOo5BWwuZIUjM6YhqRXbqS25quWAS
N22DAKQnltHKAF+v0b38IBDj93bwHHuf/Kt2+AzQqPzb2tMf9T1yE+bTobnLAx8XjIp5jQlkMZfl
xc0GQuY6s3B21OmE2ADsfWKLAFngNNz9px8rWW2UhxQepxhpfAmMbeCeGxt69JewdqP10YKyUoVd
OCAPfEX1qBTtM9JSTqIG1XumShw2m1ibR6V8PdjSDDjNyjqcNX0aatRlFORau+IYMLd0j1sLr4qz
lejw6dW4x/k4ck+51jdhYzgJj7FO42f8UnLv3Ww5BzwufIgGiJ98Jqfz52IY35kQoL2thkMU4c4O
ms0u1FnTb0LmFC3oPZWVg8xkDbMMEW4lXmbtfpBV3K4e3axjGv287AF8pryPspQWZhWFxDg/a2NM
nXH3+TJmzEYjWhiyyzj/y0uLsKJHvMIVSjUipaNYsO8bwn8R8IKI8dYrQyAux9BgkKWByKDVU5p+
85RKZTmcjePydV15cK/+i0rNCEa0Vg4MgYUjUragOlDEqD0e4XTlkpFybCxmZtyOCNn16lEsH6+x
0qAP2kd1x0IAvYi8UgRVE/FHG4vW//byTprmGhdwub5VjlqEvxIWD5m0bn6EEHwEDQ5P753AWmo4
jLGKPzwdvI42zLccFT2FUqKBZKm8mR9OZtAAKY2ioghtHLAhQVOjI9FoHct5COgyMQtC9OWwQsSH
N4VCddjNVuE20x36LNG78KdEQstzKv9m0PyX2mALGR7Hy30dzyQIjNMs6QvBtxFemRBqcowUxUvO
vkvIa7tyj2YOAf71JPvSXR37w6cXZdWzetmH/o9fU5JLO0b+m7nobucRlkVc07uLG6TGdIWAv2do
jvSTRjZRs+x+62L6+eij1ZpCzYN+syNikQ5RZmdkv5zBG9KoDEaJw/ulqs8DRbZWgyLtjV9aLii2
EuUse0VbjXMmSWDy5YLDf2u9m3X0ZIVevmZMvooKZ6BjHscIkdH0dQRyqzkZ8YreldfF5KA/xlFL
YF2VtcTW/NYXLsaHSSnvKO1b5cLbDCobqK3wAK7APV3z0jtLZYTj0rERK9gDgzsh/6QvzTf0Vz1h
RyD8vNnkfN/cRrAQ9D0MIr4tuMSWV1POBupM7aTCjpZJKXkrPDoFPF2qWcj8xg4FNLhtwV3y9JXl
hJzp18/KjAukqmc7pWhHStdUjiMK6TQwvaaK1oh3X6wdxwzXjI2Ku7fFh2m+E/NcGLNIGaKhMeNx
JTZW6Ji+dSMvWv+oVOIffXUXp/SfXotwWB9w5ritkHVnmQev3oZs7WdR5L31Ou33TiuPyQsR5gQT
t66AIOfRjwRdRh4UfJe4BnckquCb5nTFaIBIueL0p/s+VR5LVi2tVqGHJncAdAAIbfVx1qtPpt5d
x27f0PXQV8M8gGVRY9CMNQszEoMoNxkEWUVcAbOnpQEp4on/MuGqe+3xT4knuMK9wy5RJcvkZja+
C4NSsr4GyCAtOEAe4376dIUw6Bw4F8kGqlCkvIm1ozYw+ZIpxJHeV06CWsIIRD/qpA7xEu7M/Jhj
rivOeFOdUnhnr14o2rvuQsMJEm91fdnRX6l3VmZNl5dtosG3hE4SisXVqnMrIGFGjUoEZ7T2c5s2
ob78TfQp8maIFLtCbU0NeJwpPkX8X0RCsIeT20rxgvs0HuEZ1kGl+SEo/ZTJcZX5hpMYL9CyFAms
e8IGAUNurn/wNcuej0T6iNznEMPLEc+6X9kMjNAg+fXsuAvKGEsFK52vTV1r9gv+K7l0Q1QE5HBB
rwP9t5rS+5mxAqXp6kIBUnGq92Td7ORInsTEFNa/Eqf+kdzCFDOhzvGONETbDXpFPmZ8r4Ztx7/K
HQskozfKNsYwx7sqPr3bzMXQubwpHw0ngexHaWc203aTF2PvZj6tYsNb1u/yCIz6KFftw416bxKv
46UX5XYwFdfkybIXHlhw1zGjF7UlhhI90Nsm2+xbcCYi8kEh3s+56yY879cM29PU3GIv/iWdI9hy
IXFm3/1gVoCwq8I7OPVmfCoYqLjrCe/NvEPKufR49dBkSksGXO3G2lxLwsDt6pz6yaJ3nhf7JqeB
0uXERn9ei08Di1VaQGIYBL8V9yf1Qzoegz5jZYSsGvqbNquBCTeYvkjfPrPQwCKoMI4e0ABT1ES/
t0NAdj6NA40p9LSRVGrcMb7PNTTLhgAIxIigOBHiwYGjhJVOeWmBKvXF6U2An0bDO4sn3c7U/D6T
cB2Aqm0+yyGmJFrO+HJPG9qvmckkxtKL3XFp8ebnc6olBLrPOeQj8ElwqfhqGPY5F+SpFHLWP57L
+maMDWZtnUrzCBfFwt0B2V1D5Jkud7C+AY57mkVLwGByE98hKvUhmemePvQN0nulgsFcff6SwAKp
S5Rk841/QtdZ4D4PSJ2cTrxBHF1npTXosW4Z7/VHRgglFDVv6kRKJ+4km1Np/IIQhZibwxX6tMpc
b/96+IuZYaGeBufFgWAoG9XEUf38WRWCT2Xwctvieyeij+eYW4wJmPpxL9vw9nkYSuWFKNRBfzP4
GVAQi4oTT6V/EpOfzaD2XUhMYfmpduTUWEfXXLbGtMdcUHyQMWbs+o/jjLhlONPoUC7uHf1h0Qnk
lpcVQnEHcc8pkEViARar4/qIfO5lcQv32PmUAc7FcedOzTRXOiktdlv5CEEDT4M2WYCFxC5Rt1Zq
yJZ+uANSPIh+/EMNym+VjmMltDmvk/aWk4TtjviEu0XyjRrAcbkMDA8OqW/7hPozZaOARmQKkPwJ
NR6oBmNSRKeXXMzKi24ogY4dauShpm1LrvzPsHTB+8BZNOCKhg56GOwoRQiDTy+XWzsV+dMYybY/
dkP+rn2EBLU0Vm06efP/Yc2IZs/+mOkZ9zd+4cnBjZwcm3dfbmeUrDSimS3HaveVnDt4YFg2EjJr
7IUxtSjzhUpreRu6mbYn4WbBoH1CXgqhJgdL0YZ2HG8Xa+ar99iIDlYZ4pAv+sqlUvljwvUhhvMw
dj7gfn5Th4899kyKCiEZmkID8TXqOVqfE0ncALtC13ITxgC7WNT131aZOfc+Q1RJSFmMWiA907oD
nccMq6jRI1FjjM+2BEDIyqrX4ep5Hey9JKKG0tIGUnxXbIF8mbDIvL8PCCYLZH6seCbe0EnWFPEa
SaEJqoXHEC95etUkEH8N06TB1jsow+GpzeRgNN94b4vRgTxEBxN0xyFGHPKcCgkwKp4ARweZnbKS
IwT7joNTrHtxslFw3WLSg2QPuetmBYlKOzc5EX0Ik4W2GcOpf8zqdWhfBEjGmNHuz5moJWThHUGT
Nx7+12VpaTwppkuYCzVifvoir4S6A5h/76YkJk1eSDeHkxm+DHHRTiq5Pgkc0WRI+f9CsMonSqkw
zlMNzhF1pmFEc+OQ8ISAQzHdDvJk8SkXgN4kA5YnifNE7+3gt4pwlM8fc4hb3jqVhk5RvLXHKyps
GMKpW/xP8ERsBmiHp6HLY94P/TgOauE89/LYQAGiAQnDVCTILYJYk5uDohaZcNJBL+lELg18CXsW
wHMzhRrzn24f+/VRkLVQZN2SZOQ4wyN6gOMM/ftTUqHYjc3skVeVQ3OH0ycWT/+WjXc1g4/57Oon
uInB3iernrIcT9lYfI28UhH+NOcyOvNMEp/Y67dG/qyICb689QGEvJtVNWTwngO7bbf3sFnaBAFj
ovFNGY4zcLEm+SwesnJPdy8k7LWrf39+ju7DGHzW4+/gpxMxAaqerf+M9IbYbLy7vzt4Bf2QEOmf
PU92JrVXe5zNj44G6FeQ5BdNFJ1Tv4LXNtGDE64el7JBWgllzYtd9L0MWpHXLboUP9/doonlqk79
WvC7J7avhWzTzC56FgH35vPgtp8DvhMtL+HnFhurj8MUyOZHwEkjoO5K9FKVRPF9ygTT/7VPpsUw
TRDQq+P2PS/ZvMeVonkqLX0fV6ZIk5rXF5Hz72S8pjZR3Hpfse6EZgbMRu2xL6HLTXzlPZB77vIx
DB7HiUV+abWSgsv7ttRpzpz3DwCkT6d9AIGZlZ9INHEl2MAZnZMWzFsVbFC22FolGzTVy2I7Cri0
M+97E4o37EiPTpJgGVdDwIV8FWouZyOawyyB8x25f8xhJ1+10Gj5tlSexlx4CGEklFMH0vgIARLw
8v+UoGDlmo/w7MoN5zQoSn6zIqL3w8aRmg/R344+pvJbdvuSUFSUW6v5jp0mIo9VdvyVpAI9OH06
j1MQHosGy6QdiawytmUtZ3sdMFTQ3dN7bOZWAKRJLoZF2IaeOEBrTVw6dVdAqZNsrbkHoH9VfGS4
BaX5+dj5liOLg7ACYwqkh/6FnLlWPWmM2RpbU5fzWnhDP0/OwMM17RxMA4kgDBhfmhw+ZN141Omn
wsFlHDdVnx4qovT0UtXb9fPEfruTif8XDowaWyqg2j+yalxW9bjXScJ+gJNIIhNRMtU2GJuS/DlE
sghshoJ5DK6F1EjzFYYAW7ce3yh7MtOBDz7esf7qIYX35u6Mo04FPyENvFv2IB29cSdUzWuCkZk/
SmgNKRhSxKRQbup5o+E5xbkGVjKMVNLCVrrvQhc0KP3Oy1hNeqYT/VC7FreOwlbbkv2CcbHuzl4I
PPUVVTlm7kZXGT4Z2jExNJoyQwWSTdmvnHJtSp7yY+xN6r+jqE6tR2l2toQxBBqRi7xBAaP0pZVt
fvPux+4ttkdm6srSY3JBq5TfnAPf+hddjL/Bi+rccafNM0HF44/Tk94ebjzYG3nkmMcwvwh28Heb
FhAjIe+4jgizxC/mlrmB4BrOfbl20+9tGhCNuff4G/ThiNmBV1l1y84fObuBne8nXIxTyOZjiID2
KZ+jV2JtA0+cZ5wJIdCcI7lDBZE1aG7djI7aow+HPx2G8nxpqLxGDQisvsh9hotViT21Fy+5OhKH
DorfdRkAYheDFcvhG2Z4u6Cy29o/I1tiXR1mu1TEaU7dUgBDvRl5E8xAwkJAyJgAQqJ9BWuwTh+4
/2Rhg/5sNO3Qjvx44nCz8rRnHG94fDdUG8vzyvzowYamUVkjwJg6JRtyhmTbyOqs+8a0++czoy7E
YlJJUrhJ6pmHNWsX7Qm9mguDPfQ+I3Mgw1bUVN7nesmxZo21RtzRFaZn8y98WRuHiXijKPw2+Tj+
U94hrQorGvZ1LRWqXbcPI8xtNBts1/Z+qIsOS3I8ycbr8HeWxzgtclNfCuiOSJNFF5KXsZUNMHyM
cB22KbNAjNmqeF50SRDjlAdbhDSCaBYl6snV2y+qiZyriytOXM+9GwAQK1HFxV+OTpl9jemVc1dL
sgl/9q912qDWd0H5BGySvGCA9uAuWXjKWuRAhG4SYBd9ZylfZrOT2x7Lhs/6aFJVoIb3o4Etvch5
MoTkjiwnRmH43Zt51MDHRomcooxlcVNq5Y2QutE3GwEtl/DYNJvOnSY0OfAJovXcfuLGsVBYYt5S
WlOQ3XwqiKkUVt7O8AdZmWMNLxyh1ZWrNgSKBZDhJgXCmdeeemvRRDRcJ8VtoJmF4icRAo42VhOR
ozThLOgM/fyl0+H3oIKBvvrTBboXn8IazwIm3FoExPkI3TjudFQJ7L3ySFjAzY6AibzA25W9fcMD
c3JUqY2H3RHLy3iDj/cNOdYhHzf/xLtNidFS2ihYc8L6GoyzeX0HdQVcppsDiIrcuVTt9GcwgfX+
uBf64MZNKREs8fd0v/RpdYnz+G2X8S2nPH/KNymCizazjYn6mEA8Eere6pkll9v+Gkb2mlQRNffW
p4cZicE1eMlZ8+8HayoOHHp0WQ0u2q/6O1GTuDN0B7OCk30xW8Vg5pZjRe1uL/8SPVw286Rsmnkv
gPjWMf+h05W38nxvXMGjFmdx2vPgdDe5m14++Fj2wwAye98pLURFk0w2h/WxeBgloF+hcogpYXLs
Pi3WJVO/cuOOjQKYMrloIvdte/hBMdwkaSHvvNAoMKmekHgjc/ZEzC0bRIsWrRsRUxEcQV8gHKUq
PARmpiujpfyn1Qp4bRRgKzafeFFwzjuCGZA1LQOt9GNNGbDiZOnJo+5eHNhqFSHlbU6IuQSfks9D
WW209MOzEioeW1bKzjQoyjuscU7njHuhyDEOi+xUe5fIdZuVuPEnQDHvRv7aFU6RfmlJc8CeQ4mW
MxOujB6wzRm8SamguqY9ZUTXIw1DJqJFnmujhD255e/i7Jc+K3iP7n6qUtfAKP2lOwypJWgOjShK
vJpYlmzi8OrlawmYhCSZhBbzp41VXMmVPctK7flVz/JFOLBePn9uEDXE6MuEcHJtuvMRmZAdwHUf
uTnJMDKaXoJx1GF4dHzi6J5j9TEKKfF9Zg7vW0kSzkSAVpoyDaV/xYNfFAzXzVwpjxZnSTDDP6DR
nTC9mIBr6OjcymM5y5/QCajG86c822+9ixcrABJf1SRK3GJ2jLM6yYi5gfkUFmpXsobTaxQBm2ll
0IcY3tgx5VTEY6DmdPEyZDdVf1tLPHN4xauTp2ED8jYvDEpA3Msd2mTjqWb7e996KfC2Zz6YR5Gx
r6BNCG6jc6frJiFxMZNEiJUEKPK04/diVwuLF3ANKCLDb7voNdvKh9+Rkzz23oTZEovA4FO2mEPo
z3yVjPaMG9QaykZc4pOVU2ufTiW7Qj3y4dAYhfJ79YQffLccQyn6c9Ehb2r1bgbQdp7E8zeotzHh
B384wOevh6J/m/RykrWKbx/YbL15Yz8ciwXBe1T88rfmuI7zDjVOusLPM6e4w6pp6WCc9Pv1ar5j
+3/BAz7kv3L1RUXQYFaUTaHD8DHbW6v+PqENywZug5LvwvtBcmkNvALeTduHqdYIVMAobkgLVAfR
rox58dTcGzIv5xtEU9Kn8LtrCSsv7Bwos95l9aH21V7m513Qrh6ach2SEH9tROl8CEHI8VhZ3P0D
ZdyMpXI7aDspzC3oKbnxduCs3DR9QQ7UVZUyRT2oWF/SxT//iI9SHzdQtv2fbNbJ1tAv8xYl0Ogn
tA3MAhZ6451OOOqRGXQ23kfhqUeYpHUByaul9mvpCpaJQeuDfwDtQxRzwr94psfeD/9ba21S+3N8
8DnAX6C/UxK5ZJtYGz6aBTnwmAUGG1CkAZjuerQknc3jwws3Yo+mX4Y+jmgy6q3d8Mcy8jxv7pJw
tSaKGLu/2hUcT/gVAuGi4TbFLHzlRBlXT8sEQ0ANg1C5uWPRv1BtS84UfsLgI2H4hvy+2AnIuMdw
WXDjtWKak+Dmv8GLGduPRxx8xHauwxYRtMARdu291EFvecdO/6OE1esItnMtCGZe3D3mvd4uHAyc
dAk6RsOa2FgInxwY8TPwvE1Z/HADYqmMrRwv4QDXFYReKNBWAh27Pc6IZ9+TYdv65PTAOgylQqqD
RVybysCUqqPFMnY6wWDGlS9Y/WPV4RRkNbFgDITelrJ8qno4FEbORQ0Kc9OJ2vx2JljOBrlObHys
a8Vzmn2odrio1LoklacWYEu3KyVMgHu7jmSosJWVAhDlBmvSzMWWndUHtx+KbVkqKSz04Z/mNVku
3Vd1YRhtFFPkKtHzBMydZBWQpIjSTE43I7mzfkkRDVX9PbkR4RN9waezLPELLWRZiGyk9mzQxlTz
7RCuFATdqT7VI9/bqrjGLG5pLaxfYElKf/5HRt7eRMzAfn9afrfdM4s9YUp0QQeVWtYtL68YYacc
3CIUOa0Dg+Czk/5F+QNREKRImrchCz8CifePIr31JJIZEduozdK/brvruEuAyEa0eXQeahsBgS8N
ww2nd9IyAP3ZalldrG87A00M3Y9OCHx374uj/LgAHWcyrXFB3/CbEwRg6MRsjLbRxS4RZDIfKd6K
Z+3vsJ397zZJpij/dL0tXFmGlZ2Ci6CiapChli9wb2W6MXd+uWBACAZ6+2iYbsj9gEQrGZL+Sq5Q
Iruwzml0gtlWTyxM7STjbu4dFYkdh+RR1zH6Dk8pzOQIX5Od5BcCnvkBJlst6FvTWfqYUXnvND2o
WmEyh+F5aVXjTcvVRNHQ/NG7guCpXKyYUpdCrQBrGnsxg9Kw6JqJ2pGIGPzFc+cqZNxYtT7eT+1v
eLPQygj/KoljjrHK7WaCzOPLreTZ/drbimnuX9EI4XQP8x0ONOiO3xCPKXLhjkPBgLw2EjcK4sR0
4At+OF5HkC4MUBYwgsA76t6FoVvqr7YDCQYHuzRVK5SfPzIotWSEqXZTZmuJ2tLeN1oTbgUi96fG
TfUa3XEtXyqGlFX1nHEAgrAwsBIo5zYmJZs/Am/VZ6eUWimiyuBU3ii2SLlHqqatWItB6nB4gy9C
lcYJsu9sHgVFahlkdoz4UHC/SDW3MpQlg4iVckPwxkFj6mKcJp1Co3fvkiGr0tWbl2z08WUNgNXl
JHbT/UyjugKKOiuVZGi3ZvxxpvLLjCEhcO77piafe5Y7cwLG1UeIOyOQ8iq1lkNuVFVbBVg98vwb
ROiHr6HIPAqWWIb1AWR1XBCHB63i6pSQeb1Sg+Zw6seGRsfqmLWxQq3sqUsAo59Tm4To9BHi54AQ
P3sqoqiXOm7WppV6Z+jXn9CaEMjwH4rZ90QwgvjttR946ChKOpngaqXHGLffycaYMd0NxxyNwSN6
oeN5/67hrb1LEQ1wnsbGq6mkYfyWpSnM3P4z2CbCPLLnvLqI50ULElMtkuFyCunIByhJijJwdSPS
JZV6AQ85OeAvaj6JGyPK/GVLg8WRcYa1tmpRUVhaT/K8tKj3+/bVuxUBRkA5FUBR5KCfwikMmu4B
1L/Bo0UGrQ2uFG5RnmWRoyQSGgY058uvuuiVIqYIgGwV0N6h7v5OWEFUY9d6bNm8XC0KBIC+N5ig
2SBzF/mGewt1rsEd0J+diUJWfpxfngB/zBNz/87pJrXPFnFe2+fm6u6iKTdPpVxuWp8wdOCvTdK3
///c8j7pHdiZOgCSYIprdjZvFTyLE6cKwHJFmw9CHQU9bdENgfmjnuBNnco0oPB2ul/H8epFSF58
uc3cFpv/S6/cqRoTYkYdSPEOt6CPKIyiyRbT4iA+vC3U1DBzT6smqqpHIbJ9hIbFHxkWYqhi9Ecr
yQ2pRZqSWvok9ffwJ+q44hYE9C5klLJoDObJpkMJNrEL4F+wJnw/15UUIYFkF3TjbUyLFxXNegll
BkbU7hn5qC8BaxRimEso1oeaGllw2ytS/mC1rbXjyS2CN1iG431hyaBXvaLuj3z52JPrni/UAZqi
V4S/8bYCtlLRv5lKezP2sIIYSG4NLj1fZ8/1dj0Iw2DKuiWFiqhIQdLdZenlgmjkBRx7c2Q75ksa
7ZKjjYmYGSXp/eyaC8pzNRMTkoDoGTEZ2xhvGGMZuNupHs/hAD98Ns0JCkKAFhR6BQIQrN6Hl4N1
+cwVgIHnUn4iw0A+sQm6qVnqiL2TD1YjTu9NrcXnYziAWhi3HE9YRPBNsGn5w1bc9Z5+lf/YtM+W
v0Go8y6Z2IuVM08+RFcn3hrax8Soxkcjv4C7ge463WRKPjVldWidykdlxzanU8zTLHeFXtBGqW74
pXQl2zSsfhKol1ppr7qPtAp2SKtf4x8xlbrH+IFiwNHJxBN21VYSyVE1Dx0y68zaqgdIcb0Jyc3R
7Td8jW2vBaVxUrgRo2Zzkyd3z6FElUrd2c9An58/fyziYhVEB52gViOT9Lp+tRAvI5OnOwDCDA6S
W72fD2Q3RInY3qaop0JaUz1npDVhfpWdngpKQiu2KYWp0ciHQxX/9KiQulF37eY57VhqfJaT023r
M67P6RfG/qyXcHjbr8XHupR0SBUUvbaNAlz5kSVwFb3iyFcEmx5Ys6NFz42dwg96Qkzc1Kt1jStK
HpiA9RSxBwzJkxs3lPxKDSoAcy7AwMPyQdYeeEcE8YOS4oJLfO5USU2o3OR9R1ihyxHub+UrgGlg
+U8ckwdK2AEzXp9kvamYV6mR3rcgxKYrK7aoTbEKh3VioM3Md6rJVsy5vgLPLvPRdyu6cuNUAGp1
uDILh6Bt5GvbgjH2YbwZ0cQY8Rw+9Cwn5sNAHFqzDpBhpVc4JZTAXtvba2cWDT+g6L3ROBgW+BK+
FM5uzRaZqYZmUclt987oF3FDOU6iIvaGUirCKK1ipS9Jip/2DG+9NU9lcNGkZmjN79aR3SyC8c0x
2IloiJ4H2RdB/2r9SSZ72yiXggucJwqeNyqpzQ/04+Ocb8LWA0uIMy31OaPDS8PTWu9HTxtpSb8m
9QsuGLwIV4n6qpHvoHKkdLe2/hI4Il7lmK9wmSWLIQq8NT+tzcnNsXV66qRjwykYZnVq0wQDu9PQ
ePc+oYqPkb8vjtWZMIAThcKDlsH3R/IapwVI/YNedkxTBc1BTidA7Yen37zUdPFUXsUSSN9hr9Om
dNMBAjht5wy101iW1OALBxebjXJcpzZ7M/qVOIPe+XAov0x6MrnIxSOlL5cipiIVW+D/2JoJxF7X
f1N/0qnxKrNabB6d6R1D62+88kvVvjG3qlRcTHSUkUFuDn4ytHwu5No4S2VnFbQk3MGiCJlNS+UC
tkxcmDbZG9SUNFYa07up1SKaDh3iYed17nL+VsCZ9yuTdWX63r5HXSbXNTXC3qjzszX5FL5b15br
pqzEnFf0F6I6VbGL08cTyvfouMo7wG2nfY/NkMmOeT0gmd1tj4aBYj3Q6rVX/L2VtlNv392gZkbN
Z/RVvEDEcAg637jkjS4E4vBwGnAxqaMKPACaiVoKrNm/+M9icRkCRan5vnUzXEeFgG5zb2cTxB2u
/nycf1G0Nm5EAR4HOtlY/wP53M262PNPH2rziKMAzp1ilCYQ7rJ/NqJaCUlwKLgaObs3wv3PtZiO
zkAWlAKyffPSm6vFVhCe/Uy/Ek74+SYnrwXoKuVNZry1AzW31VrbaxnSSax75UC5U/QpbrTD27wy
LPkGpqrYfY+eF5GU2wMDl896GdqqmkSMm1INeaqHhfD1zgqBE6OUAgyu8mFhUf2WRHXWOCpqEDM+
1IyH0x9Ao0dfIVXPG+/VaqeVoPxOwcty989F14wt2RZn9yYhaQNmA0H9gUYDKHn98toos4zWOEOy
s+cmqivf6AdAGuM9fcse6rECOuMYhQK+/5r1461+ZpBqqmji54EgSKbgx2IeiOyZH46F4A3qSQ20
E9ENZArXN8WBhx6wNvqGIzx2dnqTP+29cV92RF9IOTgrqE0BSKOxwaxLaYvHZexxwhkZ7NwIP7U/
YQxb2q+yTNsTFaBurJQtwBJ4PS9Z3aagARlPUvtFuWokj1BzdK1q+ewwPmjaVd4P911khgZVDy6x
auvdxL3mPxkBxLB5n6Rfkk9NqgsSrrDRqps9G3cVmUsHvcUNs4CC9Xd8LvxUArAQDyERVLB66phD
xnIiEN5UD5WM/XgFBLjyNll0rB6au5aNBXYv/Jt3dNJT5qkilUnPLjnBlnOgr40gQU430pQ5v5hr
eRxqi1g5fN/XVBfnHhKoiGLND5bK/N0H453uW34/1vtJIb407D9/88ifetFrVtw9P/rt8eQY/Gn6
rrhpP2H9BzB4qtkmrZEPQrJjaCgHBl2VzzmQBFH3Jkpx6JZMFgUlyiww+H5MKwTBkciCO7TUbJr7
TSA9GifCW7WjUJSJ5nz+yC67yK6EyC14KdLIM21xPkJpBpvXolAx3Jtm2/hsZp0MX5Qj+RKE+Qtf
EEQqMO+B60hbi3GThCQ9BnBkruqYMIiL0YuE96m8k3N+M/i0rHEecfGLAJSgw2j9PFEOR+3ENxDK
tw9o5GDaMprRuBGPZxCawge9XG2VAIWhub7OsJRcmvn/Z4hCcl5y9z7rvtvOYNySFH9CQ4JMrCR8
+z4QmvkvdPDwlEOh+WHAclec/YmCKV3nQb4ThAdOgoBfkedIaVkRfznQxAquhhebhqwzpXN8XHmY
SJqpAlyfFM4VcQ8GA4BrhYDNQoeTYd6e6PFWnv32iLoAPaLKgT8jqNDq4bA+oBQlFHZDihTplOWD
gikBuRJwHdU8/CH8UOMcyRh1tFL942YouqneVFW7b9Z/ChaPwR2iX38vPekGeoEaHbQyTNy7lViJ
f7KAYjQOj4D0GR04Q/rmNPssujsLy7G30Fpg2UAbnUurxfyGEk6JTEJSQcr0dkDg/j3zK3vH22BX
Va35oMewLEs/FAYRdgbOEScnB01pGjJmX1EstJVIvImGYOthppnPgJuI04WEv3KFhAz+/BmlfQeL
mZ/nh59eItEZQ5JYpNA/x8rEVS5Ksea7D60ilLytnSgcFhyFkdBgZXwPpmxlLyqQA4eKzCmkT8fR
LineL9Ww8QI6t4jmcmTULryQIXZlMEoRjLXGehnAPuH0k3XX6HfAm582qWCYVjVEaoFc7BZOMKwz
C35pCw6FUQvacGvBnmPE3tYt/FgecHeh/OnqigUg32u4UcMQ2/CsnPKyIn2DDvbc/GGWpMxp7DS2
2f9Y14QgiD1iK1C4vwemLn2r3C4pDyJxKdFxAE+L7TBwdBFvmzskRKqU1dkiJF43+cglLMDWnC51
PhkC4aL3oWNtRA1ZGFX/xxJhPcoMEuXtzLmpEsqjzicrhDeGM27KOnXBx8GaDwcSgBkKDte6GwbC
2fzRy8asTmS+SZRPbbP0pvwD3gwPTidU9/WUcJwlpqNZzcKJ1XUcCJalbNMuPp/X9ElcBLBset1t
7PkvcDjBH/Zjwfxq/MpjwbCch+7YHJY7Ho3QT9KzTPC5Ot5M8QTma5SjRedCx2aKWmG3jyigIUg0
nFOpzBKCUyijxcCM3QKy3c4nW+pPDOVr7x4M4JHvVttwbiiae8J9b+3qYAl9Yi97BnFq74/jEJns
AKkSCR1WJ8yd6+RVR6iacreWtpSt2en49kCOtFfr4sG6kUW/qz7+E7qQRsaa8ffX5u+hka0vkdsq
TY9pF8iQkHuaFvooQrdwu1hm0EG3+1u5cXxfcrmaH5J0ZlPKasgvwmCWESbLmTgH3mru0ZMIgGjC
zWEXHKFWjMGFcVsh7isKMfhTVKpgaJH8z2oql1el1ojT+yIMqgnOhJXr9+UVICqq/AW+gUdO8Ife
ppq3DBIkHOaVemqvlI4fTcOyCX92ibDFdZ1bX5289T0D09m39/UYOyRlxZsdUigDfKkqqs4kZ4vw
iDgss54iXGLNqGjDETixkGNA202fG9v9DHyM/1su5gSmCcv3P/y77DkQ6Voo2eTFgx708vLu1mgV
7HWTiJDDgpH7ffZnhoUfAAttTqGMbDzfFjlEx45b9og32IFbY36D5dV3/nCK01ftwpZTZUayhgSp
rd5/f6szP8KIkcO6uXZXaWd+CleEyiYXnVAuBT254gtK4v+7CDyeOujbWu8JuGZOmoPfkq0JZQPa
M1ZY+gJ2gQRrG90m4Ix2yWpB4zMI/dZWO2bUEz6TbgwZ4H8z23rv6Wu7gUyZJ/VRqpCWE6S5DjZN
oJbD44OwQdhceoiPvHUQ4pVYufqmCQrlVqINJBbm1kDlb2XGuiNYEcL36ugRcUbnL6zRXFNLui4V
jDTWB2L0aioFLomknDUaF7+9FoZyvvGvhxccjgt2A6GaXlrW/+iJ++Cay4IRMVxbMiXCZAS7LIrq
j+4UeuZmbhrGc1MM5fYYCsuYDZ4xG7sm9zMh9KqeMG77XXmi8OJzfEEobRYVDkH2jqD//EKOc4uV
O6ViXibL3b1N5yU6n3404hxHR/S/ZaTwzdayMyK5BcAbmZyrimIB1MCKSZWsJlwNqKicIz6sc9p4
Px7pI6SXM2RqEYGmiZeSq4Klmpw3CKrGK8s9FWeNa0p7RRp22jUtybp73KsXSCFB68uAlco2U82e
wXAuH8rctO9sEPXO0lLpWQLR3DuXlJud3jp7nIcWQMTZ70UxxkokQxS97fhHhT0+0ev9r3L65Mcb
MYUUxp+YgeOK7iet36iQ1G/ngHHPVXLiOwGAe8IYvG3+A6K6x1hxv1P/0af7BOHQzyvAaPpACoia
/siMCicYowlKgn+Uq2utRuh99N1j327jyTXQB8OlS/09YU9oijdHzOSfcKHSqxf183b2q5Vr3TBr
tLXN9gvLPIlAGf+2RnGVlCs8FtjhBtjm/e1/3bBoutzdC2NJuWw4hXtFyd41mbXr3GqvdRxj+qxE
mXCbHdRFnGH2F9OmWhW9/qzTSlHnY72cnl3JBG8Wha4p+ZnqpQqvOVQv4sjVXdyefgEhMHk9hV9g
3IMmPZdntgCM2nC4fu3rWxH21ynhO8UDxpmppZMBp/xxwo7c7L67r9OCQUIHPyjWd2zQjCZcSRxA
JdTSisInJ+JjJqIKO2roS3U2QnU6kVxQiNnVX6vXh6FbZMhbP/bz1Gr28OnA97+uC7DkED36Yyes
0hwJH/UtTJGaGh28joNZAuaOn1ZVB8dz7DJ56jfKKf/dYkSkkLeWw5OA7Iqwu09hgw7h7TeqaI3v
GbiKlm8DjOD+iitRbFj2KFjLwkTBMxKibCSo5q/qRJLVmpFykeVnq00XGUaVQ32aGzjczYK5spvG
uBZhPBafYg+f2w+S4xHbsKSzvWDi5lNXnamL7ByTDeTZnNG+NmB8m7hT9fmKzj7Wy0kBACg7ecGh
l7c0EH5No504WeIoDJzpuPkhmLyH1Po1OY1Eiv40rkGf2yvkVLy7ZehrI0ea1DHQP8qsFVzguQ9S
BQ/ps6YzK5IoLPli1Zp5DJShXt5D+SOHX7aFjejSKxzNiVZ/VBAKuB2QUiP+s5c+jAVszC0Hyuau
ATi+rgXcs3mmnycuf/++6WdHAIXo5vd3yg+Y3xi3IRZYs4PpoZbNh1xVFTY7CiStgjTWTG94Svm7
e/4rW5h+vao2LFktT+3z0SY70OupWQuNXO4ykJ7Cj0Ho8HwEgnvhqEQxtDtnaUZh01mliqG6gR3G
pDqdoUPCPtne9xvGjb5lEG/4bWGy4+T26FY9QcivKpbAZFOLkDeky1zLrZu5AJ2hdriElV9yYN5S
Q5R9XUGi+cUsBScedy/04zbaGA5YQlOW6r+4UJ0Bv/WM/TU8u3jNBiS2s7vbdsVGQgEeeKU7X/zI
d6rEiiklNptfQQYf71zsCzKeqHTpFunBuehxGSnegL2NAgoWo+t8UPzM82OdMhnz0Rko7h2Yz5AN
ClU6mTeozPVdoNVA8Ru3+jbcBsu96fwrTczDTxRN+1wSyPyPu2IBXb7+20u7kg7VpOVvFaftILD+
jUvEaKAHmUmA+WclMF0paP4PC1/9QbXRDQLbSJjx/3UmHYxj6b09YFSB083GEfrwx9G9bsbJ04px
loeQcirkoHEOEiHYfTP9OZ5uG7N3UJRgtPHwCC/RaUMQ9Pb4LQZPZZVIZcll1ar9hZwOtK8c3VOv
okIVFKQPYoCdBUbuRwRDpnoYeXpIrMPo5eME0qZOgphjIwphLRviQGnC4H9aCJ8fQe+195nVcTOh
5Sz6JQVvXDPC/aYNMPhMQcL3YKaiwaGb/QHBcQgzE875Srvg7bYDVn3byb8Hi87ko8o+qrS4kNI5
vSXzOVGUig4AK85vrkwEnn/+5hN9qnH3wazAVMKTg0beKr+NvCDLGqXwKlt/DLdsAO151mTKhNvT
9Y9dEkKz2ugWwRW/MvvLF5b5pDbfNLehvK/RKVt/uF+zt86QYEBE9X23zXp1F4FpQ5s77GUWcK6k
iB1J9CR3u/qFtIYCs5DYhbZ4e5oRoNg8afNtUmcQ3VIRvlilJV4XPKVaW7G4Y2semeTRykEhyh6C
J8qp7dxodUXYsjp2NNQ25ZPdJp+tM2JdEvTm8ZiWFBH1JYaxYNTXg7fcXJsPXUTtedEm8O6Jlhg1
HuujcMuIyQ7cATmdlnGaT3Mtb1iTZCE/cBcOJGpzMGNDiB6+mvx7FbnXT+ZUlvr5fzWP9Zak2mNA
MQVG+tHKabCRRPF1ukJc0ch6Som5jLy1ntS9Aw+rkL7LcGjd065EfuahQ4qiXkn7VEXm1FmnWwT4
nMcMyg3Rv4DJYYQE1whdHoy6tX/JOJ6X51prDsan5iY+yTRAObwCJs92+ishLmSvTsEW8yg/esKx
YOfxMBRrRFZLXAQqO87+/eFQqfPRWXsz6WPxHNFckSeTg/KG8z42OF9nLpmF13yuS+/Na0hGuz7e
RAoZCuRza0KC5MgVMgkifABTt6TuMz3oMK4RO9uM5nY8ALBuxSsbR33aAEEoVXgtqCSH7/6mlU/W
ccJJcEihVbEodyB4AvMLsYGhM2uIVi6rXDF1qR0Nf50EdHPuK8Qrz47U+8ANA+Y10YfInk09bZEW
aEiI+ZkygnGxMU2FwlGPbTWc3D1Jdidajb7vEo0UMRPvvv+dl9VfAyuKByLKaZgm1gC0z2fNOjvq
cqIIvoXu/cqDFwjQ9nstLQsxm/pH6uPPIPxkpuf81ZFGnY5LLEouj7kQNEXP5RTMVQgXQrEH6mZa
dbKqfAD0ZYgIJ2l23Nmfch00TkkCwt3VFVMvc71gfItW9T7MpztH6IYMS947DiYelK3xontSns0S
hlr+GVHUXh9RF4pXbXaz4/5MmZcCDWdNq92CCqRo0z0fu69Q8afC8WGbcJHe14FiBnoLM1qASB3c
CPzOU4cRiFZKRSg2pqyC5Ye2miuBfdXTdPpIzRABGG48+3UqU/O4lhWSwhAEeq9LYYa75It8Zwdy
0LKRsNJXM/enYpzJQX5nziQzngIK044ErX4TbCDj6o07LHNMW6nPqJMV03ZhrkdQVAZfdF7vjzby
w2xjXOn2GQpkNbIFUVeaBa//RLEOK3eQiIMUi/8L2+s8XBNpMjfspToTnjhMssV4C87aMmb4I5WA
i5nMPB6JtLoqsa6kjJwjcd8HJeAp5KjgaRhFAx39hBRR1LRRU3TY7986giaN3gLMey5VFtwNV0oc
HMSKUQCDtjq+84/5EweuMbnjkvQraYesNTpQM3+1LLV9N1XHza9u7Q+Xohf05vYHPyorgfeQxYTE
NhcDO1Qr7KnQT1YAwspI1LJW94eu02t82qQquxkjBTXUMeE/UJuBoGqTXOWDejmb/AVk3ca8z6lY
44BcCB7yivhLaKGpLPFgQTs8eTH4m/jtUTGnUeQsmtN5IlqDis3HVcZ3ciC57I3PGyIjvRoHcakb
vL91SiQSCH4BTZRN6U5/af7sE/pgpVOogQZbR75qfFttki2HKuxmHCySUjK+nEjVEU2ekymZtEWA
7TI5OoYOvXPvIrh7nGWHdgSa0XuXsI3737+Pnwx+pKvbInpfgYKYWbksUTZySvrXWFTUAQA6zYhk
tkq+PUxnyS162DEwFuNk8Ed+P6x27Z4y38LAiLHshCocBNbhuX1l7oZJolHsuUgfiU811dPBbgB3
kXG0yN50W0AU+/cwzoh2pIODYulcN+aBCT+9Mno9prEYAKPrnVvTuT6gI6R7Qfp31Ea+1J6ZHZe7
TOSiF66jZ8/DlVF2dEi2zD5fEBFgQETu+Y68HvwWQpYYmeu/9YG9gv07HdDtTODY3NVytVjF7GuE
SCE2s2k3jCKCC51dIOyTIIV7xn2YdME9RZQHiJgJpHpCbOx70l2pCP5A/1fkxNE83XsytFqjx9KN
as8/kod3w4iM4w3WKd6FCU7W90mZiwrj3ElVYtTgFdqaue9fFWRSb6+Wxe51TMCNeifA/mCJ5aV0
vtIQBnXwe8eXblASKSHS9kVivXD1Y/X2Wqq93ZP5L2aUmfcAOR3AEMUamyw4VM8Il+Xk5Z5vKBhe
M0EBRAk+qbhDBmdRGueR75cy160TpD8dD6FAuELSc1Q4+Aim/2vYGHGUE+1IBzU5hU3mHLddUsci
ceYY5pu0HRK1VWTyUlGm1Xovp9YCp3FLgVbcqnGPC/SBFcowyA7Q7jgvIK6W9dAVHlrqBfj6AcIF
spV5sD3jwVeCfrkmNjncGFG2StndzYlzjMRc4FfjnTcTrTY2SwXGYB2Uhu6Dterxv0lUWWxe0dJ7
Znf2G0gIhtlsH56o54HCdWrutGelPDDO2e3rmXZZE65LYTbBfJREX+UIMcreMmxuDgrK3+DwRpkC
60lYL1QFMzNT2hNcSbCVC/nJvSz+NO5nf+5c+hFk6UmzkeTBIwGdeP2RjYRA+hfatvNJCaxsc9wn
orN3K2H8DD+EfNMu6PJwtSwKeKSds+Wbynsu7Tqq9BHU8kwLNG4c+5EAd3cPack+C5X6M8TZklCV
++k3cZNosPG8elk7adlyVJs7QPR0UD/g/anCSmXtVpns+BEAL7FI/canmCrZzYA77B8ME3KXHUii
xyGdG/wav2Y86iYSuqXzeDvcFOivoagYeE6Jw2o+FY5dw6tYheQwbW6PrE+7RqD4zYFnUT0fbMF7
/VmPMEDIRgUXoUi32f3erbf2HvfPeio5j+ReaqoH6oCBsFIrQra9Ge2aE2+D852r0Viofc2JNC0d
U3WYdptHMO2f41MNSc5se+D7S55WDUoAiFcLRsK9NH2Gc2wU+SmR+SxmD2VFiaxkye2UJHXII61M
fOxh5T/cto/BtdLVhbT7ogKqzO3aXoCtE9ZYi8MjfZEVtZ3S+bAH2X9ZQx7W60/hZpY0wxY1rWBK
GY4w+syeoMzTft+v3+YlNy4RI/mSBKTKMSAeMlElNa07PjXvYyLJX4zV7b4CClggBpsqmfrE1VKA
fqtAg3lYvdeAwOF/Gq6HtyphIrwgDrIIdFQmm3/IlHuRvPhsTfYzAf0aYICYwakmbaiDqfLtfD2T
GumPfVolC6U7X6bX5RDMgChHx6YmXt035tEIiwIdgpZB06T631PDQzlpbDG/sgH/nbWjFt2hpYyh
mzZpjuY2Ugb5k90jGA2h8S1kqvSgRj4ELHytQPcNm8we4AA2+5G1sPj8hO68rDJit1A+xWjpqq/x
6bByFFWW99cvX9w5NhaMpnxq1kbvHJL4ZerCxtGC3YOaWmWUtI3VeYImK9QmAlvzQdwGcerr8zsK
4J6y8MWhEXnMTEPg4DCNo9OyQnfrZorNmY+RZAcpVtg6xnEuufkpvoXV5eLnHgbXk50+WrZ6oN9o
3imh0Et14KGYoGKOOUtshCtQrTEZZY3kFJf9hWeHYJ526FnITXCAy5zwf5FUWxMG0P589UXqHJfT
qP4Q+lbWiEVKbVgRfJb4b9oHfugvRTtX290QNV4iX/jJTGvpkJelZSRZzefBcVemDK1qcTzaGTQB
pCuPyuVPhgMVzbjBvy0XJUDoGqUgsblqhDLGEcMWc6MxAxsGAouu9M7v4/zf7CCs1qowRg0KMAUp
lrsMeKDSLj1fgFllyhR3IPyzHXzUsOioG8N6bBf5dHRzxviHLkNOl455fwk9x4wKMnTd3vkOL9s+
7aSxW4J6ON4GuWQKPvOa1ALxSaVTomQP+U+NCRELho1yK/CPCsYLKc4k6BNNIBmVwdpTm56VmAC+
zUdjI/nbXvoiRClyJnIYU5Z+ua6811nj2UptIXBnAMz6yz+Ut4lw9ytKPfS3wJQerEZFkDEKlRl1
HivA6Gl51LDdXpjNjhNB+qgzHwPmIkUkZ1LXf5QxiINVKmU4KFTB4Wa0UBM6liFyT/0+5nnOA7Q/
v4uTz9PkWl9vOVjM8/NliJguZbW5jnYDoganXYDZoQqRMCHauY/i+l4xsKUOGM5+Fe1VRwVUVXdk
fGRdfJjECTvGFwODl3w5qBjQb3XLQkZT9jjFYtJ6OgcUKI7ZREKXpMDP0CiTmKeTyKnsLwlY+Qe7
AymKK3ZBcvVYwYn3za2vFldzKFXw+sOrFR+XkwrJQQ9vk47vOrlS3srfEbPIg9JIO/hk4+CXkYIt
i2cqzoSTkvqhL09Xfw9h3t9836Dm7sWGpGB1JH85+cCpipnwJ7giLTD8W8uH0SxcMtK4FAKqSLiA
csH7xw/6v50Lu8xpGinRHeqmarMixE6Axvll/xuKC8hfgG1ZcM/tslOLNKorvV8ZFnUrQTJIQJgI
LK6cC9Wa8SLW6nlnsZwEtvAnW7A2B0WqHfWsolz2BAJTqMW3ZpxRnj8FLrZHIcaX2x47zbtqknQt
2IsrGKzXxzS3DTx4wmJYuDMRslPZgXI5pulAfsjHcV9jf2P4t0K3pI2LRWPn9xBLq4pA2YPOU4Ek
0S4uKFPxhXHhTyxNDXaZ+Nr+7YunO/x6D6IXzKg9BpXGXZoyN195tCSNrM5SRVUOvvJpnbXcFP03
RiJYwbvL5nS5b5FmO8xx78fpHVaq4wmeKDCB5gUF27WiQGzNvSkf/mRBUuuE1lthcWcqyGCtet0U
Ekf5YHdXWgnIZGR63NpSJnbqLuMl5k+ZUN1H226sXGSYjNi/5pu/0mc7mLuetEFC6zHgI/EJmFO6
r3Y4jHea0Hx1+1gXsZWMPZ2GGtu1pa1zgD3/YXHVGwckRxRSQ6f9frOGehFbDyKwEOTeK4Qw0nfd
w7jGS2V5h81p1osENq1McFYNXNDR/gM5NQUHktVNIzT1a0nd5svmbV08V2J49bEUrm0ZqbSrDku6
fu45j7vZN8epaQxwezGv6fi4LaJy1pRWNZFv43LhAcD+0ZT4apm7+75OI0EAr6/RzT5A0Cx16yaa
qbkmYDA1iUOhepwYxTrN02RrolIZGs3ZCLJtyV1gxkUET53dV/Xos55YLZWcO/yN0TonFpVvwSi1
ynAAElMD3GADqvZIkB2GTtNve/5ky1fBms+/QuDd703XlxP2OmXe5mP4810Zya4faJcQnhuxcDDp
RnpEuaOCP3UCsejjbuZKixGGiyNbciTkKIYgTJ9c92g3oWzM47NzcRJ97hwBCUh2mHFb8b6SQfiz
lQpC41gsgihVpgnxBFq9BhzPfdEfiqO40rCgAetA6x3tXlrgUa9wPOY8OFUZ3DqtfE8hlGW6hzkU
zKgjsz3EchrnjXCnOn5PYjo2xCYpamcouJfWKW3YkZu8o7Yr02CMl8acrL6Xx/eJeLJ/QPGO2ovn
zmu0u3cMbbyTSw1+nc6WwzlpbOktKJTn5STh430ynm3qjRdqNtgUdJxgyzxRVUuT1+CGkcZAL0Eq
vN5Kle5txJXMEqeKjjMKKNw9N3f/7oK7lnhPxUo0uFOuzc1sdNMcySdI6DSG2TzG7Qcvhqfmf+aV
2nE7DH5YZsE+Lr6hjPqoukFKHPI409lWgBPKppXYVjJi1GcAc3p9p2ia+GtWpHN9oLmTVf3fjf09
brPBtWtyonLsXVV3Zj/WdeoOQfTTU2LcOzVMrZvypn5h96od/j3LrU38Yx6iLwHMZBzDSoRnwF5L
WZoBKAWfer3l1IFzlWdBzL+hc5PJMt2F1cx7LlKGDW6odUIwsFzf08pcdgjjLV8T8dmQnH7m+sIr
VUhYupf5cmtYjVEOq+RSi0V1zrMRFONd/0/IjUbV1GunEzdul4rt27yfYQklUKDbBnBlWnvEVH0P
YBPiaUV88qvWt9xGc24p/ADT1qtvbIU6AIOKOw/tX4x9CAZLMmGYVIdMA5JM4AMjJ33aMKtZjnnL
dNBmMOvqVj70YmTiKYLYKiNbsBBV/VFufvGXl+9qRnIn4CMHg8r+LbihfCRA+EyIPOMoaxb/y8IR
7Un+ySb9OfkVeHIrGN7g4IrKlsgr8+D8LHfGk1wMH692hNlkRGFgB75Wb+lgr3SneHZox2a9sGOz
A3jWKxQy4rwhFLkXGpqms4D+9VdoodvubtluoZQKhLgeOwxFLJg5QnRn7oOzVkgsQgn8gTmaoyNu
JZNS+mubke/HZ3Vq9cwNc+k1pwoKFzsTUWcOdjofr5caNlnL06kwzZHQeNs4oiVUQqaUE3vdtFy2
XeTjfzCt4XZ32vl5DTuGNO3v3igY0iWl+6BmkZ3Tdw1cyTSjs8LZjX3VdkRbXKQlfMX6gQ4HBodJ
+vPD9MGOPuuc7+tXiBfRc4otP+P+/CWkuLYxPpqTwlu2SQVDWKaIF8e1DpurclozAcnl9iYWNIGp
l4rCQeifelYYMYQXZmPTZP+s1Ii4WY7TL4an0joZt0GWpb22VPET5ui1RV41kBSYJ3RA2YMrnQbo
CGJ/HFaLkoEVYWtunGmJGT8YyCKP3RBflKI7kbjjNQk5PLlAkHa+0qUunEMmCu51TQrDeb5aDCEG
GQ9XoMco3UJGe1UrxOE+ZaIxac/+QHb+xVY0JDOmxkBkRkKIcgNeKNe4bQbhYUUdGO4IyNaJQd+U
RLzx8BjOE2j0G9P/dXT2ch+2jQOmStFiODfY6Wj2kVXrDJkq0WyYmFc8vN/KOM7Vlx5tRtR3uwtw
jZXV+heCY70mNId9x6rlhbNj+79XacHs2EeQOXC4XhD8Q47P6aTo0+NPh4TxlzpIsz6yQ5MQBiRq
+d3LAEKegLkM1iCcrNdyxeuXeaV5rIjXX3zWc6351l/IkNlCrBmwKnpWat+cTxjeL6NKDyHMIFUp
Ku54oCH+zYAgILdqQ0zZOfSk6S8qmKN9ATE49B0rVXN/lWcQdbqlp6iWBKMpcqwG+HrOmu1Bvn0N
2CREXQjSt8RkqMhaPiEzmgwKBYryil6cDAKnBVQ54EFZZKaFDOy84RlKENKQtKrnK/cpGO4ILq8I
lUXS9C3BYNK2r3gDSaCySIlYrOyRjeog3qO71AGFTGb58at5OsjynCB5BoEwVz3Bxuj0p596SGqy
BzLx81HNMEafT+QvxFzKUZwIMzL4JiLNrGVbXDm/Gq/Jzk53hgxvCXO54mWk4ifWNmi4FJwsnGUy
e9xr+HIKcRWDHFJikXyuJDphuK1l3zvw+pfIo7KBy3AbAZm46hKsAc0Nt9OB84ze7TbmPmlEbdT3
p0LyUw/5/2o2CS/JpuZQ0E7ji7eTqR7ElL1uHwzHKZX/eBRdOhlpHkkDBlbac7KKSjYMuuXPFInp
+wDUfJL2ZbCH6kUg7EEvlQRDhmJdIdoy9zACBcVE49JuDQo+NOnTZJx4WVx9k/VIb4VBg2EW0Cnn
w3SFzUy6S054yCsKVBzOJQNmC12yqIjFjMQkAW+004kltsrszXa2mSZ9oAgGI5y1TPIsfIgdzJQA
D4hOeb+4Ms0ZMqNM6AgDIthfL0I5I2nw80n5C5oAK9ybC5q5jusQfNyL1pH5j/xCPuxjO3CMs0Ji
Sw5lpvNsEFnDAYipAxH8GuyTzDABi0XJt9q6Aw1f7weyoM+3jXXIJ0d07u1oeTcCVVVw1RrLblqH
Ac2GvneN4PiUVjwT+AjRutLSePzPL1j2Y26rSHtNSWMZN4YI94W8Xy14Yf6pRLcVQGAdGu2oNp/Q
a1R2zsRZ7ouni55L+RSb5Y4CtPdWWF+MKpYR4VO/qwHuocogWYh+iiO04kbp7kGue85sNRnKqUYI
GgGl50iEATP2T7axp4eMDZ5WBvMZPAuI8DPOtliYYLb33cyDYPs/N3YKsm/r2pLoKrI7yzdjj8bV
lSDUQzYU0bQG3NGViEFNA+437Sw53pkbNU62+5x7em3WOdyj/vdBrCnhewbAJUsopDDK8n0kbV4R
yWFzwiwE90MLnVdHSGOSfAqkTvo+H8a01KiA/lrYkGoxTBhoZ+FkcpKObRoUzj3X7XCqyuFWF6qg
Mk3eAFIqAUApdwfTHGsqSaJY0frNg7LUn7ypxg+AixVkEf6ttWbGartLlmCjm0SivVDbmwSNci3q
6ppmWf1cJSRI1lEONoK15wsB9ZctBJVCBOsKJNzMvooJtmqmY//v8LXSq/2mejlGV8qeXdyL5uJh
NVEbaghYNNqjMaLMAdMyxdDteKFw2N5fK7ZpFaPk54MYFPnMPfqsgHHqRbsTkrrA3xTXauPPHHd7
WBPQk6Xe4sEUG+AvSUI4C1Yvs3cEoNV7qtaR4KPgvP4S/LnKGUePp2Ay0AEJHubB4Evc+5en+F+U
qMMZ7NS8dBBzGHQFdyia7zO7+C8JZm/IWCZS+ZhAcPbO0sKK+b+y0OrK9qwNQdsZJKbuWSKzJ/L/
bdOesttWaGZAqXtc83mOM9V6Iblw+RQCudp/PqkUPlp6FfBprj8A8Esircd8n0ooBZdE40IuPRtD
2dPmfKn28ynu2HgDJxviAb9au9ddLzderR5/XBI0GP19mi01OkN1v+ytVawZ55t+MX7FPgvbxrqb
p6RIhusoFXk/JXRplvKlgT5/Bh946Wt39VVdaVabiMmesujCq/cqEnsGvA7Cw4cEOdef9HBlJVEF
Ar8xmiw/gppg+KxthToXRGccv3tXXFsJOTYPpG5O3Shga1qo/vQr2zxLQ7u0+XgaW6gltuIE616E
T6iFeyqvbnSMWnwdEYDpwxg/0z1n70EiaKb3xUCcRFfPXwjC0kqi9c+xFJMO8i1dDeTGQ2BdMV+F
9NB6xqcon1mPuT3ROOoWmGx1QESNN+Qysqo4GHrMzSDSd/wn1h4sCXkWdmMwQxceuMD0teOzLDmH
wtYT5eVQ0CqMxS4rm4xQbFKAcRaErqIeMvtNs517bFCC5Xp+uBMDxYSnLGcj0eB7kryXWFXXUAcq
ie3Vwfo7ZSKHMpJjA3pP6cJzlj1822pkj1pOukHAR/yHkjjIYBcSxLNRjCGksOsFLTQw6tZdOXPE
oofC9FrO3wV9cpaOuIpNTP62VVZoDnNE5Tp+BKf1KxBbOTniMnB5KIv++ep7etK7tPpp+pu1mnvX
Vi2f4sc9Z/pSwdlMCuU2hLOsasy4YZorNlXOreBlVrCcu1Nlqd65/Z/O5FsMA8Ly/C1imLqqWUyb
9GyY9f1G7oIdVovdj3sMtdk2TEsbWpsEu1Kgn2hDu4otFLfxbsA5/ZJDdfhWDSxYe5d0uTqcCau1
kad84vlbfyB3SQ55KqcDAbESwhIzh+aeVB//+IbW/gY/wFxxj8TMH4wog8ODCiYWd02JArp2fYYc
DC53afc2cxvYK4+7YLCFkH6C8wZD/pWPDZ3fEagdV3vFaDsD97YmXIleX6Ep0sSIhi1qntrJdILj
dV6CF29O8IkR2yThR8oiWoUUxqLt+ox/VP7+49J/M4Yd2jPWfEjfUWHqOMcwZdN7uFkOG9FErLAY
TArWiRjB8c57VYLF5k62CkQ0w3OVwoh6UfV7OhRNGhD80bCJUQo/VtZEG3rM4uOotYnbxyP/u03N
TlEvRB6e8haEXsKXVwK6xtShtozvjUx0OLk5Z1Zcq4yL4HKvYAgew84TNGh0u722yOmVDDW37YGs
IoJjbsNaZLn262nZXZct0yOd6XUVuR5CmNSv/SqGTFaKdQkqNoh2XxVUFipPwnG2utnxtP4hURdH
5pUQVvwhsv9Eer4XSJjGL4QXjbIFaB5Us/d0i5e4bWPxZg6Wu5Kd0WZbGDMOfgkcC6AD1/o/oUzd
WjAn2fJolf4TBmmQwnu2XOX5RIoRDEiRDefzUrjmc6Xp7KdTs2xvNEtHhxL4BOkbLH0A5fqrL9Bk
NMQLnYK1/OArUfEkEm7aWBgDSVeNRGvfIL6mYGgOrrmK73fDylNzCIWc4hIoC/TunPuJDMM2TOJ8
JqECyDZWOXrOfSLzhX3NJRdH74eAjJiPflU7T5dORw+zu3LnaugYPH7qIaobFLo9AmzVsYxEjvTB
xK3gi8TBonGiiC9RSHldIUrWm/igt1vI409mZZRyxz+cz29sF5sdOvi1TaK1oHosTJBWjR16nYjR
9syI8eX0jvyEXrbuG+iZhhreJU/VC/iSuACKqeo1xSFVl2N/Kax6ow9zPRL7OSRWkk1V6dodZ1ZK
gD909O+GvltsG0bl50uwKdNwLXH3r2e1F+IJ8IzEjrPcE+mcj3p23Sqgw4cE8C8UVL9J2H3wNssp
XvbYto+hXiaEHBnbYRe6iRvUAKyJk0wRJfu+LkoCZzq2flGep7Utau+HE5KNkjtL9kZnVXOGOQip
U0rceHRMJO4sTBbwA5I4WvRjI84Ty6DmMs/gzLN7Yz86ZGSXPfwzIz1ZZCuLLeaCOoUSp7+enNm0
tlIAHO/5IsPw1OGApnmPIx6TTcrq0wrF/PoUb8NbvJ6JZc4wIlAGXTB1BQJ5Rra3u5oM3FtUmpsC
GYhQnYKELEbq+DlM7O0JiLITcPkGXn+PeiS05aUmcaDZQsP2yaAm5YB156bBZ2OuSehN+0QdhVPP
Eytpt1wF0owYevBUeDBquk9y9ixwFEcraMJr3iUyE/zP+R+zwtC0LJnzjI+uQciL1lPXT1ETXIhT
xbg2PzpovB/jRQIGimRk/cFK7ZkamUy2nJRbtFhDJl/ZOLUPB0UTASkH/384aam+arKilinI7I7n
+sNn6QQDvRcT/GqI9Q7HZgp6ZjdXRcC7wLhXozd/GkBuwrYJ5QgsuOxXOKNcAcGFml5PHV+dex8v
JBJTpj/kbQE6/3MmWNHXIoXkdheTxUgVpEl2TIZu8acC2oYM/a07wwezxb3S9ldt2x/Pl2wR7SfJ
FVltFjhfpX8Ax7chUpQfzA+6AAOqqonWeV9SvlHubPK7uffXrXpmCcaPs0o5Z29hQ76CLsvwahwK
nhB5UNVlSa+/mfANWIan6euBgN/miAGN+W81sn2mL/LO2GCQhEjXwdlem8zD14L8fHpsJZaCwAYN
/jvr2yiW/vV5YNZX6ej7dQVpdh4wkJTTv0sbMOzxtGHCzKzefBIMhOeQPuA2uWRaQylEN+Ha0MC0
ctG1pvvT3S9n+zLvK+ZuxodfM2z0WCI816WQsAdP3d5C8FbpDjjg/DYg7KAt8347wvuQxW8ug3PB
iz+5WSps3ByVCkjK5OGHfAwTJBhMH+Zrj54tB3pDozWPgC2mgbvHkzwlid0rZAhKVAc587XgBhqt
w2DJKnAyP6gcvt2fTGjqhbvEX7XMdsgxboD5CMFtCedwleIGZ+bHF4WRECU7PUU4Wr9OsOilcg8K
bWcpqgtCIE4VUKxz1a+h8jt/JLgWiJZhb13ZfYol/7SpU8w8RvDkaC4MUsxNBMvGa74XaKEeXYf/
hoGNu5q+2/DjDT2Hxmr94TDQ9+iw3Qk0KDSjqiPVQ3vJnCiXV1sKL1cwAtHMW+DKQDL5rsYcf9zj
C6T0CQCSZj1ozqN8imzafNG9ucrB2qN3hzf8dQ2xNZvRcBoBd2zS6Oyvrh3f7W6avKTTWxn70UvO
P+9xV23tHZ7rdJ8JyPbQTI0IeYn2StzyvFU//JivVAKBDbG7LxKlTK4N2YPNFG7cigcfYDTFvhcN
/HgwAjXD/GkqezvkrDdj7SqKjy99OzHyhy41Y4xQQHM3PFIJF8GvPL6dC5DWMhw28HC9c2TwABC+
wTbRfwZ4KrjuB0M6l+jAtaPLzo3f2l/+WgSlCjC+UxLxS25QDljGIIb1JW3zBi/GvrVy8wb0RmTv
D4+0WmQ82aE9H+Bu0T641tuRUvK6qCxSr7gAvFxSHPbxtiH680bxKOd0oahV/hreY9xvhdAyFmBD
lL1sUaKEVMh2jJx7UwcXSZTnrCe/oYDVlwzNpu1zq21xOhEBtMh879Fyt45uYKbifS8mITfqcXGa
AmZnJYdz4A5HO/c6Lvkur8En/ZX3O8hg9doiVhBbl/DWEmZOdxjCcLBLaKCgRzU2p8PRvbcVih74
q2pjmPik4/ovyMH7R8m0NwSD3axIDWA5iJD1L0R6ICd9vY4iyBIObMSJu2L7jLN6qBoW0Ap7DQdW
l8D/p3BUZGehR2PPnuCV1fAWtqPgr0RNkpio5bHp+g0Qn4yBUTSE5ANTCiLbkdluQfXWVQZyF1nT
xN2n8QAsr7sIafwU84Kaerm9pjPwmx8oIIPe1DVQuRMx9PorbHKMN/srrhxXSL/aXrVBXEnry6LB
tyb018Gc8b54aa687a5KY26qhmGzsxTWcvqC4XQAus2vHYQt0Jr9M8BGpMR/b86XYkKFNnj/Y1ro
tLxZkAmTdT4Ye7SRlSuSpc4n5lGIak8o8cad4uon68X2klqocs7B5lPHmwWGGbToo7zcpHeKfJ1b
/jR/apidEH7JqE2ycQEQUue3EJyTVOS5HiHWcRC3bsCKQnwEDVrfiTazahu8tlpNEV9orQHS2T7k
Qrt+U5LiSS7iQfYVHmI5mvaGkJrohj3czGLthiTATlWaFR8vMBITJmOxM1B7ybCqNoNaf9Ez9CEU
tfzefzZdUd1+DlCLJNrSaZNcUgZYahC2Po/83heNtcouTQkhvQFXDC/NiohWawz+HWTZRnjRye3x
B83ff74PrGvAMnyFqXCBp/tDNLRgFmQX5rAqYyNAHwMwFC+a9sh2jSfGfgbOBIlzh1+Tc/C6/HbZ
HZH4QTD0eiAMvImPeZUDaXq4WGlA6UkWHRVWTJWTgp4pHxbra2zcxO0mNXfgBBfsMTKObZJS5fF4
AsWaqT3AM4JNT8DJtTJDAzmK7ncjFR81NtOY6GEUpX2BRjq9FEpQ5jdHnbedOs7ZjON9nulprXSU
q9HCYns4XMn6USymm8IK9PAm2vULyTpp7OeCdvAm6vhSfuNTCiNw6bcwOt8hEg0bFeuTdqQHQ8SB
zSurOvieeHFVrcdeVja2oIu/6p1ZpL5g6Mtmy8kjs/edqMME2aqUxOsnpFQsYYbpvjWxhW9aBk14
Imy0Q3iQS/oXAUauSlXR1Q3UM9tV1y97g+7fNGR3WKnyjwfaCLJ2c0Okm5tKcqwhPhK+1bIEvkhi
X9qXWaqaZoUA0+JIZzg5BhxMxb6k6sLbqL2fhU6XJD6u68JqNzbyWd2zWbSnZeqbuRaFZwATuYRm
9s/FqGGOT1iN5+v3YzyTbcxlnsg2UF1z0HZ4dfx6TNJTjEhqwI4VjH5oflNNSBk0rhz7nTgtoQXY
+vmCuR34IN+eu38dRXPbTYZXnDV9+UXbhTTP26jt1alYrmdObig6pX9cTgGTxiWyaBnP7NUbmuMw
WH3ejpIQJpfCMn3lV5AdP4kI8MqBycJmdhKeyxkkffp5KySB5fu6RqG1Xqn48uTqt0oH6gW7QZVh
Bu2xA0QejWBpdErX4VHHUA3OAWprteC1a5GH4TAZZIKbYLXCk/a/M8g6RAURGb0jfT40qPZ0vpCU
gdwa2PmBHV9a/bvJIBduWh1lsFNUaBqgRHeTC4jaaXDwcj8jBSmUwU/61qLnYsC59+K38WssMTRv
pcA1UsUoRcH9h+UKuYF6muai90Fj4F4uCyoQcq0mdGtP21F++/DS3YUlR5Uy4UXekDzqmKKYOzk7
VWvw1M8Wtxqk1imScsINnZ8mVQKfeUnNtWXqnWbx30dtxe0LwrCgJbDjxjoCWDkCJ0DR9k/VotOd
uuVfbWO2q5hRFzXkKKEI5qkKDxU0lILtrLu+3rltiR0fYQ9azUq9nIoQxGSER0gn9zyqzbHWeGKY
CdAQLzAzqtalfRvc8KZYQkszJ7pmMr80qW1RZ0bUJeJ1hKyaAem9PG2ciyPhaD1UGqCSwTSnkVLR
RT3o9ALOo58bHRHEGAoVfDdZYTE8XDYHn17j04p3dJR6dUArPdPo4i/qAfxu1iB3qThJrgDWBjhv
/DN/dIB+o+Jd1nx1rs3eM0KYCrGsEkNOMtCdTRpxyt5aw9MRBiaBJUFrtLiuNcqEEVtvUA8a+DWr
nWgE5hoUei9aCTsEosvAlcW3EVaLpv9m5l/MQiMCRR4SYkfSxs2+1WX0g6ZvJhuY8gTa+cP/5CjX
r58vST6oudk5CPVeahZpeUKJsHxi7bEgMPzOZiUCvzmjBY2qpVmX4P0VzZpT5r74xpGOwyc4csxH
T/z1ByZl0x70uiWE70Wy+KyXs8DxZIjuNa/JUDXWOonh6XeucVN2Z1XH7D6TtWzSy+ym0xNTnRPC
zCmTmFHYOVwA+2TGnNMbe5NxLI+u6XI2RR9/UiHNGnTV3lvghaZyStfNtn1KHEiyUwtLI1vmoIEj
k04eElLfs/ShQTsi+2Ci7mSWRYrGd38Vl4LHJmdRP3Ts+MwrtQqquhoZKkwvmM2t3CnZxuWZO86Q
qgF6ESvO+5hwsG7C9f9mbUdp61fKZ3rRl7Vfq1lgb4oS7i1426bwNqN+fHqG3tRoZOemnLBuFTAV
P3pBv1NGhYCdPfPAjN8Iv7M2m0OBjfVgrZbXWG9bUWSEUkAdaq5PzZSfViy4d2thUGOexBYIvi1s
czi2U6Z/m9H+FVwaRXwIWdIVxADkp3hrtlQvValwUp6CJqFQOOYoQbstMDkR4rqb5htW4HLLPCNJ
APK265uOK8mW4lfxJUcopj8uK1OeOe76uoC46uCUdGJ5coO0lu1bO2UpONiQLIrKZAduXUBBuDXi
sTuzdnF+9Uj6EXPq6rAQ6UmOHh0+axKapit9fI9CHV9XwzILhWzDHx9VT/WonyCE+145lWxKiSUj
twQGlvOpgISNHFQVzVlUUf1n9ANPITvN4enWMfPLLbj3OY5yc1VXytUrJCFYtf9kfVcUY0hP5xvQ
5kkgCfG2XzIMYZ5i9J7mSDdYGFdXDNXyqMBhvKeKw0I8zsuvAo+di2zKVt10VSTL+FymvgMLq5E2
IrmQVEPKo/cnrvfDQMQ8D8owXsA50XyCLwnQTBQIRaI1NO7amwihJNtH2cu54NO9pMXwO/x1USzW
4+52kpnL/FGYOY9R8ecPGz6/z+0kaQjsnXAJEgEkjGcdX/q5hPsMDXorQr1yOPX0u4jpUy80PS6E
8jkcRy0dHtRl28hHKU0QStYdYu0R23zgnYKEZ71/52kw8EYfW9+chB6eXgB/eBztXuecWhTZUpyK
2SdQ3r+75j7ePEVpegEMoI/Xrmk7leoCAEq7KfWf/QoTBi/3qIuWUI6w9ZsqoOKt/QVW2GxEN4wl
QWoS3k3lFHJ/mjeDzN0vsvTNQw3ZwiST0FrQ0PfdJgAfCeqkyqRdAKkTfS9s2apyY6GnWUbc8mRH
Zsb93nj/ZLjMJ0RiEP/psx7cWj2c0TMvee/izfi9vLg5MCg07nl9bt9UfLvVJ6KyP3uS70X2Ws9S
tnkda3NG5bDmLG3qbBaXoUa5OTjMpXPYNn3snFZePhOOCUC+xzalpjNeiUGpSIcLPa1dBAex0Za1
BMUXE3fFQ4MSi0XTw2i7L4QYOuMxvqH63w8yVwpjXZ86MbKz7DzXhfoJpvzSEiMFHADp5/3sY+1I
nwYHC96kwIJnsyE842jGLUJLRlWKO0v+pEcXz2PeiUGbQDLvqI8buLpIJ8x9wbpVqZ9goTri1waf
nZ1I3j+tfEORU90GxPI/HESdxQRrD3SdGkYDdoiniBnBwiSKtoQo0Lm8xZ7H/fenh6/WGRBQoAUg
3ihsmwgV6zkEjxmJKCk1pf5Jd3Fm004nTr9B3jAsn+vGPnYAG5UldwqPIgWrWmeeAdvNMQxysk+X
2QoH2UieAKSlWz8aguj9ehbEU3zmpKWsdzEEYovIlZZg4b0sJNQSNAxKwdzB70cW2ABnSzJtZwq0
VaxProlUNe2UHfpElkrzgH+cPo0dmKDmUcnJmPQKLCb7Bms3UAzPyND7gJfoVQy3ffx+TbfTmYa7
+I2GhrMd/GmGkwjzpqwQ0/EtRnTuxr1a8BC2ycNWMQ9pI8wf+KLu7ILHjOFOlU/FpQ4oRYn31YHQ
JreLscVExK4LLFl+eCVT3JpvfppKx1rSjIe+6oD6Ywx6DLdG8IyNevyppNNMuncmzRkQmq9R1MG7
e8/Cv/Tz/VEOdHVGJ05SqFcF4Ik73kRfDSqLI/DYFlwI6I4KaLoXq1DmOGOdT2wZIz+GNERCRrSD
ggqJ0Whac8F6MM4B+jGU5mf2owQf4t8y9865cSsmq6jek1FhOgSfjDeYqlAqRjcvTBBTJUdp8KZR
uJC7U7VK7geSu5TBmUKDxN3LLqtI2pTDHNSie3xQ/qa8UOmUVy9Y36MD7fuecND1Cno2iYUrC4tN
PKNBKeOykbMu8XZvvuJE2fJ3OqOWuBDxxFJDYNpF/CHis4Bo2LaKkG3hlTArksBFoxNXGTR39FWk
jshBxNf/wv3mgQ2nVf7e1KwoxHlCPqAJM91i+jpsyYDOpHDz8l7cyCkfTQd+uli3jghlDIWFsn6z
v6zmgLzsY6uTZLqQCdZtDoNcYPA73qLyyLZ/7P6qiLWLeOJjO1JJc/Wau0u7eXLVx0QVp+yzEsl9
Xy833EJgwpRu+AAP6gMpO7joDyBZJmGCQ9WbpLaEVd6wmlbNLL4p+fJpPL9IT4IyKdUXR/uh3N/D
t0bDHNM+X8mBZ4HCaY642bAJLMsgfVeYFMFSuOMkROpeG/aA5mp4zHwc3+PvN4/jPgTPOKIIxqa8
v9zGZNIVPX/42/V26XPrN7/f/A1CmqH8oYY45h6xCJavtk78hConwxKk7tp5YauKG7LT4QVj6qWQ
UERHvaq/+NRlCdVNnodpjF6u8bRa+ltRF+lA+SkQm+Uu6wWSinxB5Ntk9yZV0Vunq3UN8uUdwRoy
jW15w/0Cachd60TDPVLDh+U4Zw37uwCFWjG8NFJL2rCJ22iEmls5H8ySA7bEBlGjJUp36N9KvkUl
h5W/mbzCBR2IJ3QFkaSPC3g0+eD8ojwLayxTbuhNsz/FG+kTNDNA2wGbGgM2LKSnGbmbsUg/bGVF
tw4yNyLAb3delWgpznAHCyhPjT2V8X5s/KDAHrHwplOmM/pZdl8orACQT7pD3Fh1CPP+f0gMGokq
zKCiBA5VA4ePmipZ8E9yPCNTdn4XmZuoUbzr39VLXVoZQVh6MKdbKl/4uo5OT1rOzFU8KEnMnxWk
Hi8RucsqtqfzuTJ+0tHcFNAzaA6fJ4HCbKnW17Sg7lGfIeQ0MO8/+nK9Hdkw0LZ6i9JtugQM/hi3
t4YDiklrUVaIkM5BXjFW6j0ngKvrPApxfkhVOBHCeDqQErx5jPM87Yjcel3osjc3mhJTaL1Cx1Ee
k2qF/7jO+OA4Cp1H+ojLSl77uRiIvGF/gp/60lbw0GyMzTlblyj0oZIxUzPs20ncEuAPLHaT+PES
YlcWeieEkc98//p7Hh6Imx0EeQ+gHFo6thPLP7R0SuFEFx8n5WPuQx917feu/bGoxFMfyX2IhSnF
idiiRtDVggR2vvU3IiWWiBnzoXVN9vavqgtnZhG1VBVHfEXcdw+jTuGFX8tUhLF59yBdWNJ0lAUW
jQfM0xqbR1x7gaHIvZZBFpdXjtbrEj/M5wFEuRislrTMM8N8XDQYaWSmQOnT2b+n1Bl5CFcvq7T6
ceJ98tZOjpiLpLBOS92nr8RRwWHv7P4VLUNVXbvCBdWcdrWIFjpEUbJlI3T0xBfAqNcOkqO1hNZZ
PYtI0NYOv2ktbxX6FBQ5M3DsFsiWU819YjnOdKni7Wqt+IV0b7mv8ENa465cNElM3kk6hXDUY/do
jdmG1F6ALfnZUUtR8ecGABDRiXyoOmAQ/PkCqTuhkHAt3w2Q/NJ8yXB/Tn7aR9br7gFX31U5d7AZ
sgi6+eI0RZ9mHfnSYfhGJBMliggaSOHEBZDqtrHn1Wd9DrDqsiTvk/99dKwcSzCsV7WQkEY2mKXQ
oOYOuftjAe1O9cAnpqJy+KuS6ko2yJneRuFHmccb0GwU1dw0Cz19Gyjs6mISerVjL5oHltEbqCvq
NfLWIvvPzNp62oZgXodQjFRIw9Q/lchNEW7n5EFEtmM+uXafuHua5BI7bQdPiZnyauT0xztwvass
6639Ys7GqMsnZFDNmKb/Gb3Clxz9gmYoCK8kqS82EsJyckrs7gYUCwGHnHroA1+CsOvIAps+hK3x
tQSgb01ZQExy900DY4dHHE9LfPXFoCHDRVmqP5SdU/Uzk0pXAjMQ/5y1c1ERybRpDwbATxS58iIf
ocRJh5iPUJCAkyCAEUU3ndcGS8y96aMOvHHtlZHPTN1WIiIL1irx7wt888Hf9l/kgSe2bYMZSyXY
B3K9YU0ZuVxs/qWp5XCRDwD48YMRij54k/gWtXn8otDPcwaWhb4hwHLrfxtNcgFsFtquuB08tXCq
82jm+mQ1BmDgeBpimIA+O0MrRvPXdiZiA5JQ9hXPc3VnqP7HiYsSE5auHgkKqooosRZ/B1w/XFT/
nIwBjPqYzk10ZrDuPc/LufZEMeYYT4qOMO+y2/IbyXl16jz97gWTZHkdBtTwMWtX9jb75dAsGTyA
a++Qh+rkbFek9q0gbK6tfmJClGnJQbs5E9b8qqLIcWIVnF1zUQ5ReEFlMx9mgoYZSAK2twISST0g
25d7chA1giyRk1jcpUHwzDDP5elDlZE7w/asYdKvfhfloNbMfn6MZECfr1Stu/TCc8Bol9JO6V7w
t4fB2qq4bc1ARg7rI6jFB1pqKmnYiFpfTSI/GwqkwGLDWgiYyDwNj5k2qBkBd2UE90RD0O9hsqiz
Ej4W20Iwsk/sX2u87K77oO0LznMvBithk5FBQJB6aYujo7p617KGt7OgiFXajYSLqMfFgLHT8Yb6
uqTgppOwzSetG4wOfTaElA63UItZ4Kya3Ov9dbe0/cC3EwZJmtx2gIbm6RPa6qqQIhXENE1m24z9
UppduVrh39Gm5VRRU5vnQq9mhXzfBDqsG3XTJx5b6yK+m1WI/EV643VLyEBlzF2rDohcGQSgznTu
PkoqrWWAJakBn+2LqO7GuQCiCxvcgryAx+EKz8T+ZK/Tfv4VJXkAIWI50aDZHwcAR+Bjc+8QnSRR
oV7Af+0e7ZUTAUqLy+EsORsrFo4VvSsTzzRVCoSX1ARTeajtEFzCqr99IOTq9PuxenE36VWWp2Nh
3h9L0TN9QI2ieKz6MYLSKnmnkXTJ1DrMqmo6t01C3iOfYjDSDzUI5UrXV7SYnflIxDUJW2QV6g8k
UJYeQ4+rKcYFNo5mnreD+auKa/KTUfXIqwt6w5BXxZ+2B7pZk8yftvZIFvLc5W60pyPaPeVRc/GP
P/nfC8hswXfEK8r8UWFopsIJbjTvqv/0ElcEhnExPPGcU8eF5lLVMt2kg5QqOd2XAa1P6qRLfZcC
mouZqvwP54X65RIFLBzGCXsXHn1oSHr0cA3l+vnnN4zGdEONWgwARH2y2rUyc1bBxdAFs9yK41C9
Lxa/pn5k5R/m8/QX6JseGvl+EWiPEh7N4Mvzs2Nb8XrE6atbKnVpOSBsuFbdhTNqZR7sKaH9DpeY
egFpHfEPcqPTsmmWahVqz0AKr1C6CNRgrV1hKVs1lwUo8k/0MmQcxilU0a/9DrZG4GkPuvcn5zA3
nShyl1I0UkUqwh4RBrzSolqfNFOlcsiBTjzQt8hfHc7hlvitIGolHR+TP+ATfYY6uP8jvXmqodIx
qSvntun6eibsGLWQpjZc6rg2t3nwOYM/Dl5WCP9qGLOHPmAvjzV9gAwXlzIF69oVcRZWnsTWUK/Z
16AnIYFZRh2cRoAvZBNup3ZlA/cuQGdwkM12UewJz2aXKDSFtPk5P48mKnFBIpcyYe30jxRubeg7
w+oXXuhk6BP1OSESxz8jdS5FG/U+fdRb4RcvmFU8oouDPwzCvw+6LSjhJbGLMu1UQJP9BS+jAVrt
gVK6eWi90potCT9LK/oOBZ9R7wubxCuCoaOwEsF8T2gVRg9Le6wcC3zemJLzUHmMw8xW4luc4QuN
QnPl67ym8s+OQKzQh/bkVjSXW3sJ0xRs6HRBtCQ31rdJLbnoi+2MRVy+HmVkRTIkewQ5IaLvqO1O
O0rjFvVezNC7rr/w2a3jvhImBnBxPxKyA+76fxaVHRXR87fr9weKo4Xi6gR+jh5dKriMHDio5mhQ
6+IS1mlQ/p34msk7/7zI4/mFjE+/RohLtmAiP9yNBdpd/kyUqeWVR0pBOMmE4NY9hGNQzTScF/mi
w0NfCWxgVEJafK/b/IAzhO6aASOyTe3u2G3xG+n9O19VIS5eK2u6kzJDXm5MqfLCc/B6uGpNPmKs
KsSh0Mat/6gqH1PA/ABM108LQ9vy5RmuaAFKHaBIwUdoBUYWExDxyMaH7zDDtEYfeuXcPBdZ/V5i
mVkOYh+PLI4V3IIaXCcoO2Mhho3oAdRI5hh0Tk2pclKdRpQ5C8TsC3v/le4MQKZzRzdpMp4Xew2z
SD7c3R3X5pWTHyPwmok0aipJYklK2zIO9hzUecn8pWDAZMueMk2Petp8LbphZVlzcgBClK80qOvF
94s+6xx9LRijjVUe3zgvyoLDxds5mV+gD9nm/xtxGeKNGo7XURLzdHotpukopTwVIAUtijeqep5+
G03goMd/TdHFR8Ctn9vN5o0WG2j9TP2flZ1se5fY++gNilqgBKFHvraOHlw+bQPNyh0QGB+EClDI
855BDrcCMRMjRjhpZ2pl42G6+WqWmxLbzV3ybfs2YPdTBMHtiNhWESUFTfzOZmvAanHZVfC/ebHw
gAdLg+pzG/Ffvb6ySbfogspO2EvhiJwQ8BmMIFtZe9ufRiukHUb11Ozq2U8EJFyYlPKk9qlhV9tV
GdXy50cxAfjlKU6tiAMDf7aDK4nlzdsYYM94jlAkXaM9V3e5pyKQ4K7cG5AiOhcCY9Djvge2ROtb
xp9wCNPlndK4u6YEQ2DEY9wvw1ITwiK/xE35/f7rgX34+rpEVlArWATQpqt6mLxa0UJxGKO4htnb
x7rjLeoID0yi13iPChqDyKd2UcZjY+YVVqGOS+GuW642QGsOGlMKZopSjNWqXlnLCPR7k+i2i5yK
5OIi2K1FGtLbiRqexZsuR+NnAIZBguvmE9PaVjCSOz41ZOr2bRTIQkkjWb84quJZmjWGQTZPe40t
dx13v3sU+B8ZH+2lOfzTfAg5BqZJpBenTOFVd0QwVWBW63uz5XuKwRbQDNwcZv0HIcj8cVRqN9zV
zvLNfoo6A8NQL9Au5g/migCCornRFQiue6ziUz9IqRshETvCSU0hT9KvoxexFIYwbq/BXJ9WxVTk
STnNwkeoXWAuMGXxI3fG3eKtbXQ6Bjj6ZQQjLtV/DDGa+BNzV/2bmjjgj/Q1ZDUJjQblfrGdRN3H
+w5Cu4H//fziHSMzK84x1X4Z5BlgtPIK+BJXov6xuykA4rqIZhEKjWspslC3PKdv/rSqZrHarzLS
LPZF+Gd35i8DLABA2hl+ox+q7tht/fuhvSD5gf6dtSGib2uq4iS4RC7MAf5jiz5OLLWfPG/Kpxak
fJUz6/fTGK24PE6tV3u1UqwAtHKafzDK5suzviejM6cHXG/fR6jcSyBH9jGujH4OqBSZbBIeBJs0
2TheF3kg4JR4p3618eQiNkuiE2OCFUXOLTUIwtk4fBgx4TI6xAzWyPQnOox6H8hjgH04SfTXxfY2
qeNL1rY8CHFn++c86yO+84SdbTnTM3V+HdWWffZk38c0ith5imCY+gvYHbLTDdGJKQt3ZBNnIssb
cHb5Kd9+H22YFZFPLS1fe6qto0RnmThPAG/Z95e+gueK8ZKTkAwvOey3GuIOETyURWfE5Tfoxgm9
aKWShoAhl6zEpOedaIcCUMh4mQcUCqKukglbtsBNXDq41yswlNFJOrq9kJxPfuoxZ99CrIxdhQg5
YA09UPnaf+jLsMYa1UZtH/K47HS+ZE04HUKRmcusqQ1qwP3v885JKAVrgpa1sUfSWjShMq6sXuQ1
Ix/Mo4xpOF5pEHggM/m7HLKRwI8u4x1i7ZZTo6FUiOBpguSG/ju9esW6ZhfqKbi/iWbdtqib1Lsu
sny17/I+F1xfc7SBwqqXTBZEv3zkGuuSwo80gVJhAPSjOGEriNGE+oA1y70XQuQVi2Mq6hwYWeBY
aOgjZAXp2fPf6Sb2R3zoUVsSO34rzN1kuHbH0hVbtc9d1AyBF8qtEuz9wMiR/HHhA32IKOEiZgoW
QnRsx1nYO68prLt1jy6OGJ1ErbXSperZ+TR815YP76gRAGZBhJnMyejoY27gwRwuxASUKwE6G0mg
e2Z5TV8+21k9zbWPaiYR78MLz4jLNXgskTLyd8WGE7xElUZ6cx244WlHBMSa6r9jzHLFiPHhAbML
7fp0MOB6w7a3EcNoMuPSIz3wbgYVzaGXkDz/sxT77xzjJ4eRCcov7np5wk4A75GvV1X74/483Oaj
21nRQFJBbd+sNkaGdqxi/wCKhnglCAYews1nHct01HuPB4oSBiJfKJO0wqPs98HoN96335b8n9VE
SbUx0y3HSG+7UvhKKXiCVac+famlJ2mYeA7LE1Zoav1YKDl19/PVK7xSVZnackr4xmK3j+kySmoc
0L5g7+9GFA53Mx2HEE7RG4we1PjgbnYMBYB+THSMlMGOT1t4F4orvgxEF9SWqYaod8RU0r/CvWvH
PY9W+Fw2g6ZqcTjDfLsqwVpMyAkiFt08UIw5OxO8AqRtMNRADdHobQRkRM0JVmVE8iRQojPfQe7q
/3F6MtXfzZvupsoN24bYzwHAFwAq3wZDLYvvseBNIkvX1vSpuESvETfoKJ4T1NZ79hQwusePHzBr
PQviCGtmA+z+4cHJF8gVkmo5efKlQ+7DYPsqqjbdIEkilbLliTSpbKdsl8ZwvSKuXLm0LED/plgA
RrkuUiqYCDVpxy0xqSNiUMv4RKXehzERkxIa3BGxORLd8HWEtyLZWXSM8jTlq+xz/FuKTsp2DMZt
iPePb7dxTlZGolSPUkYCu183EAKlaPOvAuqmntQFjcNeQjcMtEy+Cs3C5SvMPtkdtC+ygk7tI5fE
vW3Jt31OtdNkAOXA6WhYc8GXbYMxAXel0Gqo/y6T5iSd1hUhLbjsUzA88dwXeAQjfl6AE4XaU2ai
n4Blaj9+D3wN3KKrhof7udlglemgSQXwOfgpgaPjT8WVcFgPZJ1uy4QXSthRsW6jwVhe30FD5282
SAmRIJ0T1gMUFF3ZTm2SRNqYwbEX5yXW4WwN6eI9c3HmOf85XL1kLwUjimp3Jr738c0Nh1VNUs27
U101sd3XG7qepUPnYbfKuyz6IrDLIUx5vElwJk4xaetc6OVelmZb148KY0GjmgSCTkWbRiS+XTwe
2deNjgzn1YjFQrn6ir82zXX5V+qVlo1jAvkfyUxvDqgDPnJHSiRrBX98BlxtLOOx4CCZBVTPtaUC
G1yaXtgWRG8LC4JHINfkIuuuQLQ0AhPZs6D8S99DXjd/Y7Yib/X1Pt28NE6Q6LWJev3+miO/LSMy
I22eTwiFTOt+YVcOsB+LFgF0PEhoavtg90fjT/1qBydPUn9Ni6WJrQrACyRguYW+kE+QWyMgo5dv
n3I8SOym8KNUmpMGGyBX/oNllSLo0DdGe/x5TsQn1fRq72M+tO9+WBkUn126xKv+fPNey3XCsRFV
u7yJK3wmToE9O1q5pmw6jKEhO7CnOeMXrevRBK0l/vt02gejOZKICN2pVvkGiOmjibfIcPSioLav
fHfob03z6DJkBB9zzVjI8pA9a/9Z0/nS3n1TmIwOmdGe9ARd0+HGDqXDQVg/MLCN85iYDGUpMc+D
MjrJInIARJ2JUWWOijQQz+ONLuGFlTRjUF9q5Kv3ixvlX+gBicCa1mPdVMtVpwHTtMPvlGQvYkfo
sKGllmvW8lT2llPrAlASKKLexgQcbTFZk0IRp9EDcOoTp2ZPjTEHWuDMrxIkhmC9ES/CTz0rWqE0
5WkJlaSOjO9iryxIHh7u38IqOFrAuVVaGlyxht0mhivOEjgyOq2TH4ZwR2xArrbojUZuM5iki+tT
KJzwJ3xHm6BD0hX/1yYapD7byGtBaMKX8xx6cmq4TVqtgmYS7ucqzpM3W72nx5AbZxDx40Y51W6o
7BtLbppCckn6hII/4kUewcJL6pVmQHujCH3TEXQb7UkQuLaVopFScIky/wWPAcKnDsa/jid5UFFX
wav7df2RvkRbnCGWcjBgIOVaQG5imQNC8NJ5m9na9YVXxSowBtmVyN6dJ2RQL0qRNgmuw0ycmdGf
q4xHM6TijwYDvTfSMTLMOoYUnRCxuwCYRTP8SyRv43dt0offe0fJsfjn3TYAFgDMzXauLhtOPDNE
RCkkBbyTig4ZM+bOQh5QYlV897A6ayK06g9YK5l/RQdodl888AvUC7PAhXI5yIu6rwukfmIRD0Dp
r9Mqmw3vyA53dreKoKWR9AIICyRKlX1G3+tnGE0l78A+y81rMJGqv++FqtwPIHno6SeognvrfDVo
No5p7HHQdz57XYEV8UHQ1KS6bvKgIHBncy/BNkjByr11mE6Yd3L2lb14KnlYQ8+Ab5Dle9FLyPsK
1W4cLE/hFQeKmu7ALesPUU7jMpUBn0avlQzKxvuQS8t3xRRK7fbKW8povOz/NoP9X1OMo99m+/yI
0qy7SinQpUqB7lISkBYCluDI/0sTJ8gLU4tXXANxgGAzUm7zUSlow+Tv3aBow9POQBmbyuIh9JXS
UvbihSNGYVM/sQ33LYu/cpjEmDWt2Ym59vIq1QDwPWc32psK0HGND7v1mDUx7Y4q1wZ8lokyXe61
ENJegCx2REHnNAK0Cq1gBTSJbf4ZXKlQkHUtCk4qApVlo+WzpzXj3g4xkoy3oTl6eHgob6IRODpj
nWnQGbsdIMSGiDmPgbeIcSnm9CuancbZBZwF+SYXISY5rP0AkW7smpeSpsyr79Irj+C1zeOEhfv9
pSSKpQ+9jTRRwFsKIHwCxbSsAvA8SbWqXyM3J8xfXjem80GIWtMtFyuPkkNh/jnFBdAfpVyMPKFU
+YoI30VLGYE166SmvK9Rvzdl/+KZHhsJEYBGbOXV5x3a0ranv0m+bkqymYo3Ar7h1jLz4Bm1XQJH
EkgcR2EoGnIcR0XZctX8omi+AeMtV0P22top57VOTQN73BL3+dWZ8iXka99d10gphgpHMHTyfRZC
FgEOhg9THWesTovUOko8xM66/6F5OduDxajhO2pXmI52MhkY5aKtzaFpnleRXjBJglpESyfmpFrU
uQdeguaAiMYV8AGQ7+hseXHMfjneVUBLQko1Nr6gF/IgPfSsm/AoS8iGiGXmdcaec+LXfCw9oqA/
a1FlHljd3ysbu2UWW4mjm9x97wclliNKu3NbrFqOLIYRJWAERXkEjc8hZcWQTNcZf/PdouGnMvr4
yMqSDnUhs+F3DxYBkfW8eI11SVDUDr07Z7KHZ/SHlShXVD805SeRBG9tg8rcU2ye82zWp5ESCLV5
MYuVXSXIg5ZPnAM3Qwub3/vgtuT4anQAvTWJtwOd6nm5x/JCrF+Dpxcw/OrFIivkh5U+YO1HTk5q
UPybyRLXGlktkYzcpC0McmWdi4CHt5/fUqM+KZHLWPIso1wckFSsnr0uE3+6cEi1uCcHFvCu9tOX
ypYThjlwlQz74mGPzizi7NMyHG//PJ71w2qXBq0KrbpHDPSeofbSgvqdSvJ5OvDuXqLts/EY0Sxp
uZoqFpTDeOyl2S9gCSs9cv6rpktfhScS3CDNIBbZ+YICmDyvV8NrBKR6OOtmxJx0vigcqdxMQwWz
FKBb6KgH0eH6DprkL5u1iqyd9DcygoBK/t33yHxPP5TQOewTbRkslWebcQ94qIGgkLJKzMUlL9iH
FO27F8dAckiPhayWaUNYGAbFK0rIiDm5nT+HZf27hd0eD3jLkNu2r//4RpUHJwudo9qf3xwZBrn6
wYxRLvY4x1PojXCkZ8dYIL0y51Tk3u3QRU6DyE9CQu495LcivcYwvR0KsNlCnMe6idpbJyrBnAa6
yXQY7Xr0X3LXMVCdPUuNKolOhUKl0ce8fMv0SfNa50cOvAvi8FNcZhVSxbxH1M5WBvKIFWIWvXnv
PqccjhnnNHMISZsBhFmkFlzdX4EzrGsZNqxY2KrFOcBAX8ZmIhP00DgsmNNirikj/ARSkLdE/3Hj
7vjQlb9KckCRbx2X0C2c7t17cDTyHA3drQGiV7oEVj1d3FR7TSIUf5GTh6Wc01ZcvZ6oZFyLkcth
WkRVRa22Dp6EpV8lIXOZvgwUt9/x7vdVWdtUA6F6nW5EmXl0pIXPoja+TEWm/0mXkg5ibEbPv7iw
WotXwEsEUYac32m0IKPNeQ8dx3pWFr918lOAL9cSt9AFFfzfG1zAwG/6SY67MKvw6AR+UCETif2g
JmQiG4zItS12Kc+EMs5otzOpBU5Zg0EBYtZdDN4fW5xu21AVzNsnMiNTC89NJAgk3BKVjF7sRaWb
oyoeILTn1+ok4AiA9PBD+6aVty8Si2NK5i733OUlPqW3wc+i2O1kxgUG39/5Y9hwu6hpBqYntj7m
G/XXY1Kau9vG6F+tUJwDWpH3FMrFokJhZ8DUZYYS8J9x4FYgZpIfhEUfUTKlbsERCi7Xot+6aS5d
WKUoSyqUOz34DDdRXkY4WPwuH68SMuW602iEaTJcGzysJVn6npSMJdyXKCsY+roGBU7SF0x2ptHy
0uhtzBb0OKLHscfjjdhTcgtErotyv+mvNXntVNKqGADJSXk+cURIMPKOyptZXgr2BgIS/xV65rW+
aXTNYQTN/kTdZZnzMvy9nQf2QT2FncjzflE5tn+kcofb++93agQ4/j5StjuhCi892U4WNZdypebM
sDEEQRELnsVykgtTLhEGIOzYziu6hP47S7G9mwCrAlbakaeh6XQxFbSwi9FRR9+8c72IJ8fLuW3S
5i+iU7XwXorw9YwIS5iQmM8XdsMkGs3AAUzMuJii/8kHAvYybOuKCzlacE4mqxog9uI0jjDrHhD1
+LLBK394jLTcPNFEzsmMPhyWnbknKlXFQp6PvAl8mFCYLUZAigcB9Dnf3rzwVCt7/bX/GPC1PFFm
dmuX+ggDYZlPqYj5f9oXSJwkoLJloNcht5Mk2gz0GSKnL2iFyYDTpKEEEO2sC+z2V11Ry3X29jtO
8cslMM14yb2QCs7HrrpOGSGpQKLgYs69GCF03nCYqCwSesDyvg1z3emKfxtX4Uh3IYTExt1uC0Bg
SSlKzksYJYz+ZHNWcjIpGQcZBlagMqBYT0udrX+TCeZWCMmV1nEUgkg1dWibkiddCn+UQYcEros+
rBkTj1oLNEIf2rIO6y8Wv/JvfOqsgHhPUYfwX5Ok+3oGRmn6Z+4RSmJe0O9fcJUhROjPrRvG1X4T
mxRyNerPGhuKRDk9+8P9X3C1e0o/RSpokwN0PwLXEq/v4I9fEqLreZSabvZY9aBD0IP6E66lFAzd
JECC27X+5JB0OkhjE9IguXhMfJ/dLoB0FoWK4e2FKwmR1hg02Fz9of1Hkt+BUdmZvDUZqvdHfGo1
sgGaF0S+7RPEuosTtTCb7piZO8ZDJ+RbBMVd0/cW5GeN7sKHKVQw5o0yIWPes1Cxj1FmNtwD8pIX
TQ8y3rGavX5lW4DI9GkgdchjzcILzXuoE07HOE+ftKSvE8xES4CvshTh4X1rFRn8o4o22qKzP901
8vyH7GsNFXQnIoPM/4OiPq4yr7rdvR6EMwljXESa9cA9DqqpLhZOVK1TPc54K/dQ0xv5Vyk+nuRa
BAXWkhhNDMkaNmvUQ8GH61NnpOdyaKwOGl2cFan0gZ6fy+UnIDXFS7O3E1W22/Y8ZFl7IET1Qmgs
wI/qOSrSFhQQRo91h5UKuayZ/QkppMoHtL7FvNI73NY42wuccHEjNweVL1qmVo01CE+NKBgmZ2km
njDgnrecEz7LFD/EG37STy5RwWJrJO2JSRt8XNsQFBmj073wdf2n7MvXQIaDXPIWDPdMxKj7SIVm
8uh9/70AMFvkvEzq2SIs4CE/csHE78bbaZibv72Nc/GrihqFBBrrkbZsvOutpMpNEKgH05Um6z1s
lml78WMzBg6Mrd4UIfEsq46pdLLhhphoqnQQPGNJjog0KvrYIKYAqG2tS6xYrGO5UiGOc5JWOSJl
QeYaHMPBX5xERR1ZcPQEMbXUijD4TpGq1LaOrrynRhMhXNlDX2loFfUvcWuGtMP2VVUuZ+7XnC5Q
X00LWgfkznrfGD8sy4bIaFtdBbEZMzE028ZbkzUcmqn3hjE2lTi9s/is+93F5E3hhwpTZy1iPJIS
5/rKqqGq+9PXc57awFZglbHJ2MZbm60RT2phhgPhoTAiASiO1J1P18sV4bGqEnhIq8p/eCySQCSw
LQp+shJz95aJOdcb55Vyxx/wauePOzLLEVNa98kWjHUCs3AY/Pdt99EvjOJGIoIqorQ7DEH8jOYd
yhQm6vHPM/sQUju42C37buIcr0HoXEv+V8BQ6LItMWuwXKtgjIfYgJ8/3ovXJUfLwNg7BM0g8bRI
nuLFoXfhLzlHxVU/U9SnB4e3cdt5EIgAv+GcpxO3e9mlL5GCe2to2PGX5jbG7B3fd5/JJUs/S/2u
fhicorouujvFVdzgD347UEETcFEhDWJiai1O7ke/zcwN7xwncIe2dCRTfGy/HIjFhAv5bvZV79hA
QT/yiQco+vxwSveahS+IWGn6dAS2Bw7qvt3Hl+cXI/MzEEECykKGEPE+BwAnsiqErnm4fnk9YphQ
Y8DE9oaStEckKnWA7uemTUz/w9HDyVjl1+gTSP9taSd4OAf5oLpd/i/Xx9+govVt2zrSb21IgYeV
ky2RARO/a3gUWlnuxe6fMYs0lmNppu9M+SJiiiMWVa6vtmfH+4NiCSdeoLD5R+PAAdFDrIrS/vxn
pyi3N2wDkHqeIyPf6CfuvBvVM/oXWXcexXF8mhTAPot3OwcUmc0LshfpgJqfZnBQEkUiabwir1qT
dnUQNPkB1qeBUgfvy8hFk3vT/IsA4OEsle5ZyWpbdNrTtAVYXWKnNelPYV3vsz0zlU+pfpGOrIYO
sCVbrThfzqyIYmMdgjY+gX34BgKnXY7iwrqIRMtsFw6EbqxZZZL87IZH9yTXJoHfQ3vgwfTb7gQP
lqoRZv6WOZRMNAdXEYx+Q+nD+kJSOzTfClzbuSgCjIxz/z1Xt0aPIgl10g1/bfrGWHpr2/43SN3G
ReKxBUtP7HEJfsOFw5XDW78O0PtnVVu/2KJXXQRrMXDW+tTmNuds2CGjvL1HkZ69u8AvzwQ/qxfq
YSNkFNNCnotKk6BTwcpjp4z6KD3c7GDj+O/+jNaaEhDgbely+kmJ9vZ5FA7ikGFmKglO38nbtZyZ
qPmh+NoUkBXFU+4ykMDMGQ3GcDI+yLN68ReEi4xL2lIM/Bt0kMc3F2VfTaaX3tsoy+cZNPZxiV4b
XrOIo8qJCqLRbSGqMXXy3cQBKjLgrpx3JDVC5wa58JcdNEmUjAGaP/PtiI8vj/zGaK2ZejwJF1bj
bRQbbAJIqETtHpSGgKKhm2kuh8L7RAjF62Kc0pYul6QYefwjuDCcqzQLWirxl3akwYxpbp2tTwTj
Gg7RBkdZb4o+RIvNcgiSBbHUfMgm5T2wQlCY2uxvjDOJI4uIs7HhUPFVRhzoYBzK+cp9O2vJz46d
4GZzih1Zu00kVELQ0v08d30QjvggzAVB7Xi4zCBRogZaQNdFSpJd4a+tZgDc+uU5L30rMVAqS8hd
NsM2VBPrLYWEtW2hP3TNLVNtmktbAnlNlhT+Aw06/ZnnoozWOlPCM6tqyUM7E3hYxiJiHV4P+wsp
GWSiv/Y3T1Db1agJi6vHsgxregt3aQLHmTE+iF+amIGa2FvEFQzD3WIERjykqn7srtBBtKqGPzaC
wNc0lsSbuS8iER6ixVsmPmPEUqGzxFhisgv/YrKcabBfANQkV/CH8oYLJqGPzptECTWDD8l4uBGz
zYvCv3QSWKMMhOCqqiMDgUoZlKRje7cYLpB3Yx8sDPrNzKKGlMGaCqO8Lq+6stuTT51wz2U0jXlr
xxelSXM7gn8nvxXmbWArvtXj9Viiz8+5wozC1/1BB+T2B3QfCsgcmijnrikmJfSJH/1p/E56vuIR
knZ0fn0XvJCAToqtmoU0KmxVeFp449bIBNUYHmGDlGHANHn3n3mLvuTeMnI+Ia73UDgs4TwrMbue
QSxSU7t/Wdk35Wurl4BmKEmD+dHNBv4h8Jyf5h5ODsiWMZDbRIfvnTEo0ImwGUQmRSWAbEdLkuJU
xgejAlIHYlIaLzLp17ab+pVbVm0s+aVfEsCa0Savj1rbIFY7Vn3NFJjnlMJYrgKx0GmdRZ9zZmMB
ZwIUAhN/r+a7cyByioBVucieffJwAi+DohEqo0ZCEWj6rD7BMTz2OWW/u3dVXz33WabS0jW3vT4X
PPH3GAKa0GgOKc08SdWaMbG+eBMwToMmDeY+ShQTwZa6G57qjIRz2tlZApqIBG3Gd3uwz30oclHx
xEQBLN8dIyYzSCPP8i9PLMP47QpSInVUJ4PLd484YFwkPESo6vztmF9SYucqg4gC06UZ7Qih6ohp
2977MXPx7rmTitiYWBNdmKW3FxrO7pD0QkH4kT8k+zqiChT8ushNp674tCVC6yevYUrocWqqhlay
DDEnutd7wcQNZa+SURUhXPpuN+VPnpZTVF1v+JfyhMsopCifPmpNCgwDf4tO+GJEHN8aU3HTW2fj
kWOU4pS+dfmGb/KSa1ILY2PYECbkRyaTDxrO1uZMHxhi8pm7ZSAApZOpoC65feYBqSxsHDkvJD3/
QYdD0B1+8OZwRQ+08/YYDflzYK+KE4qYx+pf8U6Pe9c1uiWv1+3rsRSeAfcFFSRABUsBPymn2lMz
C/Pbbcp+K6ZXX91bXpjzRaHDDTdmpiIY0PLBJIfrFGnT+0tB1//RmmmOb7dfdJSFjJNtv5s9ELhJ
lCNnimXa6IgmxCaYZdq5p2yZkh91zbk1Hfc4LlPHpLXlprI7DCokpTopJi2oYg0nKTZwXo7LSKjp
FZ18gTH5i28qyupvG6QrPB1TDMM6ZGFaNsFBK/4hv7nXbmSjqvNDetJUVZ3THyZh7rf84ct0tgJQ
57ihbkMKE8BK6K27ydFQQ+T7qjhsu47noBI7kqSroYfPtfZps8ZtgGoYUrIgtUr59bJQxJ54DP1W
tUveAslX/Z6J01cF80kt+nxTj5xgEC8NuhscdrVkrG/ongm9Ui9XnFC/oYwC3qAFmYinoTUm4tov
HOG/94tnOCy0Oy11K/pYpiFMXJz6DCqsaozo/vbUfIvSJB9zdubmNzeScG/KEYYHc+BL28EpEn1d
fxKkahyY4EYvQFfns2F6QZ2NEF4w7cI30I61JHQH4mGoOm/PKOmDp8sbCQmbuA2zo3iefH8DtRUY
EFHYGr2pQ0JGvEo7NNSSmrDED3IUgUD4b0WEapYBK/CU2qhYNJ0KiIMY5oIyNVrKiQ2gjSA6yU9D
1GVM4cnHqN6Pt7MpbIfJ8PwxQHkmhYsNSKAHLzNSpZowEDPR1kXVYQTDsjgYUJdyDhmQ9Z0zVZTE
ww74oIKYMcy8AyzbVmGQLcHTyG8mLiL53w+W/40+ki/07oXhYe5VGxQ3o7hDyApflhxYl+a6+oIT
5lCi3mWFsYuxY7fr3v40cyDYO7ODnTw/zFnZC5NbchQHOxRMDvXTGkq5CdH6DWWU3uazP/Wy6zNB
TLyICxrpjV2XFDqCPNfrAAS/efGh3GVk+ztwTFunapRdomkbJZSd0spyOQNmB7+cQpw0XzCa4r91
ofJDwX5y0S3cJqEUeJSCZI93Q0nWzeEOrbuviyfjoIoLNzJd/7RRarF2d8QXh1Kq9gCZwl2Hu25k
WXKlOKSi1GYe09F+QgFSGLF1nSiOZ1BDN55cFNlXVFshaWcozenZUkvikKVpIPOiKqDGwMQwFcwA
gN/7ridgcXosFNBWQ2sDQJpLRHTCM81VJ2R4b+1vvic0cV0hYIqzSQDRAa1qee5TAX6ubQYIWGKB
BRYfcz5S8dWXAL9YvWqrASdF4dmFRv/AhrARs2UDdxwA7FNM/Lzw43jyp69Y0c6Snz+UQ7Pe91FQ
hFEoCi/1r0yVUoAtl+A9w/jLn7wrNav9UImSBBrZkR6G12iSsHRsBqHfYZR5W2tMzVjFsC78Hcq2
7asgD5Ems4hBSY7u5ygBXF/fzftyvCFwlEkcwFJ4oD4bns5kbEzL7JgDDife1YOt+zJXmaD1u8Vr
fsScGI9uHWtYo4OP+fGUyLKxjLxNyCR4a1A3CHMuVIS8OOISw2aTmUm8NWIHwU5eRVFfOjBwjLC/
FDkW8zpNAeAE/LjtsSMbYZh3aZOFMePZIP4CsjqS7/Gg8yL42hl6OB4FV9Z7fGiDiXz8mBHMUXaf
BFlA+V6D5tprjzLre50qGkeoRXN8/w0LsfFqg0oMPDwq/nUtLPHb5MoH5WYGhAqnm8CPb8EP2Fo9
TQih47aowt/SP5WtRvp+0gCTT90h0v9Flk6+2GY97ZeF+BQc74AKPLuYwYQwFqKcVMSzV4BdQmzV
vFleEfn3zCFZILPJvRS+wsNrChtQl1F+qR9c/yw9AzbZ7rDXVqVOy5S+m4BsQ24vbDOorq/pnQvM
zman/dqv2VwKDjYbbrCjx9IANqZlxz/kCP4HDIgSy1ww54gK3zZV4rWUtN9M+kjxtgqqxvhuj1bM
mrqXozENglbF7JUqBy90Z8n/jpKRkwpg9vOI2vE6xYa9tFO5BcCvV7Zjm5hepYR8VOeJNOe7GGGY
WpaQP6oRqsiv+6OIEt25Vj4Jm7h3XFuqOV8tCvry5NrCT1fRvpqe8BkF2G/d7gG99RIwI/4vc710
BfHbXQu2W9Muq0M8O1X9spiWrYVqpep/ufhGJFaIKZ343aTzu7nzE8bHZpWngX5IHzim61UJaW3o
W3eMAu+UtHfrJyXh1zBCp4RlZsuoJjTQBdI8yq+Z4pZNuM5TNbLN8BLyaPb2pbFAZFfTGaSuemzC
QD+GAG3hQl47MCTCzabeaaQkxOzmbd4dhjOQ1EIhpSe2ZRWjAFUXM10F2xccJur4Qfh78UKdKM/e
LntShXN0jGSWupzx6rj0gFzH/BHGJzAin724KEE2Qz7SxybyKlliTynaEtW/4k8TUQ5vYw/1VJss
4ZiM3wvDa9hv1HTXYnfwEv5HhGEYmmwkDP9JKNROBpYl3Q63lchWyPYlqyoun4GLOkd1yacbxDMk
tkwJ8ix5qK4hw1CHbBpC/kg25IvbOceywGcogNqMUK8BSYHIu4aVH7GTbFm/FmVQo6g/fS8jdLcj
6z0RK5eACNdW1Q6lw4Gvw6iF8tbtZ9c03adgQEj45XvI0w97W6YSL8zTYJJX7BtCpem+/T4hAL4+
DmmojbH9dYCmO5N5CQM4HRmPfO7NFNbYHzOQkH2xS9GM/7EtW5fw3DK7OkUuuQG8xJmRMiYI5EEE
jhJ8/Rl6cU66mWnWVDYe5VTkej6EzlCCZ7GnqSEMUJ/XPdrcdI3NwusHJP0fVvDxHrtgQ7TRZc9H
37qYARjIRuAViccVdnTZxkD7iskwhy2fiovu/nRKBWM5xy9k4isz5dUCi7FRYYKA4Ml8JCUahVrD
L+5nQjnxAAqONg4PJUvwcKdMfF0kBMGDVNc3/QnVSNYQPwk5Zqmwq1pk1FoLoY6nIuAG9pZEYcFh
WHOLGs/vMX7omZlc63xMojotBpz4hjm4sZ+4Tg4osmAIR5zZ07CK91qBoz+j8+e17dmqxBtGwnKq
M1AKDoAS5us4g1EtkizkgOfgn26yRE5MvCjoJcC7B3K5TvbFe4+5HmxTdSRjOAyuetXSeP8i3XsT
XUwPBsNPVt7FvgIEifv1KtTrAWl5lEH+UpN7trfzGZyGEo7KCYuJ6jrmR1hT1iFOCPRvXJEIPtki
/iV5DtThTRW11GRt/aveyiyG4YS/rlKg/Xttt/7npqEmlTa6TF6c8zr0XdpUCBvTNi5RA2m5ftba
eaLt++V2GyAl9czaPHWP7PI1xa6Lo2mLPOwrZ0NVAnxc9V8TUEWAdc2fvY9z+IYaH/oa2Vnz2Fm3
+xivKLgbhapfzbnba8ruVeMSL/DIPIx3QpFeesp9NIu8NeOj5w43z5FsePEZ/zcf+RHAaMkxeZoi
+Gca/0QW6BK1sFFBfaq0DVymT59vjzd/RzJTlZnHlzf+7pEy+zy1KIEquhrPxF198zx+suk2ehZz
a/49SnyaR2qU8yVWO3pJD9VX8mKiGXRk92lhPQriTAlRm+ckWh1LL/OqK7D0IOUsa6y6eF3M2A1D
YA94I/cc5FWR+75V1Yegh5i+65JP+5SSv8x6yZ3R4otvv8IgZv1NjPaPnEEUrhyFkR6buYk4XkF5
7BHOP1QMcapKmI2gGuxbdk2m7/zUFI56AP8e2zApvQ2tfU/IlTYtAdJTf0h+ZcUTKa65bPx7wfED
bV4YxsYU2DfXmmwsufFb2I3VBC0zyICEVb2/DaEU20WVS3twtB2ohRFl3C4Qm1brWAK68GfZ6Hvv
c2RNKFMPuJEc6n016vvMO+Tld/DgTlCPc0X/O2Xiv8UPVdgzUmp97R9FZdAAYkDOIoBP9VXRimm6
A/L5BZ5cAfAdZApFEs+gH06bO8RUcU5aGKNO/zmPmNoU7yeCriBebeC/aO1yTvYempjC4lH5VoxE
QjqvBkxNwCjul2P6OwAIlO5xt0AOJnpbKmXxoFqcNpa7JPhUor2EHLtKWdzZDhIdtsj7MsTmGUX6
AxvylrPrB8v6UOSSn3c3GoeImaII4QBkNckCJn15Bo+jvINXeKmbbqeWLlfcIuIhs4wKYDI+vG3G
YKmBVLBdQ2e2v7tY6vzlf+1lkxJaAdUmEkL0XSsbgr53UhrEoIbcYcnp4kDkxv56FjvejlJkvo2x
5hJ38+R2cgmI560cl4jnSh2ecT5U0PCbsf/L6KOfcMz4p0/kcPiRV2IJBf9xsDnL2qHH09mD3Uw2
WXfolTDCDelv8fB3edwaaFeWuvIceYfkfgFO4bcoxVNFNL+yJ70o0XeE7GV1xrmK6TXlDy995Uvc
0TUkjn0ogkeB8N7lssDh4xuKpXAYlOqzvuSrgOQPqYZpbIMx9LpWyZpSDWq5Mwa1FLsKD5OAd6aH
d9oluPNtRQPZFWkmR1PhBJ7XY/HO6T8oXqK+ZvGbexPM0ys3A4YcZI3dd7PhANQjGE7kzXSMoO6I
BF60DLxH2rQmVXGrxlr59L5csEelA8LRINpzRHVZvZEwY6YHejWf1o2cZLEW1fWCudHKcRbXPC1b
Du/i77RJb6lQSPUNirNu0r7+SUnClgBQVlAYq6X/Kwb4uDPCoTYd9R1MlJ34b/hHEP0UlmtZaieu
tNMHbYi7soU+MngtMchpezHes5KadGxAGv+4JDibMyZpMEokz8DsU4ClxrossALXA32PkVPpf3y7
Q5AAE9hFXuLGtCxCKIIM6RZji1CqITclZQLpqxrGcc4ANP1FqS7HkuA9Rb92e8ZaAO5yo6nOM1bD
EACKnXJ25zlufMXE8wG4LoBB2RoheTubHupfGVMSjgrQE6irdekIMu++4b0Wu/rEzQIHlt0wLsGy
9H0W2oMKe3DE59TBHuQK76XmsmpkJTVAZRcda7D99GblQfZp/6XX/ubSWHqhhGUoKFUhcFCS2mHv
GMBerwK8pGoiBBQ31XFvLSAmccaL1a0B8SB8kDuas2x5XlPQOAqy/7yTxdfxk6Gd4cIDabZhls3G
8isBh24LXUeoS0RRh6aY0J1YTyuIRZ3WknBfNnkH4wdswR0c04954AuEplDO8jf5DQdCbT5PLzJ/
jPQYLIyAgRUh2igRKar9UqUe7D3VfWNsvxj3Bgdj/LL6QZwwF+GkWD+TgSVQOe3rtClYHnaWOVz0
2+Rifrho97QKcNqSVLBn87B4AoD3EwnLwaFvQW7ZfjSm1XLvarg3IJ6g9VQOLRGPyaUwMMAI9i+D
EDTZfo3FjxB/ZX07DgrUwGihGr90EmXAYs+O0a06W2kGHYHEKghLKhSz0lTBXAcXoHpZQYGFH5sR
MGHwD1oC2+s0xT4Evo7UEbVSg+21VQNVnpObW2DPKmZgZgX3a88gTrcUeiG0M6ommk/WgAMHz4KF
TCEztu6NVDGsxlH7TEWlSkkhnOkkqI2aap4G17qsz+Pr0Lvp1VE5B+ospGi7snTWHn+yfbBq+B/G
vL6NtcHaxH5+BYwIX0Xj59rPiWgqeX1UH6y/vYQvtxJXuoo9vGdyOQiJp15Y/3T03J1kj2t1259G
d1rCG5DajgB2XXplUqNf9PltdVfpcy4Ae2VtSptq76gqzrAFJeyw6lTfTKfAJ3teylAO9hmq1ZVK
DFgczsA+fiAfo9P46ZWMoqI6ijMglcWoFycSsoazGkIgEUEkxhjKiS5+g2c3rgVFV32NeUf6lpAL
XEV1eP9JYPmKonjBo2FhLqouYCk+WAtQDdYyus+NLI0dp+XriHCnaxaA2ZCg9OPVKyjpKSancl5O
UMimuH6BxcfLhpoIexSQHGU6w068jF+kT7yWZ2xwqPwfOZRWhMjGvweeU0LntZ00CvOIJyIV5RcE
5hee48wAzz2OOEez3561ogRkJi6UzYosljZKkDazetXgQOEvWOS3p+cxREhFHIAcHPh7QzC4RsDV
Ws2B5iyMMz0xT+l1wClx7199aKZlM/IjaA4858Af97YC5yaQkHLzuZKr15e2bVybYdiOXqEKJ7Ya
0VIVB5kTCbkgK0IcmKlGJBaVRIjF3Q+P7JmAcfbLJSQxEZbrywx1DgoeqoVYNlyLuHYsm6Enky4A
qkXTGyIBkMSxcM1spDtMA/RuUwgMhlqrO644OK1OtnpMIsZI6wOQe51FGBQXUtD6lS3JfioM3wOp
PShfg5nEItLr4gVvpnvBL6+55XniCgNF+tbtq7Iw3mxS2FNPmWRs09TTmEBPGmhlmTpovx2wbGHY
YZdyulp8ocbJ5IT3izO6QLe8BM1NP3NRFdrl/GeocEzETo1JkLygZqSovT5L+mhT/ewNCcpjiMes
xj9juda/9gpmDypByGsawcATSZWbyg3PB4R4QAdOUIH+qIxzlG49QnVlBjA+521XcgtAYibM0lTE
EiGdezcg90gBmggs9nkCaQNANki95cNAyyfPJ78IHAUkHdPOv7wCSvY2tQ6G+KB/sdMbUij7l+Z9
jow/R/KhJn0OKwAhFVdJ/pk02lOH2BN/pAoZb0Oa8v9/aDeeWG+CukqzXwt4Qjr3dDKY9JNGmaf4
q22dw2ea0Ro6xNS4ZAk6wPTXLMddIWSbN70cSmAdOz5TCMEsCj65EG2mhHr5TvP8KNY9XRzBiWj4
kd4qo3/xX0++sMlt/ndhWNzvtSvTOhm0omWP4pCh68ZNEftTZ/ZHxn5r6pq/ZDBgKnCbYMO05QEK
zyvM5HqrFDBRoPM3Df3ksZSWe/LMZu8M7Mn5j0BpXALaQwC5+Ccpf+bVlMtmdloI0yCZNRGXlLVI
tBD9r7AlEL/uvXsDfAHfn9sdFM/9MpI5n4SwlhCVPXv03ijQ2j0rzcydWCBVqvikIoas4ruMIVzl
pROv4V8Snj5U1bA47bWj3XdBe0MQHygbLEcfhvIoJKcLaTOLY6858bbkydVyQegeoXrzZo2Iq1zJ
xIdLiYaxk8wKSO3yNTSAYN6VeZ/TplpOpgf9zGbSqARpggcz6Za1P8XdypiLr6H4nO613u9Y3toD
V5mBPFXdmh+oJKpjqMqm9YGTcXmtf9ghPeaTTfQmeQUSqNStAKol14JFy6r+bot3e04hUwy5ayES
09cgHbrD2MXiXFOnIsNHLnAXHxpoBxkqwa9d+CfRr/Ea1TOElBs5Vw95CgrW9cCfaBhTlxmIcJzk
kn1vbS0zqbYm9d6u0IS5vrjsLCPVEGRzujhJGbrEdlozd58eJp71BAZ7wgxE8zMnrpKG6jZvYqit
O6b8tyCuDdf0Kl3ZMhQJ0MHKS+GkemjaEtdl072MLFYkSq7mfRvXUtSUep+INiHnWF7hIFLnc80+
bCg5b1+08q5vrmZ6fqyHElQ9IxIRDdiwFcFelTKDFpqCCVFZe3PKaY1lFt8vdCBwKXv85HGlhHkh
lYZR2JuQ/xo583Il+YLCH4nNH9OAOmE6QQLVkIBuNBLkvICzE4LjcruG7BOTOwdi1ShSQmvF4crp
njmGXGn8G0FaXzLaPkI8ckV1Nf83/6s5bY/Rv2YPaKki2iVCvXo0ESV6s4fa9c7Ov9BGUXVobCon
yERa7eHGWZai4zjl7tnbt929jQ+zgwkg3EwjozVfKGX4ItaZ9TA7U3u5aKKs4W//JoxDRXZDlFtc
0aQAErFrCZ9avQvqMwwntR5j9OxfMJUX7GOM0QaKK6oTwEZOTxBpyz9yyAWouoNiV80WJr/qAPQ4
+1uC/06LGdkM9m4MppActQdJ+WR3YI+2H4rIi0w2KEnRi4qNu0YxkSVIHyNCUsl3pUpZII6VRZtr
Ozhqp+QEBwIGptnDS0ishKElj6nDIl/wqxKSDcxlyNKz+9HWNGanr0QY0vhS1prCmLJowCRIiVfx
ho3HaeR+HVTq6n/SooztCcLhC34fd1ac5hRPXIP4AHZA/PPAbfWlskB2VwwWrY7UQUWpD9gKcDUN
awCW19fxEmdsFIGK+u7/31l8aIuWd7SIve5ylmVuaa3ehMxswjK5wl9cMx7Dgft4/6cFjEMFdGx+
QjbvlmO7VAQPV8sAP27jNpS+HOwTrw9HVQdfnzWwjmCIhBlePsCqjmY21yCJnoSxnR9MO+giguDT
L1j2GNuXNLeFvqzOH/tBZ7fNDvd8rdkjQhZ7cjfAlUSfgGRxXx78bncPNmtEfw7uMU9ZNzi+cTH4
xZwTP2cJD3xUyfY/D0bLXukoUFKz/mMmcz//1luS41c0HRXG5Ny+3wGuldRloG9uciMrVrJScd6A
24MF6TI//BavfpPy5fFzr6/A3Ik+db3omeSPg/jX6pG4rrMmJzaKpr+dUJDXaSEPLyuSsG9eRRLZ
Ratt+nO5ifK3PnjgPSVtcyaNfIpZMBYCwZjE82Dw/FLURD9JLcr4OJBx3QfHmAV56VWhSPn9W6Q5
oPrFI1e5HvZMA2qdZfKE0txAXb2Ge5WT0rBfKHKW/8JdOwgg5kJSH6hkiaKUpCikb0OkFdXdAQiC
3+0FfQ6XN02RALJlJoy3v4u371U4xGVPwoDWEZxr2M09ESiwXrqnJcE3fNY0KnaQScduvcRpBlQF
6fIbwCJpOoswYQZYuScvE7H9gmghX8gvsIlTrV9JtPWLxftchUnZ66MNuxqTs4A44CFsppgqUyLl
QzmWYmDPlgqQFoFhgoU5UtK72ES/JENlEbAc/zh7RDMXEKbIK47q424pdNjJ+xHU0lpZEDUr/ovw
0tFwuQydZU41CO/cyPCv1EIPp5MbLoDfrTy/ScJH9j5V/XIfMl+U3cStCWD2vu95cfSkzAZdafsw
UwgKYaBP86r2XP1ZzXApFeBOELDwJZEz5jNSHIYNOR3CQJ2CPw4gj1xDkMdfVp/pEm9ulodePToc
erdx8iqE3i66bruxVckq9oKRN7MiPp1XQBCb8PnLPM5/mwWFKIH+lZ+/fTcoVI2Ir2o8SMIA8fRU
bANembkeXdVhvfy1WCAnsDj+1VVKCQ3Kw0fOc7N+sQrXSJIM3Qfigtwe3nHFDKASmFrYedLnkmPB
+zazZigw/yNpnbyF5BeenBm2YzJECiK7S6syvcsjMBoCJRLW2VvnBxDYC3ETX41TPiYwx4r799sZ
qZ1BnDB09DFaoFYU1vRxHZlW2/tp80XGjIKTwMfFY1KnmFIvpS8ZJ4LfwbOn0N+Bak4R9ZY06/fc
Lt+42O3Ssh5HghUjo8JEZcATwm5c2GiMHkg6g8+R8t7A8Cn0q0BJwqEtstSfmXFuL/7Lf+Ux8BnU
/7ENyudkVs7gYR08BwIF+6If0fiq/DjTFabwLmY8OlhY5BXswUI5ZH5kttuC+QPZC8AGb5vjMxGw
31bjCuiDgR1Az5ZZnmpl4+S/lrluyYLIiSzbOdgiHCVSllLJIPBmIChK9k4LLAeCrDlGuYz/d+Vk
f4YoI8fjwTIb+DiIru7Ig//TVXFtRGBzOsNRC+94co3K1x6mXmKmOk5gCTdf0w2RabcLMAoJOHhe
8l00nkL2JNvCyhSLpeTfPQSMSxGB86iDXPgUME7GyDIzN1xslnL6x3EwF+Wt3MKdf9/DHXiryR4Z
DBE7DzOyfog8aaLZ8BeJpNP/S1nCo6gEK9sQ/esZDxVSyfpd1ejK9qaCq+mTNtKl5ob1ROSpfhQ1
FaYm6jGi0PDtQhYdzC60GbdDbTOdUlD05lei+UG4hLRghkx6O9HBH4NNS2636Okuf8e+SfXM3U4j
TTqGdEgheFkSyYkm/pXEzHgjwFLk5y9HIqbR6zATCb53SHot8XvgHd/jg4tahZZm+yiYILiM/bY9
AcQK9NzSvDf+KFqX0QMUKLcGfTKl8NcJIFi3hTje/qhPORBgyZBH7RRKxGOO9fv5wRddRz1RNaTU
pS6pLp1mvl3swXj4oUPgDFUmm6z29mLychA3h3A2z1/BXDK5/Qa7jc7O89ShMmu/hpaUwl0qzBC/
zaTfbkBEnCVxETRw1U4El+Z1dMK9o0e+yAySk9Wjb8TMRuaO5u801SZbgyn4kJ5/f86V/jkSJTl9
2byOS1/Xd0z4d+ZajW7S0jmzB3zPeVp3cKk54o5hvd+kPO5MhzF+Q/EpVMSFfJw9UM0vaHX+8qfI
IFry1xWk6XueQqRzg4p1BNkF2/W+tw0Ggl0tAdZcKB7B4mgRorJQaM4o3f6jt9kzCcEkycD4GI3f
bH/UnjCh10tfc6U1+Ae1MZ2z2aTQC5F/FHVty43MJoLQZB6ZWSlDb89FEjhUTknyjhMPi9ba5zvw
Y+QoOrV1jWuM5fDA5pAeK2fvA2eapAp2TaiBYcDLvB38kxKPJtVGfuLBMm5nxdU3MTp5P1VPGYfk
eGMZGBbP8IbzDqbJo57FvRCC4x/CcxaoAibyoLyRqf7RFGvJMnmIqkYndktOXlij4FkF/2T8JN1F
uz/PfAsw3OkNMSFjcc1Bv6DyGfr2Er0QMMgSXgC8v5G+vJiLBRgBZl6LSoWNlcU9/raDBpUEoMqh
eQKzTNNxJ62UWAWdT8a9f6pOuTmAggbXB0T42hGesXvH+0P8tvDpgxxskidDWW3w2U2VMjilORFA
Obj8GvOzy9EuDEiDjEPf7weI81x6Yy6kZhz5ANVQCTxxsp5Nelrz+xppwfvounZm2eQ7MB7Vj5RX
Cj9secNZnNiVDOlONAowuJP0nY8lSjBZngCvzOLwLBDZEzn8kH7rO0S9nebMebHa9XmFxCaWtVxA
iL+7Yh6e+jlPkTdUoDDoAkgMknIc9ZXj7bAPs5rC1e4gtNLKkt7lmaRFq3UWZA9EN15OzRJ/ZQk1
Z70tDK+4j1EGWsqCJS/+yrtWQOlNg+8oOEcgBsXwpsX7C58FkRlhaH7emRKz9A/xbyr0OjpkqV27
BpGuEL7QVXpvsSOrCz4OlJtK2q3fLSuKG1BmNwWA4bQjaXZAxJGzdvwW3xar9m/cRJro3NDg70Tc
ExRXU8ph265q7RKdaD2Y2ivqTiw0Lk/acoYrvHSbP1m6QmJlFHx5ee2S9qIOMDn+TRdAUM2yE+os
TlnsStXwDweua+p2MpAIjvxublsP+EtN6gehhwvZP6o6oIRHDu3dtrwV14RMZBfN0Cfn4DQYhIao
u/3xbfI5WqrDC+mgf/TVqyJdmTKSNyRE+r/q/F9TfYTX19zz/Q7AazlG4QYxiElykf34dK7TZtnb
n39H9KIFzgR2BqxBY6XpZXuTdfUfcyCgSdCxPnop14flMJ6YlDN7bjC1Q1n+K1jQoL1Mdb2aqvM/
YEZZp8iKm3vsOHaZhj2L+IFeWitRaO5TYCvHIc383asD5uzbV1XUqHbOL43wVHzRKCSK4kvEYZkA
wa+Z+zj5XYAp/g00ydfmY1JCSfVOcJ09N/armchdFT+BNmWUsmkGbBxB+K7yPF9zWpF94okth8Wh
wXBahPChOuGhGYbu6O06OCtSW7q/UesJ2FaaCT3b4kF091FmCmgGtOXJqGZ/G1+/VBx8yskXmVug
44x084NBtmN/mw7IHof9lL//FmmRHDz6PkllPUvxmuNaxRbKMhJWjCErkATOnuhB7xf5GG715YOW
mBNGfBYtp1wlZkAgDaJhpnZsUews4EXah/oUqw8X+O3ZgRqRTxdJ+netLf9NW/owzmqXUSluBk1J
RFakB6GTpXSC42d/uyifc/zPAcY8PTvDIXNQ3IoXNvzdF1WjyaQIt29z2z1FJEnED7bX76LZukWg
tXZ6lQDs53UmQvnz3wB/bC4BjxldtTUadc+v5TNMf53H1nDvz6wuFKiS/3C/lrh2DTqvCDrv/nmd
UzuFZ+UVwXO1gOEfTMPGXHEqob4ctRMee0iMsAfq89pBu2FrlSWF6HmlaB0F8yDPXE2HyfZjyGTW
IL9KtqMFAoEaeUlTcmdR3dBFmrmbYE8oGuKSNBXumd7kog1jPRRT73GybrFRSroQLP6AA7fnx9rB
FeHbM7t7eNGvOCmmJaP/+/sLRSL+fJzZxJpuDn5mY6xtnUyMmKEjQcPMPO5e0sPDpIwPV/cdpBww
oWVE7UHVaNCQoY4xXdsaWov1y1Me1dujr5Vz7MvLwliJUrz/lZ7M6MkOVgoZX43LLOWXMVrXCzb6
k0jUHV4ap12/JhgGBpaupk1w3J6gQSq61Q299Bhbc296ezchadjnxpPcZMvPr8f3CG1lQ+L3U8iQ
4eL0ws5QgWzhd6QpQti8YapG8i47yqxdjDddg1Kt6DeV8D65xtJU7nfQKdt3OikwlFI9T6fmnO+V
Jag0yANzeaql70wwihN3Gwd3uIkP+ppx6S1w+UZ0zHwjdytspS65aYolbY3Wz6VepXRoOmnLptIN
ZCehWKzG/cRseKCfyB5nLJFzCOEkYqnx+q297JkOsLBKSpotsDzJKFsYTjl8yPucV0yuY8V5RiSH
1vy77sCYs4P18S6WOFeaa3FZGXRSQnN+qTJq4ulWDAKBsk8vcRXWlaoND6pD1jktzsmnEWGWdc+N
fErDKcgE3lz8nTdy/Min35G7ch0ZUSyWFkwEooDOS6XQKLw5+IVFkZ+gWLUMyzLXo18Q2jWjZFFW
L8+no0qO5wcGWM4wvTHlE/EsmTroJWXUlC67/PZe6KLgCPAIUl2qX8IcmqdvpQ4nB+6Sv/BSQ3Cc
dccR9wUIWysyciqHPLGSZ8KxfZlMYZGI+zb8IgYgaQzQ+639zmSwtqyO3wkw3RjNjT+hv0sWUeJY
IXZfqiqIlmcyD/zHGJZhHs07hPXmrgF8WDIFJiiivHgGdF2RuZkW1AKIkl1qVFY1CXZwjW5EHF1Z
uEFe/uZSVpBFTeKvxwZLQRPDBi2FdM2HtHKlAlnoVI3OvNd4DbG/70j8lki5rk35i0Q54h6YsRem
TH+sZ2uRvhr1rWHiC9DN9uczo383JLXKzCcDD2ONLNwQvhw1y+bRgQrOFvUJlZUl1YBF38ItWnn1
Ah4k9YODoKyaLj7sSklJr4zQII51nUGlk9HleNRbfoGb2hXHXfym7S6GwtgZIJ6ci6GZaeobSP4G
3tFV6DuTnXxXCVsCBXyuENJbAPLodtR/fcEx8ehXPs+nF5vevh3j7jHurEVfN5QzEdhsv4494/nE
T4lme6vsvipJW/8BH9ijMj2vTxPOotdS6UlbF5LGmvNAb83nBVKkBELI5dZ0eMR5JRClMxhSiLr6
TAU9wjV0LKH4WzLy4bmdd3Mz9eyyHxvd4s7Lz9U11uzctmZzAsjmQI87DdeNmFxBC/hX+DcUclr6
aANJXCGdAnX2f4T9AWeBqsaVEy1VcJ0TuMN6qfMD7eWoxP20iBcXqeqIy0s3yENO3iyaSiuLv2Ma
G9WF/Px5JQx9Ky6LES4nJQ2IetOil6vBjNYiuMG8m16kc+XvAL1dPSheIt6mmBaoDiT3lTTMaqQD
v3Jp9LWuK48YHmMzmmXsEVcz2HUAFVnK/M8oPDlzwtDRBcKiz6yu3ztBw4eBrVVEMyJC8280eoXx
HDNbKAU9Fi4tneVGUT11gUpk5ibDMQhbDUkJkV0bobYavPGPTQTScsaR0XdcMyCZVHlXKjFo5AfI
l/8JDWNGntaI1CeONw3wY2PZHhcx2pZqIcycsDflJRWg42g34L+BO83NdmC+qp6NwESanxhNMac1
qwYjG2d6xqSJ7gmZ9HMsdNpNZJBLN7fF8HbRfVO+VN9XaeOyhUnNc9sxtBSTxKb6n6Fu93Fqlo6b
b7/Ajj+Sfy8UOkHw0hPTxFW1ObX3qIm600N8qysL1gP8f1omq7Yj+EpuMNLTmgevY6l/6oCiSy5X
sjMXIMPTjahACAyYWRzXBGjxnfdr7PGYO9HsRVo3f4lWFQx21MRePmAPhQnPa+h9FW8JPwf1FYpK
M1RLqTMCJcfv9cVRT3KkFLnkGyLVsoPCUDrQ8EDXmryw38/l1hkeIyrdXHigg/+TFrK2dgCC475Z
SstoMsdIQ9tBC6jxvI1Fml8TYWuyJtPOIPwALXxIsZ1KhDoTWGJsgDZkQsx/aq6YQ/tcB0eeBHlG
zsgunK5snXIfKPCitQSVmsLffGwc7TSZVZE+Kz8/tT+6G3ZNoyG68epajr0xZCzFK0XsKby+lJKJ
91HxnP6+SJYMgxWaHet9NuwNO2qh2mFQQ/7nUxdTqCMUxJdrxW1Nv7DDWszok+z8utJXQNDtRyJe
neSC+ZqkqM76z3VXkjtAtxBuhUYqY/cTIZUcX8Psf7DQBS930xP06Gzoo7xcs38NzM6eG4Rk+7Zg
9EmPEk8tTOZc4+i5EhCmEc+fOReivgugCFxrh6SlvL5FRtSgSPMdYyAqk0AOpS4iQJ/iIpEtu78a
qXwc9nQpuU3qNEbWFgvF1weidF467PV+Ry/92zmT0jJthc77DGSQIVks2FmhN8T7cKA8UykYpiD6
w8W5enWh1njrMUfrpQdSS4zAYa+lCe8CA6kxLTmLU+l8DZ8bfJsH7wfk/KN/tJrz+nuuyFDnFd22
HvpkvfBVQodxXyRDhBtw3xV/drjDyCEjbDU4ENxzLQbw3fQDSVa1/yE42K/mqJxV88soACGtMTkK
27zLeLKnsp+V2okkQmwMnfxMVPGzROYJoNVgW3Dq62k/432jRgxIA+m4OO2BpMSWFuK1bquD00vu
LZZiF6us+eFHhI8AKbg3jUNyTT23Jj6rslosOUSC9CK4R2nEHUvH5uiP3wN6LyihAB3OJFjywY68
SMIVs3DnxYEymsKnuPugl0BRqrEVQlniHrBLycHay0PW0fB5bnlLrosV65po+f1qApFQg15LLiVI
o3rUWN4a/DGvN579x0R3DPepIsWmSCBrmxJJKvVHOXOmqG/I1AHW5JHhMh+pliZJbQ96NdqD4qOl
RQ2uIrNQ82go9RWd12yz/QdQoBRh2aaT9GuyvlVLwBg7Q1dCsR4qjlLGKRnZ/rmPu20HfJz9Qz0g
tkDbWinX3PwvndiIysqifrptFx1PB97bFf506CD73xwRUGTj6zLFcThWamrWcTDZPZ9uHX/tZ6c8
NU5fYw2bQDOiwO2nlH6KVxHSrvobo0pDriQOhLKARQcBztY7OcFJXSnxG3a3vRoB4kRUIMbUUBuc
UL9X4TZffY3xxNTX+qGJiFawaQn28mvDsFBeAJcRzqnWmWhuCJlBDakD4zZRQaNlXlpzKWRp0i4/
0n2qLXESAyA/iYMhPTb/VYxdA5HT8bmk5TvkOrhGITzKsiJNsXRMYLfzOkSssfuebJkTC+yFpjdh
OWl57lsxdPK/3/HEmbDmvbKdpf6EFzxxQkdhWacGwrt9BIUzoOFBXN8bk8oC6jA3M8ZQV97mxCLi
AA545DSDywt+hFzNPCPSRCOA5hLMQ0tG4BJDSgOjc+sQbIhVU1VEMF20q8cDTOkONiBy0Zm9sJzK
dJ+aLYPgxADbBCbFsb81TPuWAVW1bUQNYaQzMsKFOmBsi0tXHApZGynjfawtm1ZvgQfYMC1A6Jn5
RuuvcVO8fjPhiV1jkdhjGk1T9AgV/u9hLvSKKEHzkgHmn3SBre0dz47qGHpax+P/r+geK7kkdIh8
gzA+5MS+K1esriuwr9+grkODJ8Pz8xyrMrk7xUFXOlHnZZR+yChGlVQzaXbL+XIFkYqQKQKtrZqA
j9kedOxyRaXxbCXccdlMmjVrd9c8GjOrW5uw8xPPEubQfDt/UitDqQixh9ZKV5xlOGAHmpBFcjNs
UnE1aoRFo9uWwWIKC8MB8eXb/I2FwK4FnpgzWQQ8GV56Jq9xjKMg7/Vf/4yX3Gt7BqZGizON6N/Z
NcIYK4eYRRUoDFutjGoP8cO5R9WmSxXhhJWuoBSpwgxbuz5fTCNW6PI3sgl7PO5AeoDjTVoaOEt4
3DDo9hNihz19Giv/SZPp8vXV6FYeBk0rqRyT7eE6Uo5Hc4pKkjJMdHqZ2FZ0OGBlPQ8vrOcuJz4I
m27NZD7h2Gghg2RpVlvcraEr1TfNvOlAUVA2fmGC+krojaja5FbyAVKgSjGht3NdKXhC/DG88M6y
248fR1H7qwdtem/OdrXnMAt5y3nmB7YqH+hBbEDeLDZsLKCdLPAWaye35nOFD22By7N4Ske5gI46
MS7fnL1dEgx1J6+Oy5Dx+zzlbtSiqUO0oZMfpEjuaRNKG1X658zVBAL4TljgI6vpUyIk33z7QgXs
Ctv+IZpWQckjI06EjqtGJI1OUm+rRMc6ekmEXunjjZMow+F2dm70l83B5S9sbNKb2ApVbOsQE7KK
8o+3uTjRGe0RYOHE3XaeNROfl9pxkqfa6+ef1+yaCqdi7w/2S+i3Co3yVl61n3Ka+cvmdWqQMudI
2KNi7t6iTU3d4Uo7n2brEwxNUMTmndtb6Wg5gJGt6UwG0sBucBPGKzklG+irOmYfNwS7wsDzcx+w
79NpgCUhbrIj1RCNNMvst63QEUi6ehsenUmhLwS7Ou4/dGxmypzSHL8uFixTdp/gLq6H+9F2joYk
3YjCkBV/jQi6EWawuanGeJh/PfdI8f2ej1aVBI+WAobJIzH5sFdGqGzbyU7MK0zFBJ3ytJrPcfvl
w6jYr07fc8sN7rdq8XSfjxpNWjC7ExHOY0D/d3xhUgtBNtoL8HpeTlI23h9IPSlA+djH0/m74guT
9k7sP+Umys2tPa6ukK27A8axruzvqG5aR88cYIR/1N6wqQj/6KODqapl6jyK4VTVbC+SMFcPU5Rv
fqGeXVs5oLOgZhucq4ESph5Q9JpaLJZe7Mfn6RlsJGULjaxw555XjUlscxm5bMEvhut0qOFgJH+I
k5b4R1nT8FA+u3ZKNBIM+M2l5hlgxUiyIteBMbLPu568zSzuop77gLJC0NRVJCRvwenm7cAkrgU8
sVfrafdRGFXwV1hr0twnCvB/kkvmrbhBpUA8ChTdNESH3FxRMIdS3IsiWu2tzxD3Pq+P3mkaarsG
WC8w8Z27pOjQeItdd1xDe2Z2Xqs8VPFPQvdXa490mOy3eaqGS/IwYh0SPw6FGt7PXdmjmc+CoKIH
5Y773KPR2BwicsqorqBcYSUEl6fbXUS02K16Oj/G25dNQb0Y4fAku5S24qanhsPT1aRhSmRMiDoq
E6ahV2UIOmXeqHOspo5w7qioMRKCNPsIGjJCp11QOgE/K0Sbe5jldQzPl8ApCFsMyLjB/JHjKUcl
wOSNG3kq/8mCcsTL9VlMnz9273hEm7QdwQ2zSV06l444tSu+24T49o17ZwPIaRzrsR5VZGbNeQm2
jOzbEUDMevmNhAdyXQw/ZY5rZfDKSV6Cy/7UG2kGfEoVxyItCon148l6U9c8ENbHt5YDGiCETKNK
tPXgU5Sy6dpyGSFtgKYpt3wkq/Nc/obJ2s8wLBkOIk09vfSR2KcsrWrHfQYTqYPdSS/TyrZIb6+0
EBSM1ID1hHep34M6ejgOQmm7zjvXV7yNp/xzK4CMDbs3bMixLxinIX6WZORyXW6f0+h2NKrP2qWP
hByQSR2qtJbzIlm1HssQ8LzcQVkbtz0B6FWr8rjQyGZt0L7BYJniQ8HDIGNHQu1H3i1tyBiacvhM
dWfnyFj4Qcd5O45uGJ+f9PxJLpSQqJtWodfESZvELL8Bc+z49+379nptpHbI33KzrXZi3CMRETKm
g2fhMoUqzJFLvTy/MFBwepQpHX9vAuWuNhq1BElFNpuiTr3FefojDvhR2tehTLVKf6l9e0ZNgPz0
3VzFPo8q956ATk2mTHHeyCNIZ/iXV+l9bIVNIZ1XOt0tpg8+C6zbBcwZxyT3iRlXSvahcP8JAuv5
gCWGVJ3crPkdXx7kQdBDBwfvDL76FhRvW1EEmtgccEKpbrw6+ZepAH15rLtOIS7GIc8FP0+jQVAL
6plS8p5pL8hJYyCWT/3A5REnVlyoWeeVkanG7NkCojHFL9JLJD44bCtYpq/J3zdycFGVvH0aXZlt
9Tkf0ki5hEnw0Sf6F1IC7STRyN5amWhuBEncLf/MZIMM5pgqCHS7k3qhmFBAJh5nENsthqcQG52Y
QjBsBpK26b37fkNNvbKODdleRmD2+wRy9OtFgouS2nCm0fiFpawcAKVfzsFAqeaim3mKbNLNNh3f
qiYCpSvFZVMTsKuloWHi3CUr+wCpJkGvYYn7f1Uif+b8duFQkrHyL6ow0TKelsBNzWMD0HC4vPIo
BFtqmgFBtEO3vLJWTnrQCMkbT1qOkcBofeCyn7dJlsxhRNXFsHZdb33HejSD0rbxB+rZ3DCLZzer
E8jXrdFVeOa9ltyRLMF5FhfoMf5ntHt7302/WCWWJo6jI4ZEj3HOY41kvlk9M1fR91t5WhTmCt6+
JsaorQknchSChvuwBCt4avr6yteJThTCLDteTwBfUUgDAU3zRNHAherQlP5JrZo9gNZ+sPO4ztYx
dsjvkIhtZhOmDPjeZ7u+Di4OfO6HveJ0nRACsxqv9CeylHYJVaCTGY2ltudnJDTABCitWNJXWfoo
2WhtFDGLaCT5eKt1jSTwuWsXzQETb5ldzWwoEOhau+YGr56h4a+v//jnflAgUDlWbSuQOG0ELFtO
RVAM4/i649khQinEcE1pXVRIZiyF1n27MJwK7Ob+Cp4HS/S6LhkwT1XjlIMrb3XsJIXFSIOjTrxB
Z5YqXiFNMt4/vRWllzPruq30fo0NJA+uj1Y9hZu/mnAjyQQZki9k1YpQEJ2mbKg7U4YMwfNBA5M+
5LOrW6xINiSTZQs3Tuig49RqBpp84f/xs1APggYNBWhiLZeyTXOtsBcPxtkrysYKoI/AmtZrpVc5
v58hLuskknUHrp/+N3e+wkEtmccru0pGOGvH9TlGtLZqVZDsKpfHvSKXptWSwdnhW0lFxfXbyMQL
oWrh/RubdVPJxXLNU5wDXe0mnaFa/NSKnAiS3A4CG5oue8871pOTOdAS5QeM7iQMAd6tvx39GD8P
7s1sH5dYHXnUoFBTOA1ECJK9faGIoIydCyVDvVqzsv0WLgu6WOwK6rYVFCQg2ozCpBhQC3p6fcM1
ExvQ1ye5bKxz5PNjcdL4z+FgJz5jovEzYMTnp+YkAuRvJaFSSIZLYZJnLtfYlw6PbfFFsZsl0TrU
9mx2JfGgGKgoobCwQfEL7BDjL0Ftk04kf7cv8s66CTVVcvFcsDyzJlkTjsFH7fuKuEl/fwB+sWiA
an8ceVMq8VLoCXQ3rgTSmd4bPawrGjSOT0nbN9vweaeq3mtMtttCcl77Tb0+rncHjlSMEDkH7sYL
BMOL1bEyYd2IdyWjdklVhXIGvJ6mfXSsOZk9RC7hIzc6UJTTRqQ57iDxbXD/3BOhoJYw8t6s72gT
SCX2eUYC6o5Ct6omcVc5Ts/8hXCE77wGorQOX08jG0cJagoaYpXbIl7DDyHB7TSQuVCpAGn2r20F
G+8ZLpz6jxHTnmijpse9bUR/tLdo5ARRZO+hB4JNv3aBptFSkJhBf65QdknXo+JAVzMpm7hrDLti
+KlQ2/SFb1XRd6MA//VJOVr5U2VnXukoxzN0Kv0UNCpeK3LIRp5ghZVMAYA1MAjTgqJNZJ4bkqa3
FFZn/XTT0zK/Dj/QbOlMP/jSzvs5fINKjEQfSlUSt4C02f1mxWO+Q0eRjUGQea7OzPP5Q2ZJnAE1
pPq0sQ+CY+WXE6TH5eSfAPLyhe7X+7BWPX1wm5KtDYFtXIGzKHux8y2kvJXwuWuQ9aysedD0YrBW
oDKRUJTb7S0/PdYicJcMRyWEl7hTvifIsSiNkNizL3siExdfdTnNO3BEhPCbsttlt4MnzWsrB521
ux504hvfYzmAHJ9GkJqSU5SbvIwPe4wZz/gV8Brt7z5PDm1ASyyYSmZU3udcHiLWAY8GOxVgWaxs
2YdcNXWMDze0TK4sZm4J49P4KVP8QWp9zfTFOmFfwS7v3TQxdoMjdieS5U5jANCW1gTYXBtJSM1Y
hSPLWhu5/gf7Lt46rGtqainxFeYlbA7Kl6yv156by8hoPT9iqTg1sIQW6E5qLLmXvO9CS+fje/Sy
rtbf+Umklr0UKseCFPwpRow9DZ5uFeGc84cPq4LZFvejhZP8K+F120VSdEnBQPox+cmM9wIj8TGx
du6O+l3ZWZSl3Bi40gQI38bkT5s5jW1ThFwQNFt/ppygOAHlHEvp7RSnxPdT+QR6/hBVu3vy/UTZ
uHneFguidUUu46zaMt7aCBKSevP51cBed6mkMbK1PZmzW5S5T27tdjZksWiYxQ0f4w4av6Nl+IWm
DQvcUm0WQNuiNyLLuuqwOAY6E3kQeKmvDfSFlQSvVD2Xqkoo4L88QowLIy9OaV8JkrvT8gZs2KVo
p+vF0v95ni5h/Rxfqr1M8XcFvaA+I+kXlRbeRh9dksfcrmUQPwtk5YgJzoovTxvm22ITxjlsK6j7
kHixjN6IAr76+QyCNZIkOYdST62R9TTiIIuikEq8df/ledsE0a2iON3aGLrnpHAVB+EX50x6Rsjg
H08/i037xBLnpmHhVBtWOsQPX6hLIjk5btYx31lgkngTZTGcQMtxqaNYWWhXt3rRb/lV4jM0jius
uyFCJ5QYNmh8BcEVCwjjQNHfhrs/wnhJc2x3WJdaMiKOzm6IN3ybEyGBRYkfR7TqfJjnND+bWgaN
Ggyi3ZAxOZo1jycINF4rXu5I8oBCaV2sOfCH6O+4ucHhrtCO4hLV5ASaC9tx/T4TjJOk3vyVGnAS
oFCCTRJbeQBjv5MPSfrjnHoHp1lacOQ7PZhRVVG03FsCCXp0KCvoEXZV8J11+517mxHZ8kyOkXRS
ztBybeEvia/8d1XcB21SefEKHSEZRJGYcttr76VKmAbPTvQcIwBUpBNpaDfwuyJZZC+DBsjVk3r1
yepAmDWCALS9EgshpVeUhXRrCmPagmB+qQoupFSKUOBKfUp/2OXswRWBS6Bsl03tmTAEbgZUzzbk
ozu0n+2xUSLQUmIKsVy/SExFFhxYQFS/Uqw503dsDFfe3MWLfBV4xYNfnb/MS+P8ZiUVKLnS0HKf
BerfDQGSUcSnyACNKp9Gc2TdbNOY5oMjm9OSf4g1U1fpr9Snucua6RAzLaE93q4qgpkSCVYIsGh6
9GaKoIe+uhf9vvRUZg/n7Ycf5AndxUneLGkgr4Kqxw1r1n/3OP2Rctsy5d9nHLmXgCi28zJNOLdB
lthriDioqhstgPEJJYodedyei3xNJ9pzzhJWdVUE5ZZik8dTamrDP6cIouC0aluSkXHBmiCzbGtS
3H4fSupN2ZkxQZxopjlBr6imG6hfcsuIUgEQh+VC3PLdEQ23IqsSYL0WtUCsbEx1oByckp8/3f5K
BbQzpMXD5BLVN3rltCHuNq01D8JBa9vPlkrFgs6Q+SSkUr1RMXBjnS8Q4deqJdmz0HyaI1DnqVig
yVOwkTl0v3nX/VUcO8Oqke5AKUUbYFXLXNCxrQAwDk9+HvcdWCpvyswU/Jko442Km2PiVxp6IrbN
RqWbX1A4/tJNpgXH1PGhkfrOaLEANU01WMUXHqc7rMHn8rE7LdtxeBC5HPMNlrJcnT9jUIINy3hz
pTA+U5AEWfC0n0XI4cTqahEPuBKWJAV3P2P1/zmOq124tSrvSbVcj9/YUg7v51ezJOPXc+NKf8du
/nkF0QDHZZC7cDn5TfK1pHXrvAQBXW2XPUAnhtd0CepZfbXePVkKjXHMPznZfRIcfdlQesWWkl1S
m1ybLXanOV/QJdBiwrKYDXrp8pF4omH5O0LWrcf0drkD/ZdLqMBfoss01cQJEixhZAvlcF14oHzv
VfdSdR2JB3AbLNDrlwC2ZK467GGPZVlAJyVr1IVY3fOxQqTNEFMxu8Q994PwF8hDuLOq2LUfdL3n
/auGbZdeBUVGtA0kQmzU9RmnnEcSNWUmPtgsvSiJwQeSadjdzbmD4jN03cZOGhEAPu6ZfEpAaptu
Yn1QGD+BwLgsIPXZw/ybEYjRPdD3YG3yIc1KT2QtXyyMT1HuOJhxFYPFNHJnssSrOZkfF8AvPKCY
XX0QiybK5ssiPRQYfoE7g1OEQTm2xhDRhTrW+kKKO3TQgBplF56peKyaAgVCvWaT7+c8e+0ZNPmV
803zF8n+eMo8CQmkDa2PIrYf+ites5wH39B5oMJ39f/X0NrnTc8uracTK0DiasnK4l7TcPImaHBi
SG396xkurYV5nISUfK+WiLBgLy1ZfB6ullhC6ZfOnTjc+JsbQ6AvflXCqJDYZw6k9mG73+UkdPsj
3ju7S1fzufW2B429hfWMOM4s5RizhMUpdo6RcVZ2hLX7pHaGfllU2hKZ1W/W6vSaIM19Ea/5CPkW
BBqtH82R+REileNq1/ElrWIjHZTlsO9vyiJe3Vob6alEK9pXIIWrR/DSaIreIANI0N7z7iacrr5V
s+gsYHnykPY32Q3pUhR0hKrQVua8cyiM0T3Q0DkfOORDkahstoxbGB7DdBTLWpqOqkj89/ekeNVl
Cd2GYC7kePbrl4HOeQeowmQVqjkt8gTH30o0kG5Kiv8n5NF/rZanDBR8QcIeIPxrrgGnBuaqBz+F
3TBdhZ10jHvRWwPPSlbZ5ksnvm06JSV0xovgUgzD7MnpMLPFa6KDz9O1olgN0RKS+eLAhvLoS+Ns
6TVT8UNrmeYyIuTwXBmfbFoAhYqBu3/tE7Nu/8j1ADVejmObDu4VLENuMGqCUqMgh4Ygz6pjWsSn
+a44/KlkaU2b+rAjJvntcxkTgeQWGtp9Jn38w/UrGTC2ihy/COEpMA5eWtZiKQWZF/p0VEglRoxg
EZ3GRbj/P9/NtlqYSl2T69+QoI7ngGFiyzcjNEBwAVosp2sVnvKhsh8bGDTbyAMi94uM3eR9siKa
MmK3u+rpYcqo32uTESPpByYnuNjEs0bD6HRx2f+9fTvP3NkgZEHm/fhz6Vo+3U6FfUXHr0D1T5Pf
50eSIEZD7fULPGkizReeN/DHwhE3kVAbja3kWPg2ocL6/Y3GLbhr7drgaDgCt2EJnCbKuUi+ZP9k
8HVeAaiFtlKI8xeBc5UggA99Qe8hvqaGew0h7EB8/8GlzA/PXicm2x36Q2jw2jweh4JCOawoSgWE
DD9rOpJxWPOEPGzeu3NFGxG4OTt3KG9dHcnfzOeoBmIJRcoscWWIhkrK1RY/SIQCFfcaHtxIYUFJ
dYmraV8LeUbnu7HgjiE0KcTNXE1NVw7sS44uz1oZwHcXeqfbDFe1uA9Oy3CrnqUZdo/jpFzcdEuZ
SeudIaA8mYp9bT5RJSzx0Vae5K2WbH/lDbegnQ6+8X1GyB5V/bAmM3/28NdyEeTKFTiLUcy3QMl2
YjD48rlt78IZ7043gI/L13qbUzw0bfv/fOUpU1Y9dEDuDBOoLLg7GDTthuVAqMucX9irEIHXdR5k
ggHE7R2+y2f5D2m4c5Bk6adYxpOgWra68D4e4U6oBh7B+tiqWg2FVNi1bgropcoQtwIWa0u2+/XZ
mMmohleDaU0FIdHgSII9mXIpUlI51f3EmUeFZBagZX5ahmRRusjsjQ5b6T9kDDrI+8714h8P6CNn
kZ8MV5aSI0iO4PJitwD2IusflCuLgA5ry+9+Lj1kQVugTka0hg0ECzB2HfaXEaKPaJXlaM3RNW4C
BfwGwDjUklZoO2b1jqbfGJaIZo6Tqxs8XE1YWc/kljjmDQx/VM0vJR6bGOVp0Trjbw6PfebCD0h+
C69PRmAFAL11vW7FblWboUZbO+mKic4Q8Q06Jku0Kw3g8PNqp8tA8/HiNOd+c6r1VOn1m4oH2xz4
trf0VZiC7F1AYORUC/CLemyEvT8Yby3q6n6c/a/JD19jGNNA35YJF7G552sIkO8Nb5aHZuaC1y/Z
hDIcUtu1uiMUPgshXyFGtjsxicelhg/4oA5pXdN0eEeBjZTEG+bqFDCbCVNZw7IjGj20MDK6+sh7
cF0Jmb9P5EPnDpBj91X46/UH4LgxOlmkRXxd1B3qm6zBdVxNaI3AAiQ/ixwT/xCYYdRBb4e9N305
Orhvvxd91nl9cd48vD0ZVV8JBN2ZBNj5KEOZggsVHQl+gtmmWx6UBy+hxJVHVJnvXfXO7UJGe9jQ
A+rg2brsLAtf6dmegQzXG/iRDlf8aHJh8j6jHjuELZr4PZCmJ16BrPIZnSQVgeW8xDPacwWeL2Kz
QROB4wyoyYZhW1yH/RcJxk4kelJnFD5AsFRwHkLIZrx9um7Q97sfjYTvuxF9Vw3FU3uDZqqrmjbQ
t3Zev7IjJe30wNA665ORlS8ETpvOAb0JIR+U3opZ/0mLj1n6zzwasyIeb8F8MZW9NZcsPsem45nj
1LSgrlpgMpOZ63t/xVfBvjJcnwGqW4NWQhoTtnkfHNjKuZiO7kndPZKR3aUHpAkMD7evWcX5+K/4
FwkFyAwiLDYNF5pTdNMV8+bSzQ7HmgmbPdMdrQ2IAhETRFF/n6QGK3WPXr02URNCOaFhl/ZyrqpG
HXnrevCK8eqH9sWETKbq2xoNkjhiatIu48ex30S+EsCb5yEFMaS+URIxLvEXaRTzGanDvirpGd79
5BXc9zXmg4tLRq0vwiMqfNYOAnOAua872irCo+wGpLulDk4gVt1H0QjPS+XG/aFXoZXh4ENjRfD4
DbYY+dYjP9L7lo8O2uinoRU4VZLZ7ACp3XOpVegWKR1g5CgrPutLz7+HtPfAi2JA7S+q0OT1mBYI
Otihe7F+OkqQHFoqAIVBAHFoeXrhGwejsV2IA53Rrjpo5HJsXL/tUfic9/tI6LhfCD0fLZ2GYe5q
iUDZ9rQTN4pxcLlitfMdjUsHt/6FnjSWEvBShf0qlIdkpi+NLPae5LwMrO48ojGQjRHx7/YNgJIs
/vQXv5O0AEQvVBK3wS7iNEuYrNIvxx/7mW4FM2AcQURKwEYuSDm/mWnN9qHij9+/1ggYpCmnQBRi
jhPI/4pHng+8kAUz8b8P+kWFGxU7Tgo7W1jzOw/SfdkiJ7UVTxLMA9HGbRkZ5FBxxiQucdxclC7A
W6FSMhaGj6qfz03FWgHaiGXFvWO+1OwxTsXLet80f0gBQE0oeY3bN4GEUtpspmUJEF1lvH0nClvu
efR5pZBaTJMpi6pUcMN7V1cGnh7gl2jEuK7D9QF5vX4U37vl6+TKKXPxbUujt4jrbdoclJDNic9O
meW7Jk833605HJc1RG0CaJrgWF0+wgkxwsbIRnC2AqlgPSDiCANuX+74N7PJMYVDQxw9hwlqtVSe
ZJcOpZkNtNDQ5GopNiNHENtIq4kcTUv0IpMW74SetTY5LDRkUlgXCr8iP+BTH7+rppcQ1aNd8yc3
SxzVK74hZ/qqJ4L4yLP1SpVFtpUQG/rM0tOXjqAcWwM4J8b0ZQMP59Fixp4cNNqgUf0PSfhnG7Fr
NOkhcjqDVrGF2iuwl4uT2nJ+ZoPYVyDMNrFTdVveGb4JGbVRKUXdkVZ+ivD5kogWLphIxrQDll8y
5O7dDQ0fpA2V6pGzGUxQJj4V88xB3ulwanywQDjGk7qjEFLtm0vbJ9fw4yHfj2ooJfVqthjpR+dp
9DU63LIoK4axuhuLcSVkYXj6ODgJloOPvg0Z12VxQOCCPZewx5AadRLVbpf14vk0SHb7VFx3Z1Jb
Pc+MeGtX1PX3stB8NE4eCNsEWCEqeAfCBkcyqX/CUlrOLW0QUsq26P+K7BpEBprByftqBxb9a+hF
qRQbslbcmyVaUPaGfTbYVi3C7wJTvhhTiHxwoOqL0qb4pz6k7RSKNzjM1bw6h24Ag1EtRSXddGrp
Wt8zy0GsXOx4mNd0Uc/oEJtDfEhFlI5wYLpUMpjGIwSmd8gff4QPFKTojznadhunfMd2FKkjpXKe
2NDX0Pdh8p6OzNV3RBE5X+hhOEFIBvH5BVlgJ239q7cxG9VTPAeNR2jSaK7MHOwiPe796vDUmVKb
xBBDmrJbozttsESLwsw8gcxZ4W9nIDl4BHKLXDOBVNdCJm9284hEinn/GtJ3mBUl+rrE90vrJ8Mz
6lDIsNC4pNTTjzDOw+HDBDFibHL4MVwWsA+rZ8I/v+lVX2HshXlKB6weO58jdDMo7WqF0kXKsU7/
GmKeQawrbWz1XUeoxdlCR8nU+1LoAforjr5MVA5IpMHleXF0/nJnrHZbd5NwJc5rStsFd2m78a6o
oxoVQDYwBPqUfQZNzH6117yriF4qiH0xzP9+/qKT+WpYWqSJmf3dYokLi06btr3jlBV/R4dJ1+GM
iiAQgLJ0H9BoNvFGEfvzFg/c4iLcsT+PUwqUXFUvK3b8rAMhp4uvN/aDaHUFOYSKFQjeHbM1t2V7
2Fu4kF6z85oaCTKGLQ56AzSG8gOlO6xKmywnTkHE5SMB21mE1rLuBb4d9bVfHQkeqeWPpp9GObJJ
4TlOd7GACubYg6q7wAHPVonidPx7eeZkQxHbKQ/mFPANEWzsSqYEk6Is/tydw9NNdBkm0dCMxIV4
l5s+fkNACNF2Ynw3ZGo+XERSCPbUyyzSiuwItdyr64/lOR2d5l3UjLdt17mvajDjiOfeiL6fAjPV
GoiuiNVWz1YU08DPvvf3DauyScf0+MfvXQxCMSHxqKBuyGZ/EZLt7c/KqmN1bPSnNXwP4bVUb2BP
VPEiHh3xMIWrBtqIt5LQOp55RtJZnhRu6ansFyzhF+wOyIk9XVBg1WpsPQbsfR9aYxrEWwow/fS+
U+CGv09LT0YN2ufpZcm/5Twu7925Z0nkkHgfrzfujGnNSP10i7N15zbNwFM7x+NwDmLv2oZ6hpSG
qFc2mH7W+dDteW3NI7hggnrQ1Q3U4FJYVQTlXpmxVFM90ds4jMEMYNU2oUlWQvP2VGC38O/kawo3
SmyOUqoZOw80q/sego9Bdi+emxvkDT0uPgrEip42DnOwyUTz0oD8cymsm/Uc2n8B/M+ac0NChaZX
pEN7Z7RzhfbV1bqhE6NTS8zr06p+XwN0pP5ah7l/ZIxx8VJKBupTUVVTBXyLhadAnRWxYFHWHF1w
6F5PPcRG0Py11YNgPhBWUDRhmIIgpIHXBTWyPD/t8v5B4/6UywDqzbFLeEiScKxRu6JvIW87ROL/
aGMFk2CXM6EFgHf9SHXVnPw7XMaM+8YIctQhSrAeBKGcAIwzGyH7Y33H10gNwqd9/RV5GoIxk5jD
K95CT5s01djcaReTpoY/Ax3HlsB2C6W4Ipm+Oi2rlEjk/N8fAxhsi99nFLmKM0Egh9KVyR8OvsBv
Gx1CQkU43/CUymyfybLdDt9NJ0hyk7hiYpM3dUFzZFL420QtfxUeadpw3VJLBLTSf+P5bj7VsBlX
PdLH/1l6k0b3yAXbElw9gHDu9dx9hIe5UuzhmmX989P0Zn7kHsn8l1Bly3QChCWETYbaccusBFXD
WmyK+31mZUeLo5JiETWsrP92g3ol0fcK3tVN3JpmpzKnKtXpuurYKxnojl+iwQTT2iCKgtmICSG/
RJ+TRtY2REDSI3DGAU1Z+f9/kAnqFiIohVP23vPpNoTDJTwPnaZ9g+QSF2Q/Byu0uQoElpMLbtPA
gPtf7EYEdRT8ymCp1CxQsLPzxuLNPhUFR1jykzsHsmHeW45ty0+WMQk4E+tj2xKqa1qgHVM2AO9c
rdpcC/YiX43koVfoKTwVgnQPayNJy6SLhE4ySZ7Zgc78r1CIzICBiQt2U/3ST+M7e2ITkMSR/H5O
O3/jojJTt2YRZycjp1v7wxGdB1F9blp9A5/dVJEPh3Cw1BSmFCVr9h8auIFsC4f7RRTZTlFizMyD
obbDm3DfjP7V4v6LdwsWI9v4c7HteoWaVRUQ/NgNuxnYQJbDI3LzRavk9M+TDuaVeWYvTUSkIxML
nNMaxR4ZQEA64KRK4l2A5zrj1EXIEQmGDN2Sjsuis86xCugPv9XxAdZV8IFyqLWFRRIdKv2BhAnx
M8EC412Zg+kVU+tgtoa1qQK8wXbXlB4VuTxOzBuPCWFiXn9QHtQ+mUah4L6BRj7/PK26gJ12T4w/
N0GN9qyE7EZ3rLsX2kTr8KiStf3hfz0+HR7TVE6c1KsLgleIM8MWeYsYjBpEDW8zW0VU0Xz5OOFp
6UkYvBHlBt6yayjo0xmH/pqpn6LEBsYVqOE1KQ5AQS0u+qNk+lq4XwmQ/E9qDzk+NaMFyq93AmDK
iENJccX3krKHPWAzRrogxL6bZhh2ZBDZwAXSQ2ZATZIT/OHJe+r7rsD+MBeuU3DNtEFpuFoy8JmH
vuTY+dI+CINMhzQ4pWKyhY3s4VQkXtlRjpn9Nf7rutWTpovBCBrhn5RpfTPSzDLA/TxQxMAmxKIH
GNf61SxvUU4+AJ58ot7yqqj5j2f8RcH9qmXehMe/V01ywc0nYvvEdj2XxbH7U9MtTw7MqiMR/8PI
2vaVEOA/VzdDcwsM9jLDfj7SnYTwfY3NX92Ckq8Ig3F63aWHSlN3NRXKBF18JuYjjp5W1tneDOi8
0EpFt/Nct81x0HCZzGWpElagbLqlkYfHGslsA5GTg+CtCxr1cygqUgbuiuFj845kwPKSpKmodu1D
YeRqpmo4Q3u39m/LBVlgJ31S/z7pDnhw11V6Tg2HFOPcZr4WOVh69zAG/nV2zEo0ZF77hP0dlHSJ
yQSTLBWQjGHn83IP4i9HJHt4aNcltZIICh0iUqQbblmwdjKofpl9dpafJyx9dmBeIHVvezUrLsfd
5ua8ZltY1yFft4UnCYz47ar8gu2w8MGavDJiaT/Z7M92/47VmPVZPlKqMjEnV4TWEOv0Dx1nXsNw
v7xycp0pKx1l6KNRSbyZBR1aXHkAen4ArJ+kqO1ldK9K63dj+zp9xKt4BX58TRYshCz1D3e9DDfI
/n6BDySzDd+vcYcsBT0ui4Vd5j1aRquNI578+kvjNyOSHE66BfSZlMbHVteN4Mi9SYt45zwptHEr
yszVve8d9UjwyRxKVgMe/0I42T7UOx+QkzEVnbHhu6EZFcQjqsuct5AZPlyl8TzMCgqg6KiUPWXl
TpYongX/crP+6+zRl115Gmg7CSTd/mfMjpHi5aQjznQMuxrgOV511Btoq9Q6WQaZ6fWlPrxBBt+f
Om6CefUhRn2tM9lXuKq/kmGEokx6FGrirTL18+yvCU/ITsoIIRn83eQXTK/vVlqY6Zkjt65oCMdq
4K/ln8tOmAleZOTXqeGEw7GKwv0rN/cK6GckjZSOoEum5km+X8n8KB/wGQ/4mdMXlX6/dMa3fb6G
ane8jbVbP8a8MaHD3b8GBU2bHQUIChkIQmwRVhlnhwbW+mV2ljy44UDiWOBE7zBeX+C1hdmfJovC
9reLW7SHHkvuWt/AHi/J5ywKMjCIFjbLd/cIoN6vl8rMqSzdcORAMFmtBoa1QGpxA0fKt1uh3eTV
8NBqoIczrGbQt+JiZFhpjkMnovasMf0qf5725dxxKzuZzDJXWn6+DW1n1G1u/6fjm92fCfaq74Ec
858HrAH3bIggd5VX/wUtwRA/yqpteh0566tuYSH23dQbhNJ28UH1Eh+C5LYhGD2OH/ZSUfWkj2sB
ApFyIXWYxI6twMK7txlDObPSiIghloIhsWUbwM1bsIlRGiat+xAXNEXdvUNhJD16kWZq3F0Z6qly
P4Htmc2h2rkwB4gFCZa5c8TxCvXGyaO0SOYwmmfxx8z4WhvSFCnsSEgQdaRy3sVKyztjug+NPAPu
sbh37nLtVkhZMyAlyMSzC/0dL4gFh+qwbL21/Msd9m6T5Pie8x63tojeK2Wbhkxe90d9M4VfLuvO
wjtzc/BunqtR3cHhcd6P3EwCUIaGdBbMnfv7EbrMGnd1NMeEwN8lmnzVU+yTolQhy8NTunZO309y
x/JHlVt2NPHmQalUyiSsQ6T1TX6qhWyMiR2JrbX0tA/U68xw8Y/G84BC1XMpJ8IgAo6YAJMD7fOp
6NZqlSiwU4DVd2G99Jzyam7vhRZoqlkzCRatdb8vW9kn/DLYt3xFgi5bluwQ6hWBe7xAxcHNOG65
bUlJx8dO9kgkmYaToCGT0XkyTKlTc9n72ptiLxE0pZp17U0qV4TTtfK/gH3qg4QirxCBHE9ESEtu
1yQCFRD2uAgMYFDE4ZEU0w1z6V8mUZ3BQIGJdKIaccAZLa8AfsppUo3iFLpQv1pYboque3EmXUPz
Zi2CvPwaZ3lFbaNO6I0t+Kxjw53+7oBZ/Ax6DoL/nt8Ltmi9liJkeHMN+hvnwtHXfKNluwg5vpi5
CvHBFkF9KcdHJcFK+sX+vHoLWR2FGW/J1JOaGxSfKr5ePoU4BzzgX46h7MpjEYxdwYwtGjCB+68r
O9+ldM6HfwVRyQZTm9fq+oRPKc1hNK6ZY0A8fHChi25iDgvtGNRpipdrjl3E8E7aJjOr/8hOX7QO
FtCtVgC/4lMeeQkKEWsjQwgB1Nd5u8E7eAv7nNONFvCEnZ2HPDXgUJTJvpdunmuesCVQOcTUPAOV
P6e4toCQRvHhGQcMT2Og644wnLetcP7BgVMJrCCTcRq/ZdfVIQMtrlL3Z8/fLWyX3l1cCoBQ+MOw
/mdseVF42nZutU60kgouS+qzn+8o9GvM3PKqDQWYHlJZ4oFiFVfS+PE69vK/2AWJ1lChQByVnr71
E5zLesQeuNGJ/JBqG5P+9EOxdZT+1TCeRu01I5f8SRUdkIuJCFEn5cCXKiqz20D9WDuBxXj8MGsU
6BrG2snhmF0Fe3s1fiLQel+KxElxUcPYivsRP2jgm+5FzQXNcYQAdCNH898eMB8dC0RBHTTmFZb3
xAjlrO60pe/wFIWy922RHJsMLKRS2BJ8tFYQtZoT/eJxD9bXbb49teQ1O8jCjtddafu1r69IfNI8
CSovw3haip4OzeSxuAXrjemFF9hkAIcVbX5xoAmJd0slsGsYCrK6CY/OkSVnbsjEIZ+CCD5qh/Jj
sBQkABu+j4P8CHvaVYK2J1Wf6Aqp9YV7h8bVfaabZLHhg9c1PsIGEv0PIfv9aMsOThiDHZBNfGCu
rgkWJdX2Es98xwCYO7rjH+l70mee3qBSvbxhi0gGm3HFMy3qqZp0k8rh+XU1fib1ZbxaY85fvqE7
wvvXYhge/YvzLzgFnGHvydIFygxRLvpG42HSgE2cXz/XNJE4N/BVHS/0DwzSa/y1a0BLO8WGBTvJ
5D2o1oYc+uB/EfUaTyrh1doK2RT1LitrQnVKC8nfbHFq5rgkVyBD5dsl197leA21K+zZ4e9ADSJy
gWkNzqBeqPIPDUgFO5WZpO8XK6td1z5lq++JxbUIXrsvxp2D2BAMuonvwG6OVEwvuAHbzUGddmbh
fh+6UVtis3Ie98S5Xa2Fepfgi5F8dg+CEMR9mLwZMjgVkyzKZh/3TzStbEDugcw7sFte8HlmjrxI
H0+cHEDOuLKwcVgEf51sYv3qcAN+vdoX1YJFmY4yLCVMBkCozXzjlIUwrKEYlSDOtQoxl7cI666i
qgOD+GvQF0+w2YUPbp9zQn9UDGJFRNdQi6nERn/NuxOBUrR0E6/tZd4xg5g2MjnlQY94SuPmzKuH
gfgrAxXyqV6ESjfbw44Z5zkF8Vlqy7DMMUUVB2sTxhb9eCVeWK1Tx2AtiR42sHbIa4lqXiIsio+/
Y6SE1IL7Q1z4o0c6bgsNfY3W0QTjqom7yNOOYFkcav2DRhu15RXqSpaqUEHnrja6TFALzkSqKJVJ
4GKiSCSDk5ToOyqf0n2MQFEblzE8ZZHlSQro3bXrUHHm8/LxEoqM71gtNu9fnc4WeTfiSU6ebd5v
/bHdpEW41QLzpPHaxgf25RAFJVJTZnA9ghkxf2f6o0cGOu8e1je/tymYAyUCctS6XG3iNV9QhECu
jNB8lKzmMGEioAYJvN39APhKhiIOez2Cjn71Z0pwUIBgGhxUh+KY8VXbGrxcr5xIw1B2Ta0Kltcp
5KGKV5GGMitgeBSGM9u6leSZJuFeugdkMrf8ElDHMHC76kU/k7JB2Cwbx/akeNBwUzXkuAv0Dcsy
Rn2Jg+gg5u/Kv4x3zO/XZubSTuez21sT5NLd4Rql2fxt4lgsEeSHN/GbF+IK0apZupJH1nt7P9at
Fotowg4lF8oeWkhPOnYA+TnsJo5Y+TNg4wo1fL1fWQc0BgrUx2adV1cMzQkth7NYuntuiopuGkby
YlAeKw3EDGNlX7nlX9NjaPD5BfA0KyILUt6z+mwPrtkOzGOL2K9WuKroXPBDHNRa4g+9XgTF99a6
wwi0oTsYT/owgaz+ZdxypahIa1gogFkqwv8YI6i89TGbMd4quqrSBx9jKl7H8o2vJYZK162FLDMM
af+fmOJqh0PUDwb1RqxWcIiE9bBe4mxugneTLGnHQAIzByrC/Ur4f4p677ZxDvmixSeoErUJPlzp
Kzs2piwtMjRm4guFDK20p/Bj8+fqcav5EwVWIIuzl/3x0MkNofimCGnCCeHh2uVCNlU1oYofuDph
yQLCU6MGqTusTRmevTEbvRLx8zDUsDBYKTKrsXnqkgymx4ek+w2YlqbcK+WZE3TSiHFifxjvEyOA
Jw5GufCaratHs1KmQ4eOhZeDOyTKVYRuHvOVUoxwyYs6JnExbt/Ely1Bt03g9PfHhSD2uRZO2TnS
cBh6UXvDUuypXknDW+zs+AXxvrpbLDkVh9WNrRYflOCfgGpXfH6JSlOohjg02IYziZPtToaqqXxn
J0RMxxA5lV58LDaE12osc2ea5SfAW1I/mYlUb6rl5Z2VdxwkXraqVpUT2SR9hYq7LsQ9aVnpR44w
io7greh8p+HUdOgJo8okLSFisAFP4+ghoMdOlp+Y+00s0uD/qkPCLC+qYuvVR+YxJ4dghH7BxYpo
VbIcc97mh7ULf+XUa85LRbe9y/c82l1aX1sSbev7Q5o+T8CiqGgqcsvSMsNyyZfEqcO+aJh94s8D
8VJEPFK20/oqtBu0PE5m6HFyG2HfRink/HGrl/YS7DPHajB3mi3B5nZ/N77Y2f5pqWpJAZ7rNSgR
hsWj262nJvsrUBVKN8AYDqK8aX9UBdA3ehAdNbMEle0qkYwL4v+ZM8Xd5KIPb+fsgR0VXA1R53p9
SmcgGUGd3VC4IbtymcpAZvT/qGdIFJTCNArHW3m2yls+Aq3jQE2iR3MzxDQqlbvKug/WnyvWG5ap
gcD/i03gL7mXyb1nZKdSsQczcdb1cwN3cXzbCuqMUb5YW76epZ6lP9EDkgkefXccBFY/yqRZWgv0
kj/fPB8fY1aSowxKHtJFpOrh2+3+2Oq0orFMY0eF2jzU5EEWdRcHnMC0aypYNlXktw6BV1F8KxDW
vSIvv0rsb9O0C5P9XJ7O0Q8yMkVwGf3kGQMwwSqgoSccgtH3HSm57dfBiBX3Tp3NbxNyIH7IQanX
EOVS/2NpizqRbU0fZuDNxUhz2+3jrfe9/JaMPl7mjWV4PK2QLL4UZdARKimqFCQfnED1OKW+UP3n
NmrQ8z4qtiKvD2IYNmyTSOHU1w3ZlUm0VLPGQgyhEBBygU+Lc9PSDSfCQAk4Z1slAQHSMZnPWPXl
0l1NbJrBx8V1VRpE4wFudSFtTg4s+eHNpUqGFo598EXClGvrASzUp+MnajUtdj6BH1QDzBN+xxgN
YYWM6UlFo17h1dZHs42Zo5JBzLz+LYWvCpHF9ewFWREziRPVvFp/zxxuK7qXHFBJ3H2Ih+Y7Y6/W
eR7m95VZGUdKCBfN6J7cde+DpoPIsCgTjt3eJjW6yGbzEClfHpAJa5L5bHpc00hpyPKGYCCq0ezT
N986C79i2PVC0icFjoFZxeqn7ACRuj5zKhYYzn9bWGmxDKk5YlSZKwNofqMQ0uPUdYg2Vwp5uAM8
T+ELLnePKsWtfhuKFCjOmo8cpA0a4l9lsSnMYOT0JGJUhl2rLAcKn6+PU6cz8AnAkgUaCC61EFJb
fpEQZIr7pR5w/9vBQMQJX/EnW/nS5DrYzYYeGojGLrQe96rxBYXgeMf0b7zHe04h1+1hIoby3t/3
2x4PVIjYixR9er5YL9AwoFLiytu4+9GkUEpV4xD/uFfnDjAy8aSSnT4dCeijMru2yhOe1axW43I6
QAP/wRktyLxeoE6X6G6UbHIIkkKvjSjj0k53JQj7bpc/dg2jbPwx1jFAC6M/M2PSj3WSh96eURpv
DRLoFerrpORn+Xgp4EhgFWFjeTiI+FeB3dPI31THnD48YbO9CMO6MbVqKuNWKwUipsFf3sV1s0Tg
dSz8/IAE3o224mqYmOBfCRs3gPICmVgPirpx7BUtNURqRkOig6+wBy8QhxF8MEACerkLse3L2w9H
FGfrQlYUZE61Nwrwv7YOiwMS57Emz7Qq7PcXdZgWmaoZnXb1oVMUvFJRlxvkaKkAAT9nYhfS2DFw
+0Wvki3+OpcZsYCzYZwAL5KshOzlwXHj6iaDklJNXQVX4bQUmxzyKavc7uFEigYqrEOi7d6ncDSt
7U6wqfhoaxmoQIwJHvcxatsaWR7nJ66Rq2oB1YHkgI4G8ZOXDXrOJOcjWoXALRNG6tc3xrouPGvc
dnXjAoZ6a0345WL5lFGRCLqcZLo8CqYNx95MUdi5gygQZMD+HqHTqmltN3FdPBK0AmbjcEEagxb2
tb2mN+YMvJfyoswqvAlyzTfBXhxmgnLXmC3fKU5o5pUpcAuzsXDW1gMBUQ6gaTduWj0hefkCiEcW
5m/cdOrQ2Ckhadm3Biktz+U0MTHdPY5BmkViC6DrZw8U0tt6Z2a9k82xfeWdTYk0vYMzvvc3mkLm
PR62buyHzxTMJCMB+wiSMMwzrvKLgT/04p4+durM7Md58nkijjgovBTybgO9gPSt/f3jl9jGdQbO
xMfHn0aOJvFRVZctwJN7MmRQeTbekuSkWPWU9HajMz+yI7/JOR29SNwxae6VInSP7TlTYKddRTsh
s/Jnrx0MWRo3SSFC9QmDPZN/jjKItbSwFdgaDzbft/lfIzNFvYVxfVB87WMN14SNrGoFLZYrxhCS
XO2jr0+1CTX+qSaV/XHsO/ucPGVmLNs1U09C5h3EQoUZFW2JxIvMi32N2fa/+dhmTgSeVmESNmXy
06sesZTRhaZjJCOMhxriNa/e6tsLNfpbDXTlmEHyD7tOLYKCGgPJvTZZyTQKeBXKPXRMrmmw+4Hl
8MVcciijTTwcfJdvt7hDGosFEIHTFXEincmSzixCF2MQBdg4J1DT75hC4NuPczUi+XCFWsuTM7j1
v8fhAVVkgHPG6XjikqXIxJSQ7+kr3GgTOsgnH4HwlJUuyxRHPSmZMvgb8ZQUR6yfjm2bMcMCbWyE
LRBQFMO4fd1iO3O+worKdAgxVGGbgUbYzOq5Q9EeiN6g0xquBHEvymfqNs7JVprbv4Ry8F02Mn5Q
fN2h3SMJmnEGsITff/HWZLAslxtDaSPYBVGktAI4GSoKA/mdVpn4fD4iBm+0S0xljKYkRkbOP/SV
gYja8zdYQuKOEFkBZWv9Dx+CmqMQr7ENZjBOzk1Vy6wrzgLr9Q5Mp/i6rPtyuQtSEIH7LQHXx5cQ
iCMP4/Y4F8TryJkUR3z/x9/0xPHdpR7iNXVocpCenyO8FIPHX07wFwbKm1fxVHO466N9WBa5gnvA
g51pfxb+pPRWiuONrJpUbHlFutjsMqTy1fwkeFCsCa+CjhLRIS1CWQnlLuaWarWdiH3wpcV84pSP
+kTz9dQVT2qUo73Rhq//V9mA31ozXBe3mnKEJ3HbqeHwzPwZcouchaeaE62cGUZpPeUlXm22EPtN
Wcfu3JSohcEirrjKKbpWw/90fxLRUgYPBep81F2dVKITSqkMTAC3Qifil1buV4t5i26RT/BWUUh3
KxHWO8PDk2D+ALYngg0oFdRb/vosbur27PH9fngaOHnyNM3g2pvTXUqaYOcvd+1I52iWzrWD4EOs
gCtJfMnWVt8mJxfqUO/P/LT27/b0VtuEOJvWKMCXBzhl70gjgZKAuYii26M/AJ8MNc3PZIRCwQXm
4T0WFAnmTJPJ7T7NzvLF2jUXjG4TVaXUKiGPHuC+YSK6p22wEc522nvrniqrc2OxYCUx8ORO2qDW
guNsEt2sPAdVWa8ZMuhfxLaApZrcWLn8yOskcVdASivw69qCc4AdMUaTh5ND+rtmALooqGuZmTnZ
xiygAXm0xh+nxMbYijkPUdU8ZEjxaXUSOMmwK45Pujg+efD3e1h9nc1n54BXQD3W4FKvLMYzB3sz
0fBqfIi93j2GBQeCUdGOCfzvYOj0jXSh5h8RKiEgpKNV/n7+9zLvnfYNMDVyqnXhuNlSJiLvRs0m
qJA2Xe2oEoxBlF02iLeRI4m8Pna0garArCwfsLE4XWzj7F1RMGNhTK4WnSeqF3x+EzJLbbFV7rj+
T46lfuTXHkH8ye4YVNTtdm2VpkCIgip2YyvY8esey5hnWOytsbDRco5EoK+x4Qtu59UOzwC4vOO+
em2bL9lnKng7nmV1cBcSGNhJm5sHagKDXEhH8OoAESR7JFfcZnoO2VHdlQ5aarcb7gvTXj1MUetM
sIa+GkZ2eZg6+SmVjbUI3A44gPKIIKfoWnAPo1NR/63j3/CO3+itvdtz5F7368ajsHTbC29ui1Qs
pvPKQsYWYDrNJnsjBLYhxX1F4p8i5UKDPYM+x4nzqWebfEzVC5VtA8u9iYM98I92AttZEGNn5oPN
mBgulI3NTZJ2hA/DhQKk6M8u86nHcqfXnxYnaFaNUPkWmRx5pS/n8RhxHRrd1Qc7sKfUwJMYPGra
P/bFyUgRxwW/5KcH5Z4w5472hNA8YbnQRnOf04JWgFR1Oda0Bg5BkvzbsMZ22WnOQ0Xr0j2XIL8E
IQXYeZ6WiZom4PlxJUvXirUqVIpW7j6d3vORMGHrbU8+0VjPjfAA6DNGca6BRq4jYcayEXL0yHUZ
YpmIc7K+603L5BBZBDH0s4okKUTECKWzNoDMiyevvtPCcyjZPRTHCjmkmmtG1x8AwdZ6896c1Oyj
pmmeDKYs10nVbdUCNtkEQbkn7E+3JxGn8ZtiNEOcEpdpV4H+lwAFEOddMEAw7H6JPRnHHx7TUQL7
Za+yPxVdeYEbLHyprZOmElp1oj1x9oeqmFtLME6X3m3IAFPm/M8JEYGSBrBfIOJOshkWM9B+Qh/d
MI9UuFHzLz4M+vXdyDYxnUF7r7jdk1xLNfb5R1F+oeGD3ZhxrjMKylKiWpFgaxGxMdKYlcd72oj+
8ItQJQaRw2flDXW9+O99TBxgukhnVuS4VI82jW7HwPJTeF6YDaHPRyNiX87V9wnw+lwnsLDjMLwo
5J7929WAsMrIvXv9GaByDeSN+8NGuR7Gn+tYx5WcpzOvmH02Q29MU/IEhQbrYSko0MndATZqzpQZ
zMhtq1YbFTMOTyAgrfTGMV7e+3aeB7SsKwE7nx1FVqo9/s4xlnmSTwsD7hHgziGEPMCHjEmNCd2o
VqTjRe/+zxg+qAI56alsQM7lBmnzT/d/O9MWAKpQVTRHT3QNNpr/M2tyGmou5EJTDNq7tZf8pTiz
fYom2c4u6LN86WcDNpR6YS4fvvziVTkfK59zubarJNij/BvEty/DkKKEldeht9Pc513KANKxYZQr
Sfc2qwuiS1rAa3uH1sPkd9OCEhHxVg81oDHuvgkJwOdgIBio5QXTaIfakSburF2jbEL6fsJxVjNQ
zB9WB6me8Fnt4nBQhu+KImZIjVvCv+1gxQgJVHei+Gf6AeI3EOAEF8jJ4JD/stGYU4WygwYQ6JH3
/pYomBsLBt4VISGV1cQDYaA19qMg1u0g3aNPdx4HUTQoxtkDFiwj4ojTBnpJN42n1HaDd71TLbuR
/1ZLSdopnGHm/asnQcmiAkT0s4FWETkoVL5e5lODbX+N0olOnyPqXjsFH5JorAj1QaOhLCcD87tx
OaSrwiW17cUxZ1CB5WrqqVqbJ/lAUx/F/RHu/SOk7smWS9rM9ZY+qLlIIxGBor3MYhCGd9+PM725
+jyfEkyADFBFDMgt5fm5YE6RgJ+QBPtHRQfHknQBJynCpZMOwzcB8WK6RIxKVtStNOOr3qVqBUkC
61aYkw95bef2VC2IwJjrFClQTJPOk+1xW2+eK7wjPvyW3vUhJ2ET3TbU/VISSBMWvpwJ7ZRek7tq
CU/VbeE4Qev7dXSEVEtACx6q/sXtqDAtD2FbzN8X6N2nJ2mM0AStnQrpCWj5Uewzdtps4q8cxwXf
hCuGUo4nURbS+BeYDPW2q6CSqw993rKv/16FOES2d7UkebdM6Uxl2EcOkZPSyVspacXkMM1eibpO
WeiiarMi75VD9CXg1Y2s8InnQHOPdTgq1Q742Jhqp8wy6y0ElmbQfFXbZMpO7g2rONgwY0nLrM9r
R76HZL1TRFX4ZtYwbKJHvKvqtSKcOrQVk+TBlR+bq0x4Io7jkHOm870BLAQcYlzRKenaq6wA1wk4
uuPNf0++NgHMQs3xeXAxUERvY+xX5zdVfGI8xk+GN3Mt/6oTaraqUSZapwtQwgGrr/a1Anec+3/U
0WvsULNcLhNo0yXanJfrFAJVUeRLZh0AhBe+NhhwQ9jp8P6pTQpyG69f9meHC6EE5reaq80MGcKe
6c2DEgaQ9z3InmX4NqeOguoIcY6m+Rxay+jJxhawndHA9vkZdxwLWnsQN5+e7FYQ0x396uuuLuY7
Jupad39F7pdOv8I3iERWWh6kF1CllMdtLYhZ3qtnpGlkK2X/Q0hJm9ILjcOkrSgr7KdkjVcD0ILj
5o6vTe2g4FJfDw9k6YluE9HRMoSAiIY0yjtWQZ5EjDXMJyYafzGI68BlNL5/fDYZZyRDBZqzNDH7
pssyBWHCj/mfFupT11FYtxyMZ+986x1D6AYAI8iuEiP2msipOb7vVzksvHv80rB76yPe3dM2B4IO
ZNBp34j5Zr+0pLNYspFuB3j6yO0Sl1c0vt9iKS4hd+dSSQVmHZlqOYrRRgc0sU99+h2dhnlBarzy
0Px0S+AXwY6uALQ0+BI6jGYU5YGyEJenbs4l5MW6chHfo2Pz68+Y3Hf75YKaTXEGqN8eiUCZJNAV
XUTNvUyEGFfBX8ee4fXZHtQb5clsq1ZJHdHbYxJkKAv5NLpe4/B6zeKRC7neGZb0Y3WbnsK5e+Ww
07u0/NdlJcFS5D+rz8z/p2Q0F8frtT0UL/e/iKOg5CNXIV79x5QugJXX/FxgLI/BrRJq6EOwV6cr
wks056d10D3KAEzYnZVzLKwOs5S0lAHdg9Fq0dgJRm1F6A4gCHRum1MzvlNMO89MbAOsWUV45qm0
iufuV29ZcLxqbSOMwTZpzKZGX12l8Z1xMbj0hAusWzvzOeafPrwBcN2pRbKVlY8smrgcHYQlcuXW
Gq+w83SywEYKYPycrUvyGDfRiOZoExSoRbDOZs4RnsOfnZBb1vw71Gahr8X2tBkSPRqkDs5talkO
W7FDfqNtZZXDzQcRD/TB5zMTWbDHyWiucmUh0ayA+/5S0Uzf3zum1UvWqIS2CF6nSpn+ZvPO9Wj3
WNtu6JfBZWXRQdJ8pP6B1R/iOCXNTDy+H8lG3DhDPRMkx1RuHPd5xt4aWzYDeGYiM7hUgHDiCuN3
BUvhAnqfZi19CT9Nz/TXiSPCU91gZij1NNSN4vkroJ8CRApqqX/qxVnhJt2kTwVIHIFj1fhJsLic
9S2fQGyEpebGGOCr4fLqVAp1a6WHfuCFNxDXJY7yyMhO92Ca9hgQcGb+oiXBVtqVxCRGPANLVxfq
HYw8uGuYK8ivue5V90bqHh63SF+qCcQ3L6N3AirQUfq9KXKb36ETjE5W4tbs94iR6YXPLx37j5+H
0V+YO8gDXBZs/0nvKq6NRBq65wN2hqtCGKecp3VryGNFSPCuvFRhQg4MJ3cUvMd5fb5I2WPN5Rc+
+Uw2Lm5c10sJceP+1GuMd3cvTOeV8o/i2XjKnFE2UviVYDXp2nmWFT+JUjQPwVNLypQIRG2mz56x
FHsvbRbdcivMR43AJIQdT+h8fycUxhftvvjikBhJH/nfIq5vYJ5Og/Kn7knCIyrVKLm0sM9KWTr3
nms13iJOzIFPlvVRUd0g0EpzCkgyQda97JqgaxMXC7N+RpkFuLJo4j51s5GU9vQ3VGYE9P17Qq0z
WMixBri756rHXnMxLD5V0ThBtUONGKoGedxPPSK5M3qtfSoZxwH6TOypUrQ8ne/oKN8ZvZGBDYM6
jtA6H8uu8JXegdFrgPiPd1679LKJYf4VUbk9aY00w3Lw30Js4iWIXiNUZxvXnNadkN2yoDe7uUgr
aAvZT/YmKhLqjvoBBsE8KC3b4a3QHj8+FrGcbzl5kkupD+JcqFSIycABIuV5mX/NBS03/FuR98Mk
ZvZf2qocX0uFVv4rL3PT8zGyatej6usiCoONCbnvPxklVy45AeOVR5d8GoBGmJvidJFq75Ldyodb
IhLKiICSfVOFtkpIiulvaeHCcb/d9feaVopWKIOYOPK3pVICV2ejqGBeUNuabzOXcxhkiOv8Q47X
xUlwZDtXWKBr9JRrOOA6FDaX5MKU5HWoGghd6ovjljAMGQPrshSPTFaO8SbohBQPFiS+KpujtLva
fknEK23WVbG3R6fELX9utoyiqgvf81ut+LhO5UYeqBqd4aw5j9qIQE56uAIEvJHdQ6KInk7KbKQi
7EiKUHiCnurlE19mku8oFz4wHT7TXutd9aMQlHZ+mZQJ6p720VFFGRu8RhK4aKHv90ujHX4Zd2Tg
9RniZ9z1L5HYpklreJBraSO3Oe+YdYS8tt2QkUGfbLM4fA0PO4jLUHdw0zBQChBJertBEUMq8foN
eefZ6JEJ5PKBBR8M/FmJXRE1vTivm/u3/Zrxo4mONnRFcEjX8ui1hj+j8mzwYylGsqbQGgMRMSlV
k2yv7+BqBBrvx4qfWTMElmF1eYuf0t+qNnh3zUG25qP9cMZeh5BhAJX905t7BewTiSC4y6VB5O0S
THqswMjl4yt/9rzEtQ6krJU003Nu2UooZmdUVG0SJkHc2bk05pXgAGSJMHOGb2uH5lTWVaoqkRdt
q+PyHOF5DeIT9vjypXlhUHJisP3PBbIanXnRy+3S9L2FBG9gSK/rmT5UPayFyzUn4ZCJmESYKUKg
EemdONDHcHM5AtgZW3dbnkfrX69dq9c1bk6FTYZ4kYnAOPR0wk2yjvGCF+Vlt1lpqx1Ksj3bCbnf
MyqgTEiGRcNS9UfhzUcM+028P/UJLrzfW61VWnBxwy3vinCl4JWXrJcNAYiroAEJ1VDBS3mpKSj4
8HUTqNC4fx1dtfBgQdDp2S+D5DYH5hJHVayIpbL8r/uh7xGgENb8641v9ler+DHJ4CThRO3oJTR1
Yp6wGgI/QtKc4WBXnLoX8cWFMtfXUV7Nv30YnMnwn4+SID/lfYDIImkRF6ycVzHR61hi70Ms5f10
CFWD50pMQOq0lAHBWjRsX6bc6rYmFuzv8Oc4uiGJbCmMBWFcZOc34bRRq+arpgVhZkL2Et/hAopc
IokYM5uFPoYx+N7BYQKdDV2K3UGaYghoNvmW5NApUyZLrX0mTxdKdH6xiqTgaBeAC+7cx5vOw6Px
R85PXAxKuyI0V2S/La80Jr3L/HEwn2UTzjOO4+jiZAORiD5GNCSTMYKAX00c5iswcUDge26ji98l
yWXq/HFQfTwYbTvJhOmOhU9OqvgMMhkCOAy3ZlPq/uSp7xdhMMNq8PfSUrAnEXxQQIxQQ0MNArC6
vRMso5Oko0intHn/ft6K25tYJueII3mOl+NO2igTElQNT9ReXPsKrT5f0ucwKiNri8bnEdc/NvAe
afg1KC4c1FXoCYX9NO6OOz1dThHOPPXYfR3AA5PIp5QPfWRyXscXe3wJUumFTdYWKSEZgdKSzVT3
9KqczmRtv47DVlhLqrPuIkomDOe3MWa+PotKe2MCqu1R91feJGfXD4Rq+r3m7pd4LqcFoB/ke9ft
e64LVDcUCWXuGVeMCfTuDYSc32GNo9lL27htRscsDe7ze7Q7O4gEqZa/SaKvdi6yj2BNB712l/Jw
gly6IlIDw1Hg+Uht02skCOqqPrJjW+E+HzYLPAx9QnMuLK3iIq3ZdS50dxfS7k8tH/7NemjlfWea
6rBep/q3HmNC6kUF2emDmVwRNCXdi6vCEgAL2AOMigjNghleA9+CzJ/CZakEYLB5iFQSM6pDIHvd
0PFpHVPpTesL9H3HoXCWYzwppYE/oB5Mxf2zFD7GhLlTF7z/G17iH/k/QkbOm/+Jfd3vOqKTPPUm
8EAV2LqHWZJEQMT3KloN81rC1ACz7boyPTACkKPd9ZkqHdxW1OOjKAGPIZsPSfB/Pv469PSgfPQQ
c1uKhYhKK552rl0UHVKvmp/Jx5Zw4ID0Daz+4DCrwI2YNanHXVVx/PiczEeSWB5Ft0qwUUyki+6Y
W2lT7RNdZLb6p8Wbw6v5LZH4jAQX5IKux0ZvUHTgf26YVMDe2j40pkvXZM07A+UR1N5j8KDoCmoq
UBPjUlhcYn1Qkj6CaePCS/oSB/EUVNoKcHkr7XRvlg4ek0CxY/OT9DyFboql6qY4OKgSRpZUtRC5
feScpkG1YxxX5Hzjlry6yccW8+oC+2rh54YqFLjLtpw2rQotC1P0jOiPrXPp9rlbCHzEHO7xa14R
fSNrmYJhRJ3DtJpINvYLReJhBq060Wn7+8fCnf+3Lv8tnjPkbagAzkJHjt00cjf6ZiyPb0vyhi6r
qSwtXtykrLTH9wKjEHW3TyxMKBvby/YzG6hgQ92ftuERdWeABRMPEk51UYR1uY28CKjKZQBUPbIh
j1wxBDeqc9hhss4E+Ve3Hcs+2hUBlwghWi2qCd2WeY66Z2m43l/Uzw+6BdwCetwUpBJ/CVN2ETJq
JI0fJUfGQXkU02yepS1/NLdSrSOZLBxRZRaCcc4C2nftQTGDMmmHJhD9fKjFkiI3wljJMMEjQZpW
1dPbu2rDdfNat7bBhg3MeAgC6idWkWfv4wxdEqeGu98L6CYM9PgBPcF6dsKEkhMFJ1nrN2Fa0Zoe
q8zH43Nx5jtGDUYQFlhhWQqFsbvYzdkY8Xs0KH13vN4jnwkug69idauzqalezZoaHPx5iN9cwnGG
TVq6nWwF+kBP6zSmtZbY/g/IVU3zUlyHQcb17+CYCpt7lJbdkFkOAsIN7G8n+lVjE5lYkMV1uHya
4AxCEOQb46AsbnhC81oWhxW9A1aeuiZb6Z34dBl1619Ubd8HtT3aIRmQMPJq2kuCK3zP5ZVQz0ox
jt5tNzKrrsqj4Fo/sP7STditZkZIoom97wIyzCkHIOwFbm46Aolrmq78EE2jJWFS2ebTbyr7G4qL
D9ZTYqzQ3MG2l7eK/GYmglSWBaiz2VFwlrA5rqKuyoCQ3mKqJBg6TWe7s7W0+IB5CTrKUV6dik56
Up9l+9jxgTIIjwXo3xLjXFBknW/f2i2pUoJyvgtFajCa29VeY39j8NIRKOa8uR3uB6at1vD7Egsk
El05PjXI8orxkHaWVE3ovSfuTwZ2MLarSApfm0GuWqTZDqeCdZOZ0J+tZoWVWNXQpb7g9D9uYqTI
OK3yNOQzYrcNLnvAolNHH6m7jlrbx5l1Hzvr3+QJRlmGtpXxmRuQPZlwG2PMNLbhyXp/XtRk1h/p
im1niy2jbOjjUd9UMPdHxRu4A0Y9u1tToqKCgn150E1PDL3gZHmZofiD0uUQ0D8TN24MJibJ/8JI
B05LdFIbViINJMiAaSg40rCGbaig8hsbSoisIRFoEy1Jzmc4V/LmqnNSAX3y+Wl5lVSz3UsRVRtq
B+pL6pgfrY8tC8TOZEwyN7KArLjYYaRSkV9By1LnugB2T1vh+QjX4ChKYQ9Jho1U45MhUrusQJKb
1Bbc0P1x4Sdhl80LLVySdt9kA6fwWSQa1ZdmQJ8IA4/hW33QA/OsnSooDzKDICUhaA/ZL+2gMmmR
+7zXg7hq/COliJMYhb1IIPQVXVglWpbGK6PJoCqEMLANIbhdO14nVbHrPx/NM1cd+6aKZvILXskw
911/8UcyRWazUWpH8ohVNDF1yEzqhUcQCnWmiElN9in9jHGYuO/Eox70dw64mAhoWC0dTLy+e4Jj
zzrCFmjVmAyKQr2GHzHbP+Wf9fxQAaYg2uOaZRMZU0Ugesxe2cldvUoRS0/h9R2brf5aveQpNkev
I3FCkDz47+Vk1HaMnwKDhw3X0xdViy/mrwbE6S5zP+VyCKrn3qp7C8E5/IznoEu9ZvYkuXkBnEGq
BGHexcpXnCftzZcC+qCJCm1hapUcjc6VlOSVQQJeAFE+tQr2Bz4I7KI3JDeANIy62sZt7lwh3Ze6
NzjwmZIL/Sw/r1Ep5JS18ydyI8NeOEnaYU+6GtcpiqNByEkPZXerLN+e6TB6C1PcU/1EmaMMLm51
E+g4MyrOKFeCZY8KKvq7KIkwas1j80C1hjNMrGCx9c2H89PUwBn7moekshWYAfylNoRDhDtOvTKN
9ra8gwfjMyK9pgfMYExfQwYEq3kGZYdLXIPer2fY7R+e8NSmip0lBY4dkATSU8wdAtELebJl2e6C
Fp/zl2u+y0GIhVD9FeNhV5y7UlEnSAYAQngvi8wkZASgKQXC+sG2wEU0wc+AVJfSvN85qNe7Uhot
UVp9Cx/BgoPdYPloclTKZnpmI4wmlas1dW4al+zSC9vCm1UiysvJ4bUrICDvKKCyifs+5O2i9DJX
3RxmIB02/Zix+KziGduxgMxjL24mcg2lHNejbsr7lJcqKlVQvREoeCLdTdL271kID0GOq5Bf5uEE
Oe5cKJLjlzN04ykmdsnRA/vxdsSsPJ0b2hWVbqnwzPBe3f4xvWGwaDJeKW9lmDmrmOnFCSNDllc/
e9+XLrDlTgP+4S/uii0B9Q/RAYsFuw/E9FJSad6jx49gxMtH3+bzp8dMbGO0B9PdEEEwN3vFqZZo
R6fXbDx6oOvoOX2bcMFvVjMs+CYWq2UFz2coYTZJI9izBkMRGo07t6tmhWy0p7DMHZ6OYPca2g9J
+s/fh2vydswuhX3cMICd3qeMvirw1ErW6vC6wOXdeYe4sGEGOosIPQU4ENyppJZTLFk6m6eWovje
6EAHJ2dfFAABcAKdax76cJRJLVyWIZ7zhk9C04vdy8P+RAsaam4KKk/XJR52thLAtkgfuYlr1G86
K/DbNpzZi9QB++95eoXzeAcuJSADIUZyRcAjIv8IoOngnosIGZ1iPgm8Jk89Ji0wjD9NOQ/jhNM6
swAQppAznZBGmRcyG9FRX0+BDXEIbBckaOwjgkmQGNsCI51/PxYc+Xon0owFGr6AIb394hehXaYO
EPUHQ9pQJ9t+8LdWKWtoc6dz0XXuhgBVriuS+n6I6xZNj1EiZ0+f6/MQs6P9HtUyzu2dmTJYIw16
wULhMzfCTV0NygDLZs6LIG37lGolI7Mm13wfLdWON2nwRHMha0KhWbGcD6z8+JLguJMSomp5xF9o
I9+soxPPvpPfEsuW/S8/+s4c4N8ZoqKPv2HXx37LRAdM4FLFwOg1P7JduJ1ifu5wD01CX9VJyvkq
gPjvduJlzFm76fHM9Ho+oQH8a9I9WdztCzop+SuFaArw2Zy4MNEWnKYTrFBBpmF9FggZOCzaM6Vg
S16Eri1AS1NQpuBzw5vb7X4B6QFRSx8bkyqoWqQFEaXGscCUe3EvvtIma2CFrdlNbBEc059LbdwI
29+1Wt/NYXJyoLOW0xEZlASNf2nPgEr8SMUSLc40bWUfx9d01BRuLhHnKnUGcx2zDFwkDmMM810J
myUPbdFVUS2hG3t7MaMXSA9gmc3rFKhy/hfF2D8wxUhApGf4WF60XDwjTeBhNl1gG6dFM0oUEGw+
yt+R7iCw7COTYSEsP8lvDXEfRkmSFYfoD23Y64enLBM6V2E/+LDaYpNc7kNnF7ZonVBwz2ZKJtmz
mYRGh8YrpMTjxoxQC0/RmiXtNiZ3cU7PEVrcDcytD39q10ZofUr7aQXhJ7ekA9n8NKdx+VIOz8C5
uUbRwWUIyPDHsxWZPWfukpIrakTxXZz647Ah8b3s5RFXSH83rdYVc/inTq3giGfDPi9ayeMs7QhG
GJacwtUKdcbzSTMjnf/CjCp/x5n6tzk8WB2iCGUruWtzzQrR+n2Zgy43Nl7naGJYecXlMo75vkvU
GtOHhUNT6naFvSOl8IbabRE5OY/tYnzFChzkZff7FxDSIUlrqi2RrtrctLRKA3l2KUoJF+AqZtCJ
BP9svlUpKelhPNBFPXGZPwkA8IpReylIK+8WNMZfdtPsgknIdanvcM3eWT5GszdpNaicFELP0zmY
sFZeH5I9VyFsimkHJUfFzuu6Rqiz4XoxyD6woC7j+BslhcwWSdejxah08qJmirXkeDSbUSIuwbjh
ekSR4NvkKi5ClXI4qfn+0oPS9SDghxQc0eG3LQKbkLils1SLFrdzwZeb9/y/DLpMOQmiw1FhbTAO
768n7MRwxObg3f6tOIqgnZdrT6ai9K+tRirzHK+gqZdk7n1vVhH2hJM9UoYS9yR596kn4zba5X1c
tpPOLgHiZ35Omgebp4SsbcMcB7bJVjk0WmGE648agUxY8/Mo2jI5b0c9BZS6K7myPgGZIhVdR44G
diEQW49QYSWvu74GXKdweH5uZ/E8dtVjOpCMb50VtLvd7e3MP0FS7SIS4Ss0D2jiRPWhPwmlH1Fk
1nV0N+B3/P6Sl/Lw5JhfdfJ3UyizgRCGf1o3BdId+xCyxEg5OGCHF8byf4n0FM4uRwkUzhlYnyMf
qzIGtvZz3oE2B7mXooFSlCKmTJeGZV1HoA8j/PPcwtWFYm5FSyajhCshYSdsyW/hNhpL7V22u8yU
MjYUYdhHR3/U43/9URO13UF+SBawl+LuhPq2snuCHNusOVYv/AKcOy8cNTekCOXxfUX1S7VL6V3m
t26dXh6GCnwp8j8gewD79/KUTnJUx/xCTwc8TE1fbJ6/JV7r3OxC1vHFzHndxrqzSNUj2s4Nhr1W
BWTCck9buW7JpeIxkMPZ76XQKBeEWlSf16yQ0L3prKFjgR2nHjZqbaMJuUHDUcZ1j58IAKIS1Znl
qzfeU/4VJVyY3oStBwE6PzV27MmcDDTlCMy0abpD6JZ30FKm8jUpM+HxdOaxbg0Vmo5tONWAZ/C2
X+p2NcJcwptUkF271tPqQ7MvEl+yRHGWMWuZq8xY2evC8FmAcV7fyYC+uZ8CYiYaFXTqhdHPxGpk
+Ik0c+5NfbutDMfr8aA7gGU1bbkgMZmX1nzBIdIZMWpNzNEAqP3KFlQJBLJgq6gmwuFvJg5G+H9b
GBZHUYxPtvRcPXcN7CVy5qd8Sd9nV2i1le2lPDnIoab4k4tX4HyoMsZdkmrUCS/DAwehbWpXcm2m
zAPWjzpNrLGZW1Fs7XcsX4qj+YJMyy64uN3BUIvHiMESDeAduqwSxfJQa0kSOst3lBnpKL0Z9lH8
0GTYGULhwB1tqjN1O4Ks3vGpyFkiAy1r7/EMUXe8Guo3oLn2xgKHSrtot4VwhD7VxOXDJ7z3a0xB
sA9tOvKyNkxPL81mr9XnOIutzC0pcEiXEaQtZpuHUxwleu8YTjJrCCm2ukp3bll8d+y8D8QtR/9Q
0kBJYWGYwjAeti0+bjsxRc3TzNn07+ZOAXz7fBdoeSurF2VY+uRRWTvpn1SO3C0q2iKMzdXZHzoN
qsaZkYoM8yP4fP0Hsg13QmRZry5eN2lY2a4B5UnOUYZrzuieSb4zSQRI1FUgkScjZfyAwXX2KohF
o/3Eb6VHWbmzLI/NdSDV2fb9DlA5Gt4ilWW86Sn5emFqZ4m3CiSXmKFKQ7KBiVbKnBEDYCbA409O
DAJ4UP/kB7vGHSIf9h/PJgRe2ySt/vCTNy3T8oSOJmuXK8yY9j/aMl+uByS2S1LZ9y84IuDdzIoN
4hvSZODUf2PjHm/QfiM3xcaqDSTLEbDkzL12GDj7vrfAWB6Qe2P7+K1hoJgdbtipbQfubjnMyTuC
sP9MO8wkL0vrTxhp7RCdKVsYkJ1NVTobGUEXwgH4UK3S38stggMHzO27aj1Y7/xkvmfDD2uJa8wj
2pXWGS7W5n2BZOsHZ39ULSfVr2+sK1Pb3XLNTFt9KKB46W4zG1GidJWJn6VAQrEyPCf9HduY0mxL
CX/shqsoBXseH3SLlp2ScdQFGKxaRmnspYOLNqmJbcpdRIIl6dB+558xR6jaP8UUI2sO683U/kG8
gRq52gYMibTfsD8GHP0Z4E+gt98xel8VGnHCRlhKTiOqlREk4j1s4cZdcKgaUJJ64hC6SeyAxxF6
tXRMkKQK/E+Za2pzygq+DwJpxfUY5RFfmByAGcE2GxOD7e/qxMqcC9OFFi0JGYS90lLgCZMkTv5k
231MU1Gz5C9n2iCla92xkyc490dVTOpYhXHsRzt2t/RXBaYL+as3xFMBBy/ZCfhS2eyfhLfTczZa
dQM0dljhcI4NFOtx3A4n6E8mHwqyoqksczGw1Ptj8NZO0AP4SYVErkahrER+ysA+IlMlWq3VASkw
6svGz4I4oMJTeYYv/64awamcskUwCDJukb+OdoEbpUgIMPG3iSTdgPStK1RC6LYCP15iUHlqJn56
PepvTmdIDMj6ejsdy5QclkQYcCKyNmI0QbFETSXR6sTT+GJc1prNXFJKtQ6CAEnTbp/duAmbaTeM
T6F05FQztKHZDJfYE97LOzhCcVxhhvovgM2DfhwSgL3e7ynF1Fq8rJb4hzeT5p4B5hZgRGZbBXhR
SnQYXdd8r2TjxaXNsqKDFaBKKTuVbuV7hSb2snmcsi3Cq+foDhoh/aFxABkKh97CBPa2hdufKxrA
PjQAVUBQzl+HQpp7d+2rzwMd5nMooVKbD5qnZSMgOQ64iydIjbBNEMZSnqyiBjR0qt0k4KGJJqxe
wYUCTPYjrBsbKOQBb3mtj3YzBdTMkIWMSwItvhlIjDRRJ3Y8A4GUISoexNIXfhfO4+aUQoI8Yz59
MuITynLZK6K5Dqjqzx8Dm5UEzjzxnEjF9qvKa5ArwQ5VnkIgO/tATIgo4sH3g3yVN8bN6oGwVEMJ
FOJX/U25FBnUyUUYb3C0kccc1MoJmVXR+skZZpaYlgk4cgWwTPDJnaPQ+tdu7o13S+nrbzzCeXt/
qmSVl4Nfq4EuL3b5nSzt1w7LzZwZ8dY+7lrYqMSkCZvWHUjcOlEkC94qfVxL+BIwHtM7keIowUwX
FvckJeInofg/rJwnJGyWG75nyYozRs3sUkkGLyLYXrLRAZ6edb8sOVTZhRqqZVm6vM51W5HxVY0S
Y3xW/Us+r9jx3pKGhhdlWAEDnSJdjPenkqlLZ5ELGSePH+r0D5gkdkb049KMnrlVIICv1fADZAOx
xAw4PuDbdFGwhLcJ038kQ6Lyrmdaftkx6npDklUlBleMhMgN+gB9zYkg/mDqlrDaiEg1U8OFxUrA
L2iCuo2O1P3nKtQhNkxbFkRmI4W9KMOP4Die4Z5XBJgUq5rApOwUG57HH3469lAn70Fpr2F9kJOj
gmIQv/PHvDzRZq5dUvbdmQ4Yt6RYEvUqvXlYCzSr/OAItiLINw6Ry4e9IfGZipDMFw93JDMJC2E6
YFcNhYWDnkwoP6dmrle6pDI9/cj7SeN+YdFCUQjfn1HlWVTOMCXzL5BsaMsp4onOtz0X9453g83o
ljA8OWylcgPsxQa3DkMpceX0cgwnZXdFK4BSUpCooLrQ2h97uoG8CMPRJZI1ySxxtweuOUhN8jlQ
ZX7Zr+MeLBFePnhv9ud4sr2fhcjp9KxML9Ps6uIsV6mvRY0z8278CYQAdFW0GQ0e09RWfE9I8lAj
+/i+ooT1nuoXLXsgGDWX3EFV5vnEn0qV4fG0fNQQ25CQi8cpx7gvBbOtLb4QJ9Z+uMpArNh7M0nh
Fv7gzZhpgySPhpusLUqYh+MECynkvocH8+PsrWXdXnkAubG/a8dCEztaKwGumUF7ZZ8CupwKeklL
E5qcHiivsf4P1SSKjZb1DUkj0KNF2kLZklVpiFgDAxS4ff9fiHr2A3aZQMNe0VxGawU/CsZGKN9E
Ztdo43E7cdnfJ1MxeS+2CZ79/u+tqLxGdjM/6v48FEXbJpeq76enApXIZQ+7/1r8RVY6VMlLTPIy
un5Lweyk0Ew/n+6gsdjEWM2INXrsG5EHDTyRznOoM++sllF3vemPdtqXeeJ2N2umxZYsWWIe3nAe
MmJiKL78iiP90ySVQH8u/5/h44Yyy630cgS4vrlojYy8j9yHVHdALowyn2mq0Zy2EUrV4wfQXSrX
kOfooelVWTznll8gTTCFWjDqzs7OpCicr/OnkLR1TntKhXGurSmN2Ydha/UONF4dDeXlXatzNPR7
aw2rsDU96aNVD0OKZMK9ZXtV6xQoA57uN8TIuqfZeVR/5NwC8al5UTmxGKTAk7dAYnj5Z6Clwjno
XDtiuPpbDYnxIePi31xlQ9wa5i9SejF9dcAX9T372yemps49tvaanay9rMgJi9yvV0JU4Qn4Vy2J
/2A40FrOKLbhoFVuxWgB07zPG1uzaCiH6BGJLDI/MzuFnfUjuFVYnk5l9MGEF6Pgj2PQhcVBp8NM
bWUtQr1/K6bHR/ejWOz9HIPOAn9YjmIpcgBXTgx5rJFNSzilbWMgYKUNCmrVdzDJ2GmfByH0PONW
bJNyVwkqKHrUJLvx9thw4jOn78zxFJuU1OZc6r9UWXFHUT+pkNniAK7mNMQe1ciWL0ubhwh8D9oC
EmCuTR6w3U5GCXxEiqoq02Jd5VRM/qWKXTndTw46n3EbhzA5H5hv5YHgFgVt2tgOTfrhFi4hC1VF
jLKr/Uhm8IWObHSwI/AzuH7e59JS9h/dtOWlUBA2XiNetDV29e20lafkFAzYZRGqIppBhUWJDGlh
ZVOkoAK9gu9UYDiL9jhCTC4A/qtndoYO08XQ9ephIH+cnRmaMROthFEsm2bak7To94HIwFErovT+
AKw872ANrL2loNphk0a1P3S0ifsHoIChYz5U2yLhvVY8JyFZol6tQxo0aGIelSASVSHOwxDXSjUT
flVy0Dt+PTAuNB71Cfad1Qua6yQ6zJu8ZeZTcUyjnG+M/nXgf7ACrszhQwjALV4DXqbn5Jo7mBUK
WwPEUhQ5CeZuUCCazmh2l7T48uxHScXiJw4FtnKLC/SKEhVhArdiiacCfWabKKWaMnixWYH2SPOx
/3qiVdR0E1DO8oK96QQLqja2FMXNg/Mle5vbalRp6wLDRF3Opzkg0RCgCWy67NOOjNm3SbF6cBGi
rjlhXz/s8NZnjL1UZO081DYXrSWBmIdGW3uD2/oMmVgawyaHz5LAPnvX2VwwhjRbZuN27mLf9Jni
TWkhqKQHuhK9gORkALBPbGPp6+jaQMn5pezdmfcRjcrIZ1cf7XvLVZE7P7pXbNrVZtPiDwLkeP2D
8i/rlHgef0MixvKBf0IHwPrXV1gFv6/KmNKta6IJ2VqaqsTRtbXVkGzX5l5YDzyNkvNYchu5+PyQ
MVRjvgBJOe35GOwDoeRvDJXM91EImlj/J4yZan4X3PKq7HOsQIMMHn7aZB4ABITCU/tOVMRNeJAC
nsRJt+RhEQxyMGVXr2aWtPEk1wpjD/r+ZZbyotzGhP98ha6pHg0Wr14YuEtwwCrfeMqsBTtl+FSQ
MnxrnFSip1+8sGXqTX6sYqbj4edFT9r7/nTNkhQcfs1AoahbNEGUKeIsl+VLsih01kqa1+LVOsUW
sU0T/s3X2LoP6YtaIfaMTawq70YavQDc7Fv+4qHVArppkQrJ3SfeY6RRtIX5OLxH59Vr3zhx+U+6
KHPJ8376b8Uu7DHHE5lXGboyH9G+cY0UDgwd1uUVEAdRG1dDVONnsdBfWlh2S46MYZeQbkao2JhY
NwL2/OVM9j/YZoXf5QfU3Pf1JzJiSD6tsGndbBZIdxAQm6hIWVcK5QC0J0bh9jwgIiAgPMv2vUnz
Cu4HLths5jdJ5p3IUMhVK+OH5NLveRpWWXG1LLshe2s/4dhT8Ua/Gfqvt8SbVrU4+RN67kOTPc/5
+qIwXE3s1na8Tz8ZgY/RIkHMGqa+RoL4O104GPn7VNxZKXyPHy7ateAd6WV2RZdO2gZFkFB1D7lb
IvQFPq7UW2/DmitsbTN37GDHTWlVAJg3Xyk07WGhNF4v8gqffmBFfCI31i2+rNEkublZT4WGtxVZ
bhu2cWKs3sFDGeqf6JaBq7R/nx/OXQYZDlK75RE/ptHIPIVnPkVCTpPKVxwAH89NH1i/WQS7FjRm
3LelQkH1n4tA1v6whNGfNgeXHLDTUvQKS004vrkSmy3QAlItYQjOmOI5ZnC3XJY5ePuiRELjsXAc
2wpF/lrS1uctYfES5FPPOX91x6hI1EAu7JfhfPEp5lMC0lx3PT2lXfmw94SBW9+LBwDdWGmJ/vc2
gl6f0bM74tbWhAr5UC8UpgRHyrRee5/RUD3hnxqmLoBk4sqUhP3ktTEi+z6DvxMkRN9k39EnH+Z4
mHQGfIRmHslSC9RR6y1fh5LCyO3Hs+5T2WFh6BT5NOVxD7S2356x+Sk7SMdchpSj7jpZV2hs+WYA
A4M+lEZGuL6e1Bj5D5JXeE7HzOgXrBEvMC6to8EFzLRo6rU1MOwQMOxnbARxANZcWcnF0mtaGS1Z
UI5zlxDtcfHvKR3eJ6lWs6PWpYnwKdp+mmqJ59fWZkCdx0rMl/a2fuPQobWo6A9tY7cfUjR8H04b
HWLs4GQw/vn8zDqJJBt0vq0W/m9+8hYCyCUD5RjkquGqhnWuumxMIOBoRa+9c8680cn8ZKWMXoIf
8q6OG9aBbogfICQ+W+z/q8KH1n83iedNbQ0nTJL3V7rH9qwDG0Dp0SKKEH6rj6Ho+U8ushb/s+7E
hxzFKdP+2yzoYTpzZnu0jy4uVqgygJtLaoCspg0lfWTX/bBG01DrtsMjxo/v1qrlTEvL8LQu9zRP
ztyMDHsmcRJi8m8RFXwUf7mmpH86phQ2ts0nR7VwHqN4hDyRiwSENxshojCY1Ql4Kd9xVHJY6aol
osnI3258oqOjECx1t2yBWE31KpiNhXcjCKyacbK2ZIfpkKB8EN50ym4tlNso2lB6wMz4MfW1xjFQ
rXuHKM8UZiubeUOdAPhvoBSFSq172MzWzArGsZNfivUKqDw4pwRNdQm/knPSUyxLYaTzrxwhqEYQ
AG3ljP+pOecRF5ILNCGmRuUdXLO1itWTo/3DlKvpBVUJs4nFtdaKD73SnrTjq60WNC7tP0mZ79qz
Ut3iWhin4lxCo4QC9oaoUcP4eZxFK4bFkp3DyyNl3wfoRF+8BEXu5NnqJ9zhMrOyPtKVwS1ZR7Da
XeEAjf2kR6EaSedJyIlA5wyF4vM+Y3s/AcaYWS9xi7+QgV8jMavf7jv6RLfYfStgAFyByUC6ssG1
pEaDefr4AAJU8fywD5Ma6PJYSfLLImIRkisSWsoaFrSB0BkA1Ih54ePGBFDIDiEBxWz1RJyNQ5v1
u8KI5xO7iRWzuxoqN9Xgu9Zpxh6qYoEymndAu8fANOAE2nvabfsOQrWXL8V8TW2+lFBUxf1dhY7x
GnWUGItz6KCbxOaNBgCWooyk3yDg062XcSgMa5iA0oHyplebBgGMZGMyWyLxCEBC28ODweaHLVrs
+yL0kT2ztabGHAH8GJBwHJyft96Ru2Ut+vLWE/KQSz3bARUxI+wzyTTSef3c3JA+iZHWsuATsjOR
dB77e/ExkDFy/HBFlcsma6xJi4wyke65GS1iB/c9lP9NUninOaIiS3hnnvU5Jj/Hg/oq5pBZoVUZ
DyQ+l+dRS2CxEZT2uQvqL5KANEpBwT+E4tslKlguCsdzEjQL0GfYJI0LNyWW0YCBXp5JsHpiRv+U
GEKVU/lcuTINufFHER6nV92k8P19DCvZQCzUrKZQhtL0CLRnqxaKCH27U0x4rrob4igwQot96Apd
k/VCQCanbQV+OIYUXtn0aVKeYl+N8QgKGqMKfzlPSkqdEqcT+wkV9eu4Y/tkQdyKIlHvnNHMZcZa
qTF09WHOlY1JxE7fzWZpQ2ERSl/NyA/guHG2RV54SCXToQu08iU5hJz+3YxPyoVAbUicWLx0QQDE
UPI8SidXKqPan7iqrolvOxA8MBvSACvIJpC2c8QhaBQabLSzT79Hl+gc+JNAk1A3WZunVDGIgSdk
2Z2y4NRyJcVuBO3ouFmeNNSTquCe1SADIXSBsJZSCmv9nxbWUDN1fqZCdZBgXkjVVLz/ZNpNHsvG
mwiVG56Rw5hTtSIdr9q4lsLuX3dHWgmiVwW4a52PM5vGLLqPa0AS5vjhUb2Op0eqYOIVGir6bg3N
okPWFNFPhvPbWT/zv3AfD8T1n34/mqiMFDrOebxqPmzRM1IiGoj3/GYviVqa3W4OcbftfjD+DLS/
S97A5Pt8i3da2kfPNTt7dTvSxnR/f2e9y8qZBBOvXs2ePym2Aql1rgMnUxY8LSjJ2qoX1uoACdsD
fabLAUmbWeX48HJYjwvq7TBsdPCIn/lrAq0sxxKLhS5lsMAjkBIhjLtu+mBCm2EKaHuO6ecZBCqz
WqiqAArvgIWx+L+UiUZ5G5QZkT+YmLpNlK+ETJWpo8qkwdPYtuNi/lHPwc1sLyjzFN8AfbQh9Csf
ncBI4pVab25VzO9ASoeIaPMFU/x2IBvToG+ckPsHJ9pmqp/QLxej78rpOM53N2AofAVZwawgL8sg
uDqPgu41eL7a+27ozc3e6nZgLZDNiWfrtx/H6qVDrt1wTjGeboYhZqeNGILr1ZB8wtPMdg2YKthy
S1pLq0jTWR8iRjiYwsk2S0sR6denkXYfaF3UrvRo2kVrOIluZjfB2fTnxQBDATm2NXFho7hRkq3V
N71Vau4pFTZcnmVkc7iAMp5OpZ2a0ppC5S6HA7DBxLwttWhrmh25xWxgfthPB6o9jnmyOeFvM8KW
c1GYQ4xcdCqKi+Pqmc6auV3jDSTAFZEgWiXsKTjlWu0PeUjiuiyCPrXXazYa0TKei5Zz556x5PNl
zhBuIA8HyzcdmURhXEXBSz0AFeRqZi2+lu+4P6lVwE21GLNle/wewzUGZvtzQ+U33qVLrlyfuxwE
cedLX6zPZCGASheJzJOrqV1P3ya7h0q8AhVsZD4juL9aDqNO66C7RH4H8MtTE/dgtqeRdrERALWU
hBUOGjR6zLkZoe0wTtnPBTnQbEpAkAJmSTnkaWKuu+TQorfvECg3xQ+wthGXm1j51/9kaokDddRT
YF6rdXJkOtE0UMhUxvBQme8Ci7eQP9tuvxPNnUouUt3DM42oydokhDvB29ofIon9YcMdWsa66jo5
hAJQu9KXHpM/9IX1UKsk16aP9mLwOG0uO+Vm4tcQvfp14GD4D4bwBq2VR/pBJa2f08JGNiKXYMyc
BYxMy33HBZ2dymoxeYZ3HTUDeYVDHTWXYK0/I2MTfcSwhpr/+GGT7uwBLmbN5ZeJJJuKP7HXyvDV
hP+Q4l8f+3DmUpZlJlE08lWwIzxW7uK248aXUlZkhew8c+Z4Q0r+l51/gONzevqD16JbOEL/WVVL
gELyuXEY/gzoKHLmdoqvBwJFjyveYFFF+Uh7I83r7vfRlSAdvmnB2Dl4xxOjZzSNqop+Pr10voRC
2QTE+O3rhZ5arN5TC6UPCy0axakZxIqeOYLYp0dF0rGYY5EiR6c5eAX1HROcgrYW6BLNa32Ftml8
1MLMmrbsJn64sbfUiAw/Vq/7lNoQ8egHrJr0OTOrchD/VK7XVBZW5piLaws28nmzHPxOHKuzK6ap
R5dSCKqjpoHBjEKZnpTotbF9TuWdFZaEio23RmWH6Hvf+9c+l4PN8kN8lD+xoTjAuDu+XhrZGLxk
ai9ls9/pRv9H4bDY03Ey0izbGf6XT8GCLMhUtzDdG4janCKDTptlun/BP1irpfcpGb7U4YRR/W4X
0wkUedUHmEps/kXev9R0aNbSbavEcc8YQ9nXtEVx/y0rf4zko02UCHUYIHWNBep8CIQY8CE1F4VX
kPs+ogr11HLHpxH2LmxySpipv+bAhxHEAOjpXaY7X1om0puFOWY2Lmp+hqh5XdsBhQ9NUCI4od1I
YEpC+9YSX7Is8OVhXlPqrerE3PHJ7rD3MYu7wddc/l/dPt7ePDo56G8e1gDIFSzNh09VMQQQ4dAR
5hBO9U0evQD3SCsIXcabvaWu2sJdDjeFR1B74bHCoKjy0cQJes2fGWgSG1JPTb2G8AXE8aiFtDcl
rIGxHP6/w29HAo5pEF2R2pzXtYoibpfMTw3R5/yHc5tZQQUnuMk5I5uxOikl9wnAIV33MRjJP0dC
VSxLU+rY2rVcp7ikmpd+Qw+MjCD0A8Bu2DBKc4i3m+adTk6R+aTy2eLz/2GQGC5Ukkg33x33yeYQ
DUBwwJo48E5/gvKXxUWZj+X7+KnMbFW0snKaEwf9qxpzq+YxfITgWDQrjiraSmmuZivMbG29Pt/C
DZJA8EZ6ry36tHsdSqEQ5GocF9s2Np5gk37GEswEH6alDo/vqd7vE5jr4ZNu0/PI+HsZKe/ypgsm
4Le2FR009IRXaC6YHamE/TI/vn2bpwINx2Jx7kvNq0JOseBTtOzBTnhni0GwHdDHaWgFCX8XsWBS
Yfd3FTQK5lTqIKz3aMFpGDnwh0kUP+TjE70EQhwD3L4QpVd5iUIddbPKqlKVVO9+qaFsLyAv/Am3
ZglSlDi4znntB5U6e0o8jr2P0IzVDfypKVdQN3EC6v5/A5WN0fHPvbjYqOJM6DTQj0Zxv3oEVIaQ
l6UQ6X3cFZAy9J0GFRL7qsans7WsCQ/bdARLUlvDmoC1Sc9txYES93lNnzOFH7440a93dhMlEHqs
WjhlZIGCcUOYBG6OZkWRqFGRW26XFFxnB7MjJzIPRof1odyfqJyD8DFN7aO5Yod0T6mQfxYiC/ON
+AojE8YU+vO63SZYbXePtOgZctQgc/uqZ8nMt5XIhCd/eCyeN7fY+nirA41cuFzbFoT86zgM5u5F
EeN3v1tEeBLFCiD4oU2u1SdFSzEiCY/rLhAu0ysCarBt7qbUB+OPJPvlXLBdCp88EhmRXeVQ6X+k
oSdwaioWmWunK2mauRpOCRxw5svSEm7xplm0UX17lOUQwjhpCCNue0CuNjZYCW16Bj7TcJEpWEl5
Acfd7RPNHSqBd0H5cHwIzcgSKg0UAKYX4FWnf7Se8mf6QKQGwPDxhKMaDNRs3x3SSE4/6LgGr0xM
0XrU8nH2DznPi0GNnmPuTmA0kR1A7lGlZa9xUIz2AuXN/VHCiCaWMlW0tSGdb+FyDKNmR78Yvhed
W+KL1qWzPR+kXjbL2BDu4e08olEHtNhkTEGMPmDBNUtMfyi6FHe9blup4U0P4zOAS2sPHEb2rhro
Qxb1HfNoEr9Q1R1tUQEGrpTmYpZehsgIFmakgWDVl6noOwC7z5gNbPf3A4M4omHYOHUeaFb9dfsv
uW1ddgHIbFfIvtNSM6NzgdGCGEebmottEOLFXHCVAYGlFyM6iUavz1wFLk43sHgJTMcpuljwAnwV
0lo6FrNFhlhUXuUt0SnFTOi29oZWyVgEdNFZUC+0uHSam21oaQ7lfjH0gGVGHUrHTxFFW7XWQsBo
8vQBEXttWZQ+iZvGC1Qn36EnYTHuo5MTPtAUx8M8juqTMAHetnAn3O/vBNUNgR2GYgiTDnO/CXef
t9fosGMl82afXEjYnNHPXJSTIgNAtrPsdiA1om0CaOBG8KewqyLp4PQmqakWtiFoYjkIhgZJZFdP
btI51G++lW84Ogc4B/7Udsg6LeKUNMfKgXxevl4WGrtgqoe32Ct6Sy9zlDh8SisnIj2/+5eadUPi
gANt323L3Ji4CwIPtav32rzUK1K+sHi44iBDq1sxAHuqINbmMPnaQwfFMYm8h/+SJVejnIxHraOI
I387hHe/X5+u65Yg/esLO6hrmcE47K8fhr6WWh82r1E5Q3y7MsYauCF4YIFzXvebVx2git7Ib2HO
rwvfXITPFX6uWl/BZ9FaS0ffN/9am7uoOkaA8RXy4SsI1GESFbOPocSZ6B8oEVk54PeH27x2uUpA
V744YKm7MhVTGO3om8186+YLeK0/Mzk/V5RSFs2m6L7PiMl241oGb0aJgdeaEusErUwYD+fM3hUb
MNwLitrFTcP5UlU7c8O1AY5bNw1eYvJlmXnFmlCBdrp8ZpjObjD2sKLW22RQIMgp6WrAEbSyV570
Dz34AkQbN5KU8i53Xom/yHwWONvxOWkC/vNbeWAvbjrpj26PWUh+5GfcpbCN8wfZZxZEm6n8mdeV
5loBp+a4LLAsa4DlbQtknnaxaGHGqJGc+nOc64DL8Oy7KdKOPmx9F8WECXIjSEN6zjVNvYAFBIfh
G/FTd3Sef931jtU9B04f6RovQGIdzQytpFBbRyzK7pfSEnF78+K+WdM7Yn1Vi6ZYPMg8dR8LOGsC
DytvZrKIRoD7EOpHBre0ZqgojoB3wlqz0QikvRX3tx2KkCVLxbrz6GiCqZ1TgkPDTutc59QspMVU
5auji4f7fWgujlrXGp4Vi+q06oc6v1VeJglOGdpvM0xNJCm8y9yWOMrmBvUy3FHQ70iW/9XkRf5O
3gREyMvcROADFRlZKatU6nV+YzpXg8282WGBHPlt3AfTvCgF3cmZLtpZuL+6DdrDQ/x2RwC4RsZI
ql+orCOgR5tHONIE/wDF6FdItkrGnEk/fy9gmYB5mF+YkgTN/AebpuE50M6Nxcl4UmLj8xCatOSs
BrMm1RAnmKr+JdKL2E/e45xEgD7WXScZBDv4WuREVgSnVNZPnrq8bJ6Np8W0oI5UklPfa3D0Md3Q
gpGMH70wzYt+b35m+WcBBzCbWUcVPM5A/6E+gD3Np9Pk6hSG7AH+r7qKnYvpk2mVvV6lHcx79R9a
wKjPE6BqpR2op5M8K6cYha0r9/vRevV468HbuXlZ1YSCvArSI/FB008m8NEY6PFQA3hdB1lCWklm
EYfvdf/BpB7/ClawcWhh+clFCMvfjksp3yzke/mU1leV+XucHqccrP5qoSJvQPyBJZeNFFJzqQ8L
NhyMa1Qv1wwQGQYJC9VKePSvDTV6Y0qWp8Q9nacoV4vyUWrVrjZWSAmgBnYcmf8Ms0Ci0WcqtFFL
JNphhMhrCANyU1CdZZmow8tyvKHo7xe3skp8Vlhv9EHAlVXeiniSNbEXGEiDwO7ypqa64J8D8BF9
iIJ16qRUT4WfLwmmWtV6zgEw0DE5RtF8TttXH9HglyNqtvXR5Ruddrk7RBJ21VsaPNDBvooBp1St
mhzjXz0sAzm+SMhEqQ76obJ52DoMMg5UI1S2xmmrcqlCyVkwfc6kXt2rsXYI9zp0HZBPmLgZgAWy
e5PO888tTgnFFm0FHg0jk3wKqX65NNBwHXRB78qonSYvUD+RCBCR0orfc/Reij+99z9ue0L/HqeY
x47l6XHh2bnC5uRA9pHolB/Ni9gJYET9SoNfqfP1Nq7iEuQT9s9aEhiu3HnZxp9tOXhs9tKYOLsy
/mk0MOttkAPulBMJLAC4NDnyiA/RNCktbLqzrftICq/0IqM8PQiR3nmfaz4AxNJ8XdLypqij9+FF
DstL9B7jqYmQ94WAHex1XxOTQBivMWkyE3145q2KuWE8RssPSdKZYIgWfjydllNT0cB/+GrQCnGE
4/Z+AgEOnsmDM56Yy1LvqBMBiwkV27hYCA+Jt+TvlSy6miPBbjoDFqRsx2Zy7tC7ZoRTKbn+8h8H
h4XzXUsZ09SSBUey1Y9mixxHI2X9q1VMb/ePt7aaujQM/IVgjgYFpc5r1Mr47cNNruJdSapLxSn1
hoo6WZ79sJb1p+gl35VDItNztxHhAmlF3Py/eLzc5HUq2GUWFsG51++/PF30GmOH9Pk0ll1ha3uy
vVcdRIH7JX97CIid1WC3fao8v5IFuiyjHEmh3tMgiNMo96nvWLafbLHXyTkRwAGw+8s7u9l2Lpyv
3QVHtbqfixjTIwGrcVemsZ+pK6CHQLivyMUJYnXw7iOFiRFK0cCPq9JkG7IEuC2f97TG3r/xrWkE
KMn+mUFetHGl8nvIcZOhSSWaFRAm8B2H3iD8T16JdhmzS9FKwXN3blGLfdXNGPovWNfHkvKjmBuW
vWTv/dwms8XAu5LtvkYO1K5pe626arZGvM+NvUnkdfmdcvoD4ldnAGnXgdfl3sbaus/BV0sjP4EJ
+ycAoGUs6KyVU4uhx9gxWa/hJ/MaC5SE/TCAb16UsRYPGrMfiAo+7Vw/MvZPwapZPRoG4uhq5bVG
4F7yvzJEZt0HAU/PQ6AGK7AGYiFtctoTeNWid2dz0tfjfwrdeqaPpyRDTriTyKLATrcovenlUsFc
2fE27qiGCPuQI9PPBVkfBO9ezXcC69QJazINXujwogcy8yY7bV5eExAoHNH25olSAiwk2MbQP2cJ
uWgRsS/m5PbzoaE9fvrXcvyT267AVb/1Ny62Rr1r5DWpaWlaLjMV4DCHOYOOPdV5wx8nuIq3DykB
gi36gNfkDwAnCMna1603kQVgN3fbsFatam/zsEFLjqUwLbxY98WD2r5IaYpYdtT7noHvZdvEt4T5
R1ZcTDP9uTIcRzXc1A31r+3S0V7QKJC8aAGY2QDV+VkMNbHeW2yBpOLqk2cksx1QuiFPst8C5XWA
iGvOWTt1lHlSRrLGr3BYiInHT2lGuKPPFKTGARVNbgAyMCNoCEU54V3B9BndM9pL1RIsYjjj6t+8
2JUyfx+qvs4MsptNxRK8pdlehJI4IU+AOcX2woqK+UR7iYu38wF82uVk34vsEFseKmfxYn/d8Al+
GS+BJRG6LofVxd7ZSNQDJwNbGVuaJLOwxJBG8yXinI2mCPqFhDRWkqDOP9PxFcxrIMWCJnP3dWaw
PeLjpFv1/o1w18A1s6O07q1b1EnPbHk8qd44JyFkeKmF7HG3k/FWdcJoTf/mNH5iaZcNUJzHfvW9
CEUWo6DyZrdp8pG2Po4nmK890Tnw4Pa/IzZXJHQuOM2w7d/t6Mz20bo9xZH4XB53VXGru2aV8bs6
bKaPFLUk6haWOgxam1vDyEswuQRtXI6WRS9z03iGNeQV/8XrfcKx/fmoWUzPSEYV7Mzf2uJL0mZn
/F53rw5orEyyFNOCU9hpJ4bnXFbt7+/uJgvnPlWLFJ0KvuuAxIfsFBrCTpPsnBDbQEjwDB4JstTy
WxM2b3IyKWgGtGEsLqKeS+cOi4i/BjZggY7lxq9+4YA4JJv74WtcQd1dVJdNvqtjfirD+F8Hh98w
2+vMBoLRBeL0MICaeEIMnu/xKMZa4ZC+rOI0Y2hVVPaRLulG02Or1eg+OLuRW4gbjvmtMObp3KcP
HeJ9kmPqeUh/vjLeUXZJlQyaOCqM7Xb6DamekcR3PRHbFkEyeXdNY4mC0kckuk6hwVcwxIDUsVc6
PVBo2KdIsy6B7LP3fNECo9BKI5qzwE7I7WKvrLl4mfX6nq4/Wup+EEgLjIWlGulirJlFLXmYYM3w
eQoeZ8Qu3V+uJEVMEkPau+NAEXGyPbHhguEzRc4mGxI2HheJ4Be3APYcdLD1ZUmoalJG7Uw9P0X7
r8QOxswMJdsp0huDxPIPc5VBguDLEZRNa2ZbMM811QARz+0Qa/WYcZaMxMzjwir3LAbB2pyCjBfU
2DwnMxX+MwHQVAVlAddE+vLgk2FjCPewyGB67N6U1fBS0Fh6/ORVM5DEFxnQ6o0c82d+Rc+sZs3T
of7Omamt+bv9fGnwTxQIYkNTaddA08nxGRoAsx9IkySxfXckv08aMv7rRJPpIVNkPn1+AM7mNAHy
UHCHwWOAHGDOSPjy//RZ03ZU/htWEbKsYXQYLlf+TCaIUjJT8ruQ7CN1rdhazqCu9r+qAwt18B5P
Ehp8BhU3qQVIbtVt1tXCpF3m8WylsG/RkrWwpmCfUxpPnsU4t1qbabGbayGNNjyhDmZTLeFiHuEm
2c02SFCs4xv2Kc3HsDXafzpGV6y+xfjTBWW3AuN1l2ZqlRAPMkyM4iABDgRw/jIgRySQhYftVtcp
mkLzgixC/2l/7wJlDlAJ2MMJ5EJT3bjvoJCFJdXnork3CzQ2ZQ6kFbLR+yRp0f21oiBIR7mQ9TuH
y3zDsdJ8nzrUDaW71+naercUHfSpEe04kF9e6QQsOfpEvCZVZQ2G5NMp/KitpE03a20IsS5dfnDR
zjQwNBqOWLJ9tQXJ4x2sjNCn5L/gPZAv4Hvdo2xBe28TPDocQA4ey2LsiqgImPIOfk80CDHGitH7
xL6cwZutdCMAo8TuuUaBCrfh7WmdIHc2OnivcqN/mKaZWFbH+WMrYt5B6+6LPfv2GywgGKRNZBB5
h4DIVzmxV60DQlBs3gB40YxX8xYzg6RcJnmtykYqhO0w++8GY0ABwzjXWmQqfWQaAMFB03MN/5h3
Y0hryYx17sEp3qEfZHo7sfzdB7pP1Uulg2PbfTb3xsVNkLinSdFS2+FE6Pde9+zBLAPsDUKopNeT
p+NLIttupkrVU+6XTWcLHSP+exB06jYff3UmPuP7sLKtnkXAAxX9mhP+wKvE6InmUzVdO4TQcaks
MOiOQ6wSnyA++AxIaiYiUqYo/r52N8XaGyEqntMx9tbP37CV6X5zCZ5MQZ5EBbXKMrOgtlr2MQ9M
YNyggBaLYlp26PHGc+yjIWpEkbklHYgyb0togNOnlLKsZkt351egZna3N/9sec3UWYQYOVjTd2/a
0bWBXU2wqFy/r9OS2H2iWMHcmw0dSePqkoRJfeoaGNj6Lp4Jd62Fytbj+xpWxtfkLgzsKl8bI90+
RgTL5Nd9XVEFm7zkATZKa9E9S2d3ukcRAx4I00/J2HxRm14lH15fngp3FyuOJVcMrdHdxBFd/K51
NPW249y9yW5HgSSKDtG7Kgj4A2Glsb3WBkJbnrQPbY12yIlk3MRMVIpx30xXnxIKRQkP1laHsZ9S
iQr770Bsu8K12xlRKYCvnQTML1oXv7I5JM7VPvWKlsAwhaUJMtAeZ61wqRtx7w+vQhEWe1nmiUXI
HZEKa7Y/ddBS5uhYeUQ6gR0qBAN+lA+3IprPxwnn4J7al3Rxpmkyeajyoeq4OngAtLM6n3gYbo4b
F4D4gh/is+VZMWUpN6kpqZkOGxSxOf//odkgiYf2yksvwNhO9pafA11ATewKhNGatsAmjfpDP+RF
H8R3j8MlT/Jh9xTPGBHj837V1GYz7nBk7DpHTwi+MOHTl/jyKbDClO+LzhsRWMoSCVmbJWBcMn/B
F5GdgC7kQhrZZvsOz4B7X2yN1CHgjAQw5vAGvbxTk5/jU+Ujaq0+Vxc9zTEPKjaiMAMBYwMv0AQi
qVmAgrZWmDvrUR9dRwFMmkOvj6YEGT1AJalFuV/tQ8AyGwChetoTu9zkE6Fv9z+eG2Jj3yd6a7k/
TElX/T+d8gNwdWUJzfjeBSkIanLKdhi/E5hwB7jQBghq4xV4bYbqeTIZ9F0zXZkftC/ZhbG5TNy2
Z8Xt4kkswQ0gTuJCyR0KTrd9QI82XqV90hTeGPtBeIRnIAB1spY29zW7nhk7muIG/krA4DlCAmiE
2OvFDyJslZ+YALXA/JLpB+R+n6ucj42uALtbTsBN+xuLHfd19JSnzkuuW4MS8RY4LnIYmG8uQ0mF
4lcK50txWnx9de+oqha259r58GVM6nNACdzHJU+JVAHkoQkPg81xesg79KUhY26C3ik1sCl3Xu0Q
j75yPOrO1CtTOS1GDzCbTBulYDf+3u0dL74YcUJexIvwfjM8tOC08n/qWPchP3ZGi/xLdj82wy3J
uFLsyOBhfBOE2R5BcvYXHmmx9g4KStKvyH/NSxffByhFsrvoIVcATz2rbInl0/osWmZ5/yljR9TR
7NWy5sXWw/2R+OEZ1EwVOIbsJVqwBJQQaYHNUFD5ukZSPEznbjhFA8hSHuyUeNkDTtGWVu/YDkZT
oWnATYV5fmoTHRum7R/3yxXqbTmqe/5d2L6z8R+SlCfMxOEMYD9/8XAcvYhl6paWdWpAfBLHKZSU
/iYPWVLBI/kXtVZHeyFoYg+I4KpPTNG8VF8bswPj0quq7TcBDH18p/FHVKCmDMcMAtMu4Ubmq08k
B8IjNO7XdaZL3HmkzKRkP2BjwqCGZHMlPZOgGoRa5pWnrnE7muqwewx+SYm0QhwK9Xcr0dLMGxeV
hfLgKMdY5X1JbFxMwuh4si/mjISd5QJu02ypL4q6K/xNivNbJBlFm7d2HozfFzOZvAic5n5yiwv+
myeHePUB4g8r3g0TsSHixb3tTTJgqayGewP2w18L2pbyQFahDwLTJaxPj2qHsDm5WNegXDMhkXX1
Xt8TJwKERu46OJHk0KoQag8fDPqQp4OoS/MvPRivR+mJycOTbGNwOIkqpQmZBUQ4ENgP1pSaNnmu
LakK4uNSW07A9ek2Sl667CnrVoeu230UaIiFeAATgXM9LcRJTWP1Sky9tjXojEAYreEvjm6ND6wG
eKXZHVCt2kUp/4oF6HzahCpcqmmcJeh9Ca1jET1NfAo0CP6SorQuuP5yV4U8I1PdJLvKsgmHQkDa
zbcwCUmkHD1WgskBkO1akYz4jVnXNZ42S51auselmseW1PH3yvGwSdscvTc4KZ71cxx9YVDYVqt5
56cxY3luR9HzoHpyTCGLqmE7i9KZ4Azy/ig4ZyKlTOw5kifIL3TjK/lnTJ87X8lUsucdy6MrR7JJ
D3rjkGX09Sr/mGORP1qmCG1SQayBk85H+423RXuqb5JeIhtzObKmBid+B4yE/dTGcMRaBWjviZAG
uybyQpiFdKXA9LqriAzV4blT2OLrFlJFIx+bj8yzU08gI590/Adld2cSN+0e5s1Hpi6Fy6oSpg7p
3ckHRCg/O7dzxoYFxrMxGavatXaNuOx9kPexVjYMK0OmyKjXRdv+AtfECAdT+251uAqtknDJv9eZ
M5pVnPCNeO1T3RTRHGp9pIj/oCWVJJtgJYyRTkDef5uGtf3d68UbNhJnv1aEEhDdktPeNxHZKVPp
SN5bLA4tn46jeG0wvKgjAHalDXFwTw+IwfDiiuHavmFcsM2a0VgoL2h4OiId6tWGEz2oRpAxo3QG
TjwJ9xfnL94ThIXq5yvkPeG5S6rFwrctfD8yAcxtDp7cCJVK0mOoQlR5cDRODTXoRKczEgSEP1kW
7f6XAoa0bqIj1KJy7WMImAbPyatXuRT9DuWbRN0MG1qxc7ufC8Db7bDuZhUTWCoiqjlGoHpQ84gM
+wF7gQp90UjJgOBB9369ofZnzh0+8//SzAAY2Z1M6Pl0FJytvMi80WnEMRBCKlUtNtA6GgRHO3Yx
8Bg8v8WjLSP2fB98XRUdN+ayCWWwmsN6exx+I8ElyCm5RZ3lgNfRQN2eYkRg9KFUcn0+W/N2kjqV
JrPoSeK4AsNbWTDG0kdbabfzlhS14ZUxiMXul3O41+j9L5Vp/aK9ABUbCRCFWDbb9mRZ78avBmSz
hE0VVHThdfwZsmN3LLtFzp34lIziR3SQURqU6VTrrxhrmXhcOHlQJMBfMnf42IOxdZMeADSgbKXd
D2A6vuvCr5aZkFnlqC8QckcXJbDLCxDLuoC6nGSiEyG8WOfWAoNHwnWpC0jgvN+ssKWwMoYcDG0M
kfNWJ8P4f0F52Bw5DdPdgQ1r29F+gwbX+2rXDayi78fC2xFc5SsCeRULzGGvu9ay7plaYJMWcmxz
3rC6/NZX/lZAAl4ADPVnApC9nLNPjSoDcx4WnFncc3XGYcdn0OFrAVICt7tBqjKlTy+gceT11z5b
s+D7/LdzKQE/ZZ8fo25bk36Bg3t11tugx2qV7TP5WrVq3TGQCloSnMYNsuLfLDjpjXCs7Rc27+cS
0ESO/2kbTa2oJU/VrChIpJ4N4fmwVbECaCe8uj5HwfzZuezl+NnVI5L+r0PtvVbBWtL0bHYGwscl
KzpSUde0WGqnLl0JG1MPIhRs75emviIX1ywp0tPo6PMCGrdKZbFfeuLLFmYELec8/cNTGKGodOcL
A2Zb9fyNUZyV9/uNtKb/XekpbLHTFHeqUPPDK9Y+/UbCMucMKV6SJjzOGZ2eWZyz3sUCfIIkJFkI
PoAn8McbCfW4LhVQ0y+bd8T/7DRosrtsPF+RKCijh0HTney242de+hfLXLHRsW8865cs98MuEIUa
MuiCS39oWTncKo53IH50dYNTX8UA/ZetFyj58VtnhbRVAKUSAloRVcqgUIkel+IEyoxJnnDfbEfy
0e+H9l42qZ8pRr4SKZrJxIbc7s13+EiognM7nC1XACKN6LJsKBhIn44S08mdtAg08r1ljGhGmoha
iGJFfxUvtKJMOnjAzl/hwmr5qsbnJ3EDovIV6F6iffOGrXAChIy7xOFZ4QtjZZJyo2+Kvyjw1TEu
UnyuUSv+J53BsdGGSiVXHPxp7YQkHCaLC93molSLuhOgSvvyoyaOn9UezfthauVmxywxYDukM8oi
fCCyyM9O+17v8RQ+S0sVJgRYM5cBcRzk8NEeRBp09H+RZHbuAL7tytfqu3luCtiD/ezVyyeOYXaz
Ogcd+PTEi2uB/mxiDa0jJGS1hB8fs3kE3H3LOWlh+rAugJ4Fi5ewZTwaYwxvywy6xBRS0RObJhAl
6E1udsaDTUh/HRtk2cuc2/fqf+sdP45SjFk/qbMdV3Z1IfW066hE7YJ4i1uCtkAD+Zf1GbTI6eOE
1LtTWyhEVwOIKsnT97VR7Op14ffkeiAfoERAHa1zXQjoP+PwpLH5s2UUZl8OeDTAXpwV62NmwlzH
550EHLndmoqAAtXVHxOaH0YpGvXuGdYc08QAMo9F/um9s7KORuhgUg5eCNGeQaJgw2OreHUodmRh
9jx/2CVIds99qy09aFSk3VpRLZ95twDJGmObcmrrO0L7YHEeRsz0f/52H4CO8du/n1Uf6i/44ASu
FSrdhTjjxtxdPP+DUsJsJ2RJBIAz35EcutUtfPfyY4ZZaQMX6T9MXQ15sirWiQS0XQMuI7okcrl+
bRTkRfN9VIKDeadaA2nTxXOsYNFDS0bCcWzWxnMoeoNsqUvxfeIAIC85myENnAR15Z+2VOW/tC7r
Y0BNyW9aYvyysdx4Gk2wAwgjDhIW40N6dM9Ebr7xadKcXWV2pkYnjZHPHiythlxX35/P3iV16AdA
nfsixwuNDEZU4KBIgai3XD8k/1Eb+4C71e0uBCxJ9DDKINNiMqJnPyTDhlpHWru9a816jqtyujIX
CyXt6Smc0QtKxibR/7RQregHCMtW8XX4Vcn8ge2m0I8gHK5U94ml2RQ7mRuEufQlNbQ2aELPHmq6
LMALoL+KLX39RC1fZ1ICKKTUtjRwxeldzfWJrRrPxJkWS2qsARqgxImVSHJl87xm/lRje9dAw4Xc
hL5EWSwY/AjGdZ1GCv0pKSSgjw0W18v+5qIZMVGVL2YaQ09IEKjPdDiyP0IzxZOu/SLSvZw5x/iA
Iu3l1w2FgNJe020h4goJjo0eNziSHm6xHvHZOPYoDWnIZUOcowpuGHWwcDGl+LhN9m2pZiEPU0Wq
MOT2nPhgIkkwvrtF42fQYozqjZ81P1R78Agfw6R7o6CCGpRa8l5Bp+SDtk9L9aPijX5eA6GX68Sz
iVPDGlAin1SfN3vqbrauIys1zV1w+6mI2aGW2nzSl8KlDRBjiDLq37hUgyQ3u2ynZpNGV1DvcdeZ
uiF61q1iOx4BTTvxz6Jpm4j/zfPdWrL+3vX0QaUsqYPU5GEj2Zu+vgpUIPUUof4PA51hDuKZ8VmV
5DorZbGy3Ep4XJjA+GwuL21oWdw4HboDzF0PpdvEx3hvc7FxtlN7XLMC7uHg20YTbfvbddge1XcC
aXN68KJWuizqDlpabr7QO9SHuZqCAvNndsj4Z61DRndpY5VnV9pQOZiz8z1YRB8rametH+zwsvWq
8FC60J5X8xcpJGYSpHUSHxC/wy667EJ6qu4+zOJRxaExJFH6gKRFVMK8UFiXWVvigyYS9S0ANkbx
QF4r/FlKXjCTqp4aUJDXwYomPUrkbFJRarKLg8GWvXsd64ozPtCbkxoM79mQa+qSh5HUj0xbtxgD
AvzTly7DJJxe+X9CqKtiQcs6eIikFYxxcVZmXslpebgPbjg+KZv/GjGvUB/tKe5rRrSzjbA8pTXc
frRcsGYc5GYcxmgSz1mz53QMcUE/ij/cj62C2pVOrNuzp+PKyUk4L38ELcOmFCLPUWYRpRwPwS2K
xLN37hGD4iAETC0j2VYwi/LVXpF6E7eOxSTiU2xb4PZXnP5rV1iKcsRo5NM+jI0Eqmx83CsEdCqA
c5NqQ1FjkcOVvlIA1v9zIxnVGdaLflE7mbCShflnuLj8CEeYGtWms1ozFXGLlnsg2rXGGkkbidaR
hmlNNSlf6LLRPRWBtP4lLTybpixiXgAErluFDlUmEnWN0UAb56SRfmUhxol9K3RHNtx4eXPT6Qpv
wivEj34uOSJzU63PR+m67GELkPO2+ReMoGc9gQx6yGK+IczUVNlQ/J3tSi1Irs7AYDHt5rWFgByp
v0L5vAoaNhgB5pN3jPWk1fJM0KufFmxzEicvG6XPkr292lEmeq+QWGmSsNqVBeiANGYeT7VJdo+N
tIRNfPypNEjM+9tTdCC9cZetNUVAcMEYkoazWgkoaXHtXkaghgL8GG+DUE/hnzw8iiF/aTnuKq6U
6QdPc/uiqYvvUQ2dikLitxpdd+pVKkIEUf2R5GX5VS3J1TH3VcP9thAvEv8RMbzBX/NVlWk8V/F5
gfP3FhR1Ynn0DTX2N+LXp18ORmHLhECJX5NgPqGqVLbL7l2WD+aKk/NnLVPRGSTnVj2xRwJ5U7wH
eBuv7jZDNv3at6lOrY/RBTFQreasCpUl8+llEpq0hV3jjBhAxdhioKGsLHtqyrP08itYq/96Ygw9
3QiDYEUXSWOBCvaS5cGicBddjQMaKUFKTGF/4e5IUI61PEehm32M7rKVvJlyAIgI9R6VTbUws3aF
sVSdYtvFO3WzIulNkV0ryXTXxoAVCfnFQo5U13mLgPV+bEadL3qvgZ3bs66WEbFODevPvST95/Ce
J+dFuhYEU0F+VRp9Z123EJxPsCnqNWy/w69HLvBFToEdHkxiy/qupgAKX0PYlYBE3LwzwppJs3cq
sEQ9ta1EJ6QiAcc5I9M64Q7b3wP7dBrEvJsw2ZHMCjh4Z/LLOdom0YactFi7qCxJCzNIB/+/nmFg
pqX8Q7bdShnNOJhZZOXD08JQscTtGboyzSWlUk5P+zoN2D/ceMyS3CKAGrUH3LZY/VCWo7FTcoLO
S28RoICrnfYruGlYeLpoo5XLVsrXEnzVqprL0+stve/wPNZRQNpWzGUyXgIo8acSYudl7/FQdV4+
/kXlzZrYzzqt6i5O89HL5Nk9uydSFlbhx1nPdeMMPaRW0nyzs0Djq8j0a6+XcuIx8LB6YJUdtufW
ibCvfgygoweK0OtpSJpaFtNfpDQo7XwQV21d2HcGVcRYxTqwbikXw/cYntPKUH/8/LeMfg8p9y58
/YdnD8zO5U8nOa+WD4tVLzPiTpukp+UgwjP+It43WMaMimphPkvWO2fjzdTLzXcddO2sO/9x6kBs
Xgi02+mQVF9ADtLt9yca07ProZtBgt20o5e8dXUw7Yfa5WgI7GYvWyHvr3/LZJfUhedXZmbaXjxX
lZKPIrADClz9c7z6ys5Igz2U+z7ANyZi6ehrY3ImfkSAPqSREdT2iHMpLYAXrlkbSZ5hrW7oixm1
IGpXfxu190U7FY5bzCkBEwj1LcnuEJGfgMGpcl19/kY1Kc+UXR6BcXaP202bDCtdViJCtH5b3oTZ
RN7amOlG1ddXTGbVeeP3OPWd27MN4vL2drz6bsvu1V6IHVmS5zPjoCBOUXHf4i/+aQt88iSTHXcb
T7dFGyHA6Qs0wu0lAmFaSxIdM/KbMz40eyPQy1+HobpUI7lcVDwhfR0KiBMI22X9lKa8gyLtyG+/
Z/sxZKYynn+jZt5a8zWG1PW5pboCVYkaZ9ZuV7OFePXSgzX66d3vzB3IEfUs91lfg7Hnvf0/Moq6
rVgVrrvd5KdWgEOVvmSHL4Ka4XP1vf+khUh2Fm6qruFWgK1ZwhcbY8/hCHKdZtLNWAMguOuC+wMA
rhsl0P0l9CvK+/a+5k97m/yFozNe05xKAEKRTb/38LwCG452SfxVsW/twAUW7hnbE+kLWRHv5SgJ
2pBVuJeA2CAG5Q6FY/pVjCIoZQiJvQGPaDAc3kHl5fw/otcYJnB2ZTn9B5Fl3S+Pl9naZnb1kxcS
N3O81kzgJPH3e2Th4GdkWoT8Sek1tZ1HWfq+hQ5g30e67qi+tiJCCpAvB84YgiwLlhEV2NhEnOah
UdAG1bd8RFVAX/C4IpJmjtYiXO3vVRJKhjLQ7qNAFAic0M23pSrwveY1jVuieVpX2wCoyIcHAL//
zinolBk+a23ZCctjgDjVs3VHCZYWjkxt27rNiAUGRnVJtekqyQybNyU06pODY2kdmdWa0Pr33qiL
OUC3xLQyo8GetlmoGHjJNGu+QJT0Dc3kRvf4DMob5Zk9+d+KNYd4knUmMOd1HtQKwL8J2hJabx11
N1rXrwEESVdHJ50kcRvG4pnpHpwhipkREeOCKCwyYdQ61Qh0Fc0++YkY0XP2YN7tLva6w/9sl4ak
8kx7TobQDXdL1GxT2EI824fLbA29apAElFVB7jTTWEZnqiGmUeUL11V0GVUE6M9JrqYVQjveNOrV
WAs0Cw8MCuFoeJ6iRNl9dTX+yjleaOz7dd5BDjCHnzcVXIx6u/avbvGokwt+AZzxqT4Ha59mXOFw
veaQTMN1crb2xImjnF5joNIe37AfrV33Jc4i5meARlG/lcYGkfy7ERKt9H8zt9Lqdf04vma5mg0b
2GqiKrjIlSlNXylWYPfq/mvMdLMjbYsgMLzgnPE8dz7lzpzRfleUdxnDmaL3HD97WedMLiFoF+0u
iVBfKHzPxQNye05Wo96+N3s8IQ1dL2P0ERo45u/j87TIH6PMQ58waLq7QhUwZBstV7gJcZJpQbJV
fqL4Ne22Pde194Ra+B/ke35N3HiKK3p/a7vQOcT4punm3mddpSQu9WXKKauwbm8TyKHtu5gjkwus
o9vCpRs/qPFW/P4b7qV8wFdTmjyjwTV1GeuS6W07hkqzWQTvbnFo8Wzz2Ln/0JS3VGtJWOk8Xd9y
vkK6DkHwGiV+LR0HRWnX+gPqL9ndHkjoj4vsDm8Aku/kCGTsIKWo7UbPSb0SGQMk8AhIHo9yPwdZ
leMo819iiM0iKtwWtTq/qJbQfWRUhGGc61C9qIVoayNX5aVn3d8R3rZ8Qa+I57t6QRep/wQw3yji
8aibpw0360wbzFmzyotL3B8mApt+JlEc9XlaZtzf9WyiSVJpspeDF0XdJdc/zXcO7UwClW7XXf+C
vNryYTUv3TfB+QegC0JOOjC/CBKNxe3r2E/JSi/FTT2XNEm0Xay5f3CP6fuX0bRKJ9++ckxflRLa
sNprHJTXU8FHsHQt7Mx/UNpai9Zl7T+vKT2rj7Ub4+PmrUkS/eQxqbZg/YrrBc5QGAv9UvCwi718
MSNm9TQofbFImXlXg1jmf1if2lMiv4rzfJ30NqubB6B31zg4uzPCDQkTuc0JpFa5fyhl1OmoftyP
4uAKiNYWqFqGouSGBKv+/+WIyQhkMg34162Vq2WUapmiJln2Ug/DvqRQ+bpavaVyp3rKsArloVDk
1ucHe6ZM+NmKcdhLqI2Ms7Xs9gHqBGQI3hUYLV+pLtkDfLdhp+cLOytqE+Xbnx0khTjJa529N86i
rfNqEdDmKbidXB1GIFTRUfipNMLEx7JoYaKTEOcZnHS6mzFwoVWdCzF/OUijgW+f52xE22waIDTD
o1FNhhlfdwQ4rlch6A6AVt7sgU066q78bSPekcEbxrMYf762RSng/dxY1eDFatvdm7hJniRwjInr
oYf6F4Koce+mPyyCRjrHI6ARFjMUzK8M8/77Nx62vYS22b9Kb+8S86AF/GRPn0Lzpe6HBXNzPDYS
uxmuoVOhnXoNI2oEFwxXZ3lvIpfUhVljxduBMJp/uTT8q2MwY0iDnYCGTpi0+EiSLKXzkl8r7210
up7SsD27MJUuTpQ63sV2en3NXCy+0Scpyg9APmcgRrI8LM9SvSgmJcxKzu466GkJwFDL8xpOxSqW
YXoJTJBAsfWuLTku6osiqHiM8/UEjvDjW0FBFRFU2hE4wA8NQ2KSNzQmvBTOR1mXrQJD3HPt/pwq
xEqjiQNffiRXp4eF3CvToxIMeInTaLExrrLCVNntSP0nL//RdP9ZNcCZngcfluUsv//BjkojcOQ0
vrlX83hnz+Zpbuh2dsRkU4gHIWjk3bJqY21snEi/X3TpXzWXwUMi6EnpwrYT43watL40D84uz1J3
zavC0Bd2xO4NfSu/JOtSaPdyM/6CQDC39BKPSu5j7NnPnHLNNk105um6n3l7OJM6XcpUFn7YbOrZ
C9UtA0MkagOJ79e4FAcXTOh/jkn9e6gYnMhC/HfApBgDA8V73thcw/88o3D6sKqIX3POC2LFrLxm
SbYlzZiYbTtjU61zSkQPn/IgZpTNhUOv2PpcbCUtLq3LJ2iWJk24CUF0OQp8QULWBztr0aXDneF/
1IrJgpaqwlmZhyMB72tX2POKCB9TC4tje0D3nB/KgKVOxQwtuAkK6HG8vYganxZMWwc2xwNAQ1J+
OS8Rs1FYooVTkq2w4pKYGNCtX4GvcLEQ67nm1SOFmtJNvmAAXjNZKrKzahCW0YUPu5inSrE11spW
iNd9tHHW7DOjiQ646RkCvPXNnvklTRplYkOwTyaYPgW/vVl6ksYUoAln7F6r8rYXT2kjI63cgWON
2Xf2HgC9QR64ldmjj6IHxIlueRUwDolfc3zxqU2UnubOFEQepiBkumi29M+XD+Y6Fr5lqKbnqr2G
SEFsoeyb3v8xdud9kFf87g4KqW9EntLn8VunjVBnGFtMm+ETGE2XcsGjb6zPj3CC3dn8+uZJxWuH
4dxRYZ4yCCdMyd04TRfjeug8dMfkYRZLonNV2Sdl+3nEg9QiJJekixoaR4oJKbx6NLGJlrR/7MVW
Ez7lLX31ZN8lJBH9PKQ58LFwJ+6b3k2d3PL6cIn9VxWFqF79PUaT03Jftx1t6+1+WxJU9jHRSQgY
GCaVv+ikiGCAG4aF2R9sJ+oAY14YfN/eLs3cpB74cCIjONAqbVExaFv92kFUvMomDBhNn1zq9f7d
4dKEEUz9WNDm8ESfLaqmQF16uzGNISKM626tq6HR9cKzcSF5fLvTLFjMZAmFMGxoKrEIOV8V7F1w
PWqNmEiC2Z4i+kuhbH23bonHGaiF/TEg+vh9Q2UhMiBMCp44JlNS4zQbqUmavxNXT9OnPRh4KE6d
qrqPxoziiGmJT72SKdGRilq6RQ+umcjkiDLWDG+XI64tvxpPzxB4Iu1Bkcy8gELxlav5HFRs9t+9
gS6WrxjtkS9iRaCP1BDrnZPpU1voAnD/FKEErNZuiA3EOA208Iz7Xq6op9ThacMgjWGgel1mo6tW
lUc6JfcH0nnfIAlYFnIwR4+nnkGCho9BUV9C8rOU1lT36ZHOZcplQgH9Fa1IYtkoTwe02+J08AiH
17bCneyK5enYXD0RlhysLAAy+6t17o7B4yDlv51UO8jPeTAOvG9xEqatDoYfDUHO77oVCntPfY3y
hO37PQ8PA7dzTG6lt3FGDbtyhKOCoi4CxS+jjyCpCnEKQUjCDL0C5X0j94MimGt7HorkZikhT69Q
sKX0lieB5ba6InIOe9FvNaqKAXvKGYGJZxWUVrm0y+7dSgJAAszNAj/+22ddkaXnSiLvjJZ8H62m
EiTYZjRl8cgiqOEZ88TaVExiL7IJ25T6yoZ6zTAoaVFPiBCwmbMudrkiYMejdmXyr2ZwVm4NDCxi
Hc0U43O7rciNK0WB4acpnM3NXf/xJbazDQnidlrOay3I/ewx2TnceaLZB3cTNXWFbZrLbMgOzadR
fGUcRwZzl3swIDbdSK0pqiROMclEEUa0iO0nD+Ya/RJVONa9G2dsMFwBjl5n/1YT4vRcCo5ODtqM
UWwJRSSackgu4pk1TsWE9pxRp8jcVsQ0eIpPoPAfcLz8Na2Q/XRMIi4+Jhq33Lqeir84+kgAc20l
Y3Aof70QLSzzcEkfIeSFwYP7xL1p89QncdCBCXyJWbs9t2cvFg45VIOtD1FMj/qHzIDcfTx6uCBw
qJBT7PXXGFGmeXTYC4TLpDdAjTsI8bULhBa2NkK4BJ6GEiqDxmKfk680tXuphs4G6oe+zpXXYBOX
GHOZhEKp4mWTWIU050HrDnMQMcjIMho6QxOS3mpolxa8yKXDmEKxp1LccE7l9VW6LOFBD7HgvUdn
CFjwpSxb14GmQZOVoNEvBqxbiVXGD8hg1IbI/bjNxaVvCmvbx7whKpG9M9BWSxJaW+jmbTEMaVkS
QzyijMv0QimeuyarJ5uqjPASwsUtVyl6OYOhXzfTQW55Biu0T49WMcOkMjF2bbGv63gOYLDmMbPs
72vlPnVPEZXw3NlaMhALGnItwIwVNaPakcS5+QEGM3TEN/6TrkscHgzL5XDuIGmBB40P1Lpqe/hq
UHTVpoAGVX76BsX5Z6Wuer9zq1wE/oPCrAO11fJ7+4yzF1Vx+HOUSjScw/zTUQT2jUKb2IMrJWOC
rCsMQd64WC3xAIyVUq5MCGiVLmtL33HhQO506SCU8fm5R4g+faDsieIOLcamWh+Fd1nbYfDrmSjm
W/ptbh27aXuswN7X0QCYCcJrAUG8+eySYbBjYsj0JFy67yUndCQyjEWU1ge8cyH6FKXW4Dhr8tJf
uqAd80RwAMz//JBVvpHO6Md9pZp/3OkIlNq4iyiAV/nc4CzcUUSVArYr90Ti6pen3PhcKzzEwmKC
FATC7GW2nUlYXlPKeJjSVmWz1xsGvkp8IOTz72hn8ztCaX360zMYAnb1ozUmhaVR75LdpUVFrXKo
hzoiiKxl751OiH+V+cbluffbq+LXwCHTZ2QlNfHfEDO9mVNlpVho7UhMmFQR3IFos810VrqmFqK6
H6QFgustx7ZJj1EYpLXga8HYhAJZ9JWx0o7oYHW1P8oqGZG0QzQEWJ0lr3SsJjbuS3CnmNiQBA3e
LVZ6OYOIx72woEt+ecWIZqrdUqLkMbaQE87JzdXYnf4+GwVOFriFwOSz6Psxm1R4Zm5JMHm3F4hP
L56N0y4a4VzFMKdGzM5gyzp3YeRMCa2ssPkuPU5Ej8yLB9ambpgk9IVIPa8lCfJnwzE0T5wB1we/
MduBH6/H01BmRjEhUSCzW5BTSSSfvpnSlhG5HdclE0o7N/WL65wNyhlhbdfRsKJqdpMQC4dbVCl0
0lD8by8CEHFepmy453KMWqTHmYJ6KrpABN6dGv/0qO0XcJQc/bVw8h+h1ZcQBg6pwO231xOTlA3b
rtfs4V8IfrrQYOPMT824gi32Z7NFzg9U9MJdgnJ5DmUg4xDuuG1QbUz0RMg+6DT0r4WuPOchde65
wjhWv0QQwJOyd9XSRWmCYdIPFzT1RzplNN/vpmvqdLwR04CR12ujG9ykXvfu1ZwQYZ9VoDz436QZ
A/QXFJM245aw0edNJUE/fi4/nJgPbGn2KU79h4t8pZzht4qMGOu4y4kRx2G0j2sanPxOcstM1Mj6
piE3CZ9j25ly6WQPTW6uQRyXPIAEFMLxftZ/IYcABd0EcYKgLGzHKdisYvwyrlU6Vby0c5Ti/RNI
I1QyHy39oucbBAuJOjqEcGgbBA0Bj1r/BwYMUFbsWMuloa1Y9gPAhMg9zpxT8Pn06rS1K+rBCH0w
ekLg4wWZVSypE0429eGDLdYa74w30UeJ++NVB5n2MyUjtPkDX681I+4F4p2Tg7qC0fapeYUlgktJ
tT19kCF+g3d+EFZsfA0Z0jKEkNBKFyLVeyl3DrHtaHOMxMWypDx4OhVYVhgOwSWDa5HapjBtTqvX
/EZY+YlAci8OAz4E1iPGJGiv323+v2EdLjvcBxV0/JLB68P6cxrKLdD2K7snHwqZetdY2OWScasu
dImfX/OjcB13HU0m2SK561b4HUI8OrkrbDt/e68iTyUPN9V/4G+VSED3lZlickSlY2AJ9069SkZs
qLBzjCSgUNxtnKuvgNVsaHWlX7LPGkGrdKa71hNu+TsHJddyZJb0wwjespnytWQquiYL5Ioh25Lr
OtoYL02vtrMa1jwB/C6svWSJE4sZfCSw6gBjUBGtmSbGqQe8fPQVDAh/ouuvHNC83bGJeLs6hPuq
fqWSgBGO0y7h5dHpRclUUNqAZ+VN5W/Dcf0bHXCVjINR5kBLhRZEo2DGbnwSEfhe8FXi3mezSpW6
vGFDDQ2C/e2zVJjXmkKwgfZGngEKeZt7qN4KSlG4GO1klKz+8Q6KbsS3PrlmzUkI2DKMF/ppdFSz
LW6FEV0NWqBz0sUwjq1sdTWwmGyrYYo0kNBXTDW622P+p86BfpfEJRsjqTEUKHEIz1zJ00qM+f1o
hU0sc5o30r5i2FU2jhobEnzygBO5GcIh1Gb5pOL0GkSIzPuBzyBQSK8cf2LiGL8B44tjwPqXjyK6
/a+j2/oHKTHSBbZkTqwyC3dtP4O5GY3BIhIi0/vY4BWc8JL3S1PH5zYNSgzNioOA87PSXWkMRQVt
3rQPmR87lLsLeVijE5Bjj9WWr5X9p/FibqDVl5yMady4nRge7o437DOLg8uUJTcMYFr9VZrcOLdY
eKG0YIomgnxfRyeqRmXtFVYAmj2Fk3/Fu+HHGrwWEQ8yypjqdaIYKXXbGNkhnz1YBu4uqCgWrmbr
G+Bmx7BBsPF+KPcB2TtxAagFn/b5bk/wftJHfMCpnCNpQ5D3M8EcJL6vgZpz5NcbLhOu54GF4CGh
GdrZvkqz+xYtSRA4I6pIWD1Oa+nuV3TymnSZlT35sgCWL1SqPTqmUzjB1QMVbKML5OleHehLcDYj
ENi6ek1eUAgQSVGWkuEjBF8OAaTuN0F5TDHbdzxy7rGb4Y/haQE8kdozzM1XsyhoKBD1oKpz3hNP
4P0WhUbaAigxAOgyl+ipbQCdti4/+NQIPfw3YHwN0GQ7A9S4TcmsSCwfUAR5Yi9CPfXJJsjnvKp4
uBiaAbonw00H8aW8QffrjV0beKsWHfYbt8peuJDTUo0lMt3qE1Dlm2p9OYES8m7b/P7bNd2LVM6x
1piUcbtHqgFaPE/Au5nE2SPIoGuuhP2+veNwUoXB9AQKbtlja4E+iyTc2PaPKknlvIRRas1rTOF4
wJwjlKXjpPBfRYqrGygI3D2XzZZ+oMsT4tU6KYLo/S+z3osRfmo/Am7kfZWywJtywmhkBq9D2lrQ
b7rgeoA3SoHFcoSu8Ea2eziPYz5jK+sIesbLUv4Ng9Z/pbAJ13Tq4dJdzPnn/MFN5AaH7QDK/5wV
M9mzpGVMhnasTt08c9gjLANtooUBY9zODMcS2/cb0dAWlOkQIjBxpCbjzySr+M06tkiAJHXkv28Y
zcxnMRiwo3y9H3W8+lY+1SFFGibpe0dgI4zbVcltu4SR/kd+sKiBirZAp1RwLOBDUX86HcZQujdO
GaajtnZnZk2P0cO32z4i3kqiEmBWh2ocoeHsbRT9stX5KH/O4wDjOk8VHUpfUWl24/TWvEJAFPfe
8wRfrY8xusNZQiHi7EcMNpLGYHzjiAqNX87HprA3TTKk3yssD3TJcebECUeo11at1uVj5qZ0WLV6
Di6cJXm1yywfa5iuoeG8T6hNjsdJyiyE2W4+amnW39c8LdDeL/ZhrhNumjg3pdUVQFRgzZmUPzjL
27GqaN91yLsCk76heIi5F0HNr37gmvIER3wlRC+rFGk+wkM2F/G0emdU4szEozGCJ3eD2+UTsxQK
ma1OI90SAd087F8ONLPrWrTs+T2y/95oQjv8wIrocfGEJOj3AKpr/K/miPaYjM47bS/Us761ST5r
aXZiVMR7PJyxgIfphbAvcTq1Lym70/BgyHDfBHvLga49xvsSGtFmdwOm3C1T+GFPqhHv1BVQXsKS
Z61yPLKvSAhRTkPtiI6aJJubBR0jQP72NdOzFDzqkudeiE0Bp1qML80wOWQiTjpvAQ70Rpd6WE2l
GffPxmkY3X/vfMw5/VYJxUOUblbSl/sjgQDmyRoRFAFywpxyMQt0ay5Q6v2aa4foaHg/Fxkc+6yE
UyqLy4oysbEkitBAJ5XKQgzsffGZln8Zso7CnH7YI0WZhwSdjcKw+vNkYCBTMNOIs4f8/KvyJmVl
5erSWUIYGb0xG6jC6ZcdUA95AQZp1WTsG6/3lEKRUM4LCcudkDeyyERoWKOZRlXiympn2mlLUs1p
1AhB5f4+OIEGKD/jNlSAEZc2VX6mx311PQ+uCfnpbZc/Vy1HCHzQM5VmZCrVtxADVA0mb6Rl0oiH
eVtLq6W4VuQtqC8O6TTJL0YKF9DnEPw3W2AzvrzkSHhSwx0iIZELIO64ZNmRYWfHPprnHnxzIVct
IEOcNZfBWTMEkJQiiS+Qc8lxV/1jtL0H/qBKGrn7ePKHTUp3jn415abaJWvSFY+oNVhP8ks9MLZP
8if2PWM0CVV5y2cqeFem7ziw0eGZ2Xx8Zp9QCmhrZs1j0XmIN7eQOCbu+vdowJBuIFx+kQZK+9rX
xM2i3wsiAArR+qylhjNxFTcALpDIrlr0aRJTMiiEYQckWfswT9lLZaUYafrslqnA1LrZVRDF563b
RmLOIm6eCP+16ncs6vkqEFnvxFDBPHCMpZ24s4hnJ+w7iN3UunCZc+cfFc1LquoG+wleckcLThg2
8GBaFrEI83qifa6KyCABCHSDl/ach7AgwEGuDOg1RahDGvbcgalrlfoR1V9DkGvD0EcbcFKMyROE
Jdf06RheuxV6DG19j7eLZ7w7WIdYiQFLZ551xFJwYkoDfBP/Qqd40i/a4RaccLgzTUgXgL1qDla7
NbVAQxHFfdweboEhJPwlVkXYZJrdChMIBhbqnAwrykpjCSylWoDgdQLJ12mBp+sTQh9oadGi74lJ
j48SH/jRlbPZHCdVfAPtyexIK0826xilWnTsRjzIv1qIod3B6kOyxaelnJtL8TZrQBs0fQmv2Oz7
oFIJZ4A57as+jttNfMmnt/mm78O0e2Zi0cw8QwytazIt4+rzkeSPUXLN+0pQu/itZdxO+/uU1bTn
WZSoA0KIAKrlOv9YBwYBJNYT8TNDrrKHWdDt7Nd1KZ4oduIOGixwXLqQE4rLCtUaXdGZPFT/KnfI
bi/A44XbsEi8FrVcZ82tYjz+f2KUH1xXUw3CErmXNCKVuvpUisqRjyJSWgL+L9vkKAwMV5CLlGHM
wAS9wzKLxX3iluVpP6clXV9i32+G12qss4sJ6wBTE+CmZ0Y28yWWuTCe1XfaXaksVFNK+eRBeQbt
/V86s6sYY2K/tfNjqCYIn+3/UBAKqW3LFDQYQTBZXhm7LdCn7afCupdrV8jd15bTqJXO0YKvA58m
8RxAGbNsyg1p7UDLezDvX2f7312Klt4YGNS2zDQ673gGwAH1ehEbBGPhoKHjMmnJZ4ptbuhC4vUL
36PoPVz6txiHrrLRg3O1VDkct1qPA/ZNvIXG7xQXyHNOCoz/4lD0gDTRW8s+LOiobMQtFutd8Sh8
XiGR/QIhKlqh034QXRNwIFlZj6d/oYpbeaQ0tdRZ4qpMp/aJIrFwQMR2DlRFl6jZfH78gCfnQvdh
yqrJq+1gObs5EXfSbikTOf5iLS8ueqCTZmf8c//ajF3RWosT/IHz9BkPD9cnEL36z4ScUKImgaBl
VH74K8QbJJWDBRB30gXjkLykRW+lYnL2lOCRKUrqGH4HL4tWpUme4Yr9QBc2b43JPluhoIPWIkj7
PFTHEWf8U+ECG6DqdtqyR01hb31pHSMoBV4WKIeSt3L+x6KzexbCVOOSaca5a7unzVWRTr4CgqYM
ZkYKo73mqqyPJbXO4nieyFU99YQ5kZg1p9ksvY7YaH9ikk/5slPi1JS5BZKKlbTkAERm/OlGFTfv
1Tzy8JKxSA449JSjBUojgpUF8uCsx3prxHMarBYTq7v3lZoWHxHg7mwU+EEp6jeG2okPBqh780m0
6m0Bs7P7OGwz+k24adp7P4hjW3b3zW0+CA48iBnfgEhRD94eEA2jFyf//Rdtvff7HdHfGzO1cX0E
6sZvUcqZaPOoVSTYZK3+OcaSfH/pm8W4ydOTTsvNyQglBNtXu4+UvlL7+5NzMQuWQmsYP3+MRFBU
4U28+QxJu/9taJSxZNbOjloP9h3ixQkP0i3kBhTOc3AZTH6Y2DeYOLIwqa87ctYUdhQYDaBUdPqm
SVll0mu+V3XkLTOVO9crYQ3BInZ8LX4AHavzvJ90ibZfzozP6h73xlefwiK1uB4hhcGPhxBtYaMs
gVjlM8KZTD751eF1f9KoPTQ5X8r86pD4Yw4aVN13eViMBxD+o12NxtQEWW48lj/7LhVYf5iHUE3l
cAmm91VZNe5thxpJl4Vt/eyCasCWaCtzalTM5Jktk8fhHeIwk12hkz4mUjcP9XFJcFVh56ffYhMR
Ti4QyR64zzqIqsz8rAO/DXwy9lf86hBWTmkaVV2P/fP4bFOruV3ap+bQNyo46IUD9VGXJBpjA4vA
uhAcckLKhUqFcu7pfRem9BKZ2znEIIJZZiyiDpH6dNtf2LENHEwTkQ609EAhlu4dvFS23Dv91lnY
gjelgTREX6wd9ljZuLa2VRJryfz0GiQHHVTMzTtcj2VB1NQZfG91sCNiKANSkELejt4LG8oobpCo
VHTJ/RyfIPxqk0vtFaXg7VgVjFLp/GCTq+z/X9PocusnWVJ8HJ1nQ9ADPi6c7nC5QaPzyo+PqQbi
3N6blnseCf25mcXLYbxkZJpflzZp7zUEtA2hBeMHJfeIKYlRSL9QCR8rMqX7z0V5GEVQGOy7NuI6
aLoT/dEowgBdqX0dbcmQTMqDsMP4TFkbrRQXGyBBM+AeZCuy75SZ5oIMygLjOgS8bE9C3wjtsZ8r
1YvW8b/wyUpPCBkQkNrZFav8w7deZ+KwgnUtVwtJFiZQmzX8n1COB2Jgf/xFC13VmMUU6PryzUDw
gL8UQGGF1DU8cAkHbPHozT1nv+yDcGmNaPOyRJlATYxKn8hWEAOZFYLB+Dk2tTT545Fxg+jzu8SW
0q1iV4K2+pSiyVQqF3PdSaTGIKmFdMEmWEyC8mv0DJxuI8HXBiJ+XJdNT5eBrfolXaSBOU6E6MXw
LpskW/MvPGry5481Poc6dG5ZvEVIfSVX/zqiEZ9aEyrckIsy35vaeue2nVVK1L5YdZ/e3LarKPEm
hJG8jQ58DDKEM6WWFs05wYqwr+GFCPPkeEOutANi5OD1mfkFY8LXZ5DBkov9yj4XtpEmcjRbwSb0
Xui8ujVUhxAsWAU1EP7XWB0+HKQswQBCeu5iAsn+VTGYc0eiOtuEw48TaYYMRoLxrJre8hDVRs2q
k0awWYheMLvSfpAmPvAqtdFvO236wb6G9Mth4ZWluoac15Q+uGKFTpJY2MaT1seQloZczf99mgR6
9lynxkYuMvMea1Mtn5vt5XjKxOuvwc16U03MMeNWJAVVfVSYaY9RIk0CSqINTy/WATdRx8650Ru5
KrmslruuqV0s1ND1etiIiZXR9U04rAv0ZBTG599BbrPNjk7xjMpKHgLytxS6JE/ReatM2jQEoOKc
ZzP0GMky1/OThmMIRWiuj0wvP+EOxszPXHYXL9ATOnWV2RkrVNvnPS/1l2ihdz3HspvG5jwqiBD6
oMCTL6pypM7kZKoFrxzgQaEuGHXEEfZtUvdDmw6kqZlNUfTBrlO7aLEduu3+dwfdjSN9evyaTv5q
tR8ot64v/WuJ/6RCIvV1WiaKbcizq4GYPr2TV6NpZ9m9PSmW4nRltArcNi4JGj0ZrIrI9gg6J3hU
dr4bpafeQOSIqhJlP625eRkHprHMQWaPKWHjkwZfnT/poSQU6NetJJz0NLOEHStZO7ZV3lUnVgtr
GNaFwaOxicinISiTtFdwQZvGH/OsnOV76vs+wLQ6fkGm5OozdYe9ABOoLEqMldsKjnS4+zhsgUFl
+fS5yo67Fq0UoFdakA34jMQRw5bMBE+Mz4+jPG90xu9NJ4a8Tc/apTw1Q3D6bprcKoECO+/GoA8s
hhk0Kam6jyer6T7zbg3p6feU6z6if0a4UjQUPNAyNjGEqVzS8xRJ3+r6qY6swNE5HLbJDbSKt2oi
ufLeqkZ8Ylk2LKtMX6ICo5vqQkTwBd/G60fgkOkz+RzkKUzHc3oEg63AJ5bspTCNnCBvMaTk3f9e
QWLZTX+yptgcfPPzCmDaUHVJ64G+uU/haKN6M9sxUMbur0/xAJi36/8llItMdNzRw0cBRwcbdZer
irDUFq6kLWYsgudqYYqqoNo1yWT0z5DjuJjaEdTktzarXi2+dlxRcSVv3+8s65GW6Ei5lpg9MMaU
kJqEjp8LwD5iB3DIpixaExSD/R5WtKMuyuB8XKf+ZGoc8we1EQBL01Ey+eAs0o9mK4gon2qprFDF
bHsczsl53Rq7qm17pA/3GAjvEwjcaxzCaLN2IOv669SECc39qjsAEjwLAY38P2YyPpPryPpGX88C
xQQ5COM/mcCEx6j2RIl+PFdvmQYDHrpCuzda1H86h+MRtx51/gkkNQp7SGG2ktR03hxn0NxndkHC
zb4ZAc+v6TBsWclRr8tCfsB2g/pUNIiSmbnLMQabCbHxF0MLS4CEmIz66Rnm1T5bHEHXx3xd+xIL
T0gVMm4atofTL/vnx0vBjr6Vdkn5hvZxEMFeSa4ls/qSwNT4mnsrxBRi+Qjc6jHlDpEAe4ui3ve4
0Nr20Xkd/bugRl2a0sDN9tzF53so5h4vlgTZofotF9EyY1QB5WylfZr3YRZfjTP+BVn/KtiYZCqV
HXVIsbVd0q/Q0zIWsJrG3IqEAzAWZfjSogtm7/8XpS+tz7pEVKxcA45Y2OtW5VYw84qIDatTjj2l
eyusfS0SDWk77eCRwDU61X+Y9/11d18VCCfV48lUjF8Uw3PfD4sciRS+QN6SMk9PwHLrns8eMI+U
fuW+ZZQzBT03RDxLBcFLJbeJ5pFb1rEhtnBgDFwuDXPA0rGzlxbEIHgG1jUJCWtpkfMBeCdNO1Y+
qxVR4K4gs1VpD+/pNgeYVEM6EVPGzKmkjcCo2+8VyKKC4hlLyhMZQS1U/tKS8DbRgHE7Jdr8xTnD
JH7HWay6dOx56Sv6TgJ4FS194GGF7L9MsxMoOOafpB8EOUlH6Bb10Qy5Vl34J/tmi/7ajDr7Pvne
Rz+T6wozKPVNAMxYYZSuSW2HaTFpwWqjAWDt+U3AOt2znjdLiFFl9yBAh0H4rInbQT9cXdkIkFmq
obUZcX43Dkl55U4+LQgGNiVj+8ERdzm+DquS/e7p7X3pvIXLXoXMk4jgxArKuMHGvMpXCvtG3uMz
f5aUCrECdoKPhZsn4BxgULWMyG/BihBbWcSfUQGY9AzK6t3rYuGxRjNa9toBELyDL41K86xMkkbn
8mgjsvradIv8dJe9N5Ox+M4b1KukZyCRqN2nBjDKgfjvLwWuhNLsVuqG6EC2Nh41BcoX9DQ0q9bP
K8sV10MQ0mmuvWN3kMxsUr5YvlWUJ2NAgJWItR0gs2G8ph7043pFZpcr0WwsUmBdsA1FciIiDd5L
NWI2b548TIxugxPmhMBoU9f3XxCiaIOiQAcAwUS9ZoYDPZQrqjsaIOd3gQoiY4vZU0EsZqkOA5yl
W5aS03jeOSdI1KptRuuQtxBXwXEPNNbtVFTZil64RRnGvCElfNTMkaSZ81oby4EW8f6ibOM8uOlW
eNbAS6Qaxy33MO5tiEzqyL9EebcNHU23YDzrbbLGhLJ9OynSDROZfwREmokqpeDsxoi03hEyZ0V9
hEOvw53baEwa8uuVf7vwVdN3JHdTw6wjLBzX4KHZHL7w9grCfbGmrAD3QdPBOY2nMWRBQbdppLxE
kadjSSHP6c2WngfpoNWTB9fRLBMzE0DvYtX374JNU+CF/fPJ91rpcDrJEXfIXpx4Cwm0BLi85BnQ
ZqcjjF+Nh9rZLI7ovkLSOfDqNeCQyDG66ezkzY4VFvHWDCUKAftY5WmZRqTV7k18TgUW9XuqSfis
kWGqjcIVajI5YnHigmP0PKGmxr1oEpYCPL3Ii6jvRRVJaONk4vqpWFbVX8hULqUcT7IkN+8xOkEX
/e2JLrWRm0u9ESS89wRzdV+ypHVyCUF32vgwku8Koodk0RSGaXWidzag/xmtii3c4fD4u1ehFOCp
6mxdXHiHPOst7BkmXpijTHW4wHoPBJReNvqkmciufjbEd8hcyOmjLw1ED0D8gMPZbqHwadJRdCsB
4GXn77cR+6MaFENA5Gfvnmuioi25pUr1zhxpbb11H+qMr8MdfWnhOGAjRjjLlbjhtqiTxTWhn3U8
/HcFr2hZT57W2kU4FVleHyqNKwNM/jb2kg5Lu5KwUiX97PtmV4y+F0xuJ3H7z4W8jG5upTZI4pum
yC6i/QnAYeNewBXf5LTVsEg0BtjJRDxxPmBL6G0uzCgfxNCp+CCEXaYmrBFnycfa1JGL2yK8CMQ4
Sk7rBeftLSE0wssH3i3od6+WWdjO5Xo7wTlMZs6ot/RJynRjCjCHsd51AFSutzSAlTVFZTS7AkWN
1Cwju5XCP+O+W8NSPzNa+0MvibSVMdDYnhNUgg4mt+kLmnhtsRma2FKiFisa3fzvl3733p1Xt++N
sPNavvfdi74m3lns4FypDqux4aipDcjPxyPJ+FNJ/TieOvnHU+NXe5+rzVJitsyZQzxX3qNScTQu
UIYsOsMIBB0aIU76s2Wnp+O8FIA3bejhbda2XeGU/SA2bEx2DIggI6QG8tZOUQ34s0Zd9sJt/3H0
TvzxxvsAauBB0+oYspJe/TiTv+3rdcKHi6mAYApkVWFPaSHRIO3kt4NNQf3qSJ+BlDcHp79pxeek
v7oSkMGpuAwme1FtN6nZmXXllwOE6JL8Oip2KzaoZQI56dCCLv3z9Wf+DWKTDN22l5S5Bg38aYyS
i+ko1OMj8E7gOuE97p4bUYnzj/wbBF0QlVcj5PHcfNcuG1yFzZwx46G9KCmRWAnCtFUtz8WDsdd4
/3OvkcY/6lFAdDyzbm7l680DVx+v9cpOpTwxUvFAlYhHXao/cFAOmIJZRLyad48tkhT3dBGd7t+w
h9lWZb/yQkKCv8Cpztu1zRDdmOzqh+0YCxNv/qYncKzUuXkORjhrqheliyQnoBhyszbESLjq6sem
TUk+T81y5QtN9JYUDsRXtLBEbMShfz47cNGXMjCTYFIG2btkLJ7hJXaaoZKv9hfrFNlCrZqqLe7A
jUGWcLfgDoncNOk28vyTjt79kEHge5jgyy/QaVapz31cidxI1By9zWON8VZFd76DHuy7gQi8qNOx
tDAvIwGwn256eUGUUVLU46+qtSY5jYxvT6CNZubWyzVSCG3mrTxJohKd5YAIIPjTxrNo9vD57qOq
88319+l5E/o1S8XETCuJROBWP1B8NtNJg+T+4OLXSpCZZSon7ow+o+B+UOzcEHIwDGuOYkrxWT6R
ewNDgpH9VZ5K1kBlwr5upTqtnIw3Ka+AoO1SQKA53ZVw+/MpYxrEYti1HmhbIfWo60JnsFQS1aY5
C+uqTlvIPQplqybjQczu7DUaLI3FBbi+fTMPHRZ0cnN5hTYfHcxdLmLB/U3wI/ZBezzQUP3bDQr3
Vdmw8X4+JmBz1hJ4xb4wDIkBlf9WalUB7gQfTDTPIdkuNO0gIqylXB39LcW+L9u7r5uD+BhyoRDg
twtMGtmXCqXoboNb/FWZc28vLYEH4oPd/99xwWwbxSjMg4U9cVU/SBP4HZs4JEQ8zx+MXpfqp7yZ
efttYhPr6vGoW+rYOnGz71h9D/t/MdUEBUOYTxMj8LOTuDCE+f40nTJy47piFCUklU//7cH5f59a
rEiASKiI7xhBC5uIRfkY9K82DSwcQfCIKw022qy5sBpuNOnOIEHRVLlZUV91cYI0NSplb6FUcTn0
hrM4BZL0lF1Hb2EsW1ob+uJ3/qy2QgrnziabO078wW/ipXalPTTNf5Yjr6PwzMrvCH3Hcl3WiyA/
7QFtWL14jpDBxy1wQGYMC65kmryvQruv7gEteMxtJQisMdWiWlJWfcXBwGte6Ex+xg/FHcmqCHta
RffVLCRYPWP9PTK8ELKznyUWOtSuEBKoWZ1WlI7aHSa3hErtF/5BYgPWi/MWunbTe0F/nOKgpn1q
hoEH02itqjl0qnVgHVO95uL86uv2mBMoOqMeEDwHIJ2jPHHo8vYVaiGTvYwGFxew+Qo195KrUy34
cMBXZ9zaeCrmKI/spOYjjPF0YkfiD4pNOW1LEEl8kYJzKS8SZfLUgJvqG0f8fXgEIccWb2Puo91i
BiKapVUJVqCEgnhVev1n7vxraqNS/dnOC0yNIGIC4DjeomOjmyyhl4puw+98ogkwEEMnWUjnHc6D
bCvtc97G9IFuijQ00Ka2HU7dJuGJKboIisctzCi6+X1Bd2+syhag8jmvLgF3dHzlrBMBKWdPpaie
dQXc7Ot5r3mEgent/o5xP0iI8WYyAhouLVWeHjHT4x2IE8WdoeXCJX1xgQp9eBlAsPJbXMir3pkM
Klww7UHA3ylQyce7jbLB/RIG+Wvju6rZ7yVVNHx8FuzN6HxIyaNTauvTEb2n750LpaqPqPCCHJ1Q
i62lVeFKZQ6owa9I+tQdU7obBt9uWsYb/B2GK5RLp+yDkCO0Ay3g1v2LWsjQerU2YAJPbhr8mf23
XOGO00O93uywZ8x/sTKITpvOrPYU8luZHvUDcB+5DLAVxzougp4QcQZh+aRNoesjP+NokpTSzgbL
m+4o7rBCselsW9oVZbSLrGIl8mRUeKoRxsKRxUIEUc7W553Ise2ZB1Iwik5CNoNDDiG8TXGvlL0o
ALXcs+ZlMlqoomdJ1C9lxM/BRnbWinpP7aAMYCaE210JgpgsLACqpig03a+nt6YEqVdUE002ZmPX
DkEmGPTgsaAWpFxaXjUmfZaEVzs+jKPFnzeB6Sz7S5NxKGMeLmJoSnF5a9QKfewBXzr4gIGV8gTF
HvFbAvwiKZYtZPGqxsHRWyfVT751QsVfJtQWFA1kozAAgC8Oc/VdPQlUpPGc0c+vzQAkOP3hz375
dNh5UFBRfnvdIlG2gIo0YG0Cmji3KEKKVLAoiR2c5rImyMeQYedMr0YjVhuxkzzQWViLw71I76Wf
4XH7ePT8MJyM8Yai8GcUFWETh83whLJ/QbpaRCvg9HW557/M3SYl5iQ1sjt+pw/KLXs4Y6yd6jU1
QTROdFMvIuIe4O7rRFOYPD0uXlcnOM8qbFceCVmkORPf4SvOdlWIXdVgTvAfMOuC6UoHhe2ipXZ0
s2mBeEYTlioE6N1rA7dSljhX6YgiLWxjmM0Kq3RffI9f3wA+5Q41EqHagMSxTL0kgIkvSROQHBZY
Dj2DyqToCsW2gtKBevV6X5TmDPFPRg4uF+DIeVXax8cZs4itvIrMkJnt/lP66Lg1hWcl3xpErrsn
Lkw2ySDpAwBQ0YZFQoghHn5VEdlRACZCzAb7/gNDmRKroOGBA82TL2WbihVdcP9eVjmptlPDJRru
LpcpTH+SFufYdrk2iHD29fJn3fQNUlUisfbAjhNa6Wg8zCou9JIm3rLSFDWYH03Czq3TDzueoL9F
pyLUoEPbAFH0t9yIgV4oIDAWA0iw3OG+3HMlY/2eG5lxaaIJYwsTnA/FrKBeY++fyYrXzHvoasib
TlK758z6oohc6MrMZ4RWHDQdQUpKZzuYSiPqm8vJlqHrKDKXXAFlXCULFqQ7sBEx5Elv1NiprYaZ
Bu9aB03E692tL7ivfGoQQLu+6oCN62O0Is1fahyRgEl3bL/f2So2C96rZL6kTYrzcNdxJ7E+jPob
s0vqHnQGZBXYYz3QqcCCrQzvqmhU0OMjrUM9cLnOSvLr0qz70y6GDEeHlOdcKtL9cRv/BNXjiM0T
C0vjUTMoATmmCKqoz/tIJLesM31jYnjVAdzmzSk8IC87seF87+tD+hfSh0RKli5Tss9SKxUYuDQE
YqNlfQkUz2s/2iLAwC5Co+qrRVzNsiBpq2s6YL1J5U08ypqZGEmRGyQQ1VIfV2ECxEUxESN9CLms
QrXoGtiqAN0jV8FpCfsrb29U1SbzCaCtREhLcMFCVgCal7jE6UAOHCan1VNcD8OV5CXbutoa/TbA
Ejq/G5naJMyPec46l4fWX4YFqa1JSg/CislZ2t/J/tnPkVg3QupVTGdUp+92TlJmGlitwYIWDgZI
dMLUiY6bpOoCywkZLmaqt31TJ8JItZVg5a44ju0X8K2JiwvgOJVtQRczhkrIOlde5Tu+4UFfECQQ
Y3gsniQoTHWCk/862GDYEyb4+9g41teBwCnFCMoC4kgU9ylbZCaf+dXfovMpcKa3UaN0TbolZCQo
XHULnTy1z3SqZmtBwUy0n9Oflh7Tmm37RgkmFy14viizjkeUcl5anSxu2A5KteNhINjteYp6+l6S
SGf2iu+jP91UcSJHQt6GjySw2UT1T4Zc4VNiCNPKJ9XDK47QukM+dpZRfjHCcIf+1yocOpl0bxf9
FYaXsmnTj300J5cPZs3OsWH1vgKnIPsnU3EaW8DP5d8cfumXpRd5c0GmRYTIt+4rKsZeDBFupD8n
/iCcl/dlMLwMDebIBaVGVmAsVtbpcTthdmd0qc10XQjCNNe3VQfr2/Xh9nFNdH+va1TDJWrLoKxU
L9NUDccRqIWEzoTZ3PX4O1MQroK+cGYtwabWZgNF2cvhRuRA9/KjbIR2m8PZaDZ3lT4uEhHyo7TW
yE8BX/46PqO5y5GoWbDpOA7tyoXafBER9uBlzX3MFRQcqe0laDAp8zMwqfVhxZAMpURHxjxEMNOp
5em70pYvVFk11j3Ae3GIrxXengP7Tf0QQBvoWxfAI+2QbI4x84VDmB8OJAQ+dI+THIzUtdSlrAcF
0VVodhOc7DHOHWU9M/g0zniZLRIJ/oouyzBKT4FSu+jpGB9G8yTpwb2p8AlocQKkFLys7M8w23mP
AdjyTdztUhhHkzLoammXXDeeRurXhvHTNmyeZ7qx8N7igWRyhvLRR75sWmnd4EK0oFJmnJdRVmaI
bZ3zes5ztfSSSvXla4GTO2fD8CP7KFm6pyxxCTjiJkc1RXi2SIs+8wvYYS7R+f/iS5NET5Ztf7sZ
uEzWxuIMc4nhujAoZd+sI0f0rWORLGzeSOFq5YHeGcmFvqyP8M+KEQ0086pByvODIpsRf3I8kxBo
4ya6sXXUvUgXeI/7adxPhgC3Ct/oNkv4Y2XkXM81eW/xGX1ntRuqNNfJB3qMxcqFFZX6FESqPl0o
tg1DvAVWUAf6AhPo+eTs5N4tPoAFBsvHzsAblPyCc5WDYxrEyVDOeJShJf7cwHBHKD942Clr9txA
TVvr+oro5NV7ZcJ9Lwa6xBdP8mjNiTd3HrbsDpKmkdhoQkFVgbKaf3W1mdVnqd5AxJ52/zGmHZPc
woc5CspHFC+UhrsaWqJ6qdqQoFOEFovdV/8vpd/UD4KZnlMu8SfC8urbuc0pPidEOVUsBpXj4Tqr
0uJMApcR6gLGC5BhxUeq31N7kqPtI3nwZhW2Dw3/sD5/3dxGnr/6zDGx5ipoN3o3thnBcVYVFVik
RuDW+SNcudE9LrsBTfa0pZtCxCrNRShPlOlA+4D0eO/Ccpq0gK845xjii3h9cskNAVol4xnNLNsQ
vR86U0wNj4dY1mfiZaYw6VXlWS3+i3/6ykL7uwwBs5BumEIYB0nCpXpcJTCPjrRpOVWoUcbTe/mu
L3dA5oZe5BcihExocvLycEwT1AQBxi2HLPYm1liKj9XQIrOgKBpGVNGB8EQlwMWTTeKKmyCdnI9z
CWJ+HgVm8NNYrCfc982AzU8hicvfT6pYZba7vl3jzDdnW3Fdp50T8fcewmcWUVpv79QYpt30QxE7
j2w7pbGWf7TZn6TYiqhrK/PT1vauYYhO2QoKJWhXUiJH/Z6gh1eYysbTGi5fCgbYOH6s2z8GcRFp
uMxM0hEWjTXsvJaWy98LQPYBYllxvGV6V+TiQVtaMUlbyoPiaQgrTpleEI2CcoV7d57HynvVEDid
4eA+SWXZhOrFlIoITlh4m+TzSropm0LpLNhGhbisa7+IE6nlgYpJs+AW5k7SWKSlFdhJHKsb48gU
+t+XVUBG20fXQnWa4LygiprI228Ze/EqFnxr/vLY9PaMrTPiC9Ju9AA7lVsZWPe0wUYWbWSJJUUi
cD0gbBe159FOnG3pE55ae9TUF+4RSoxF6dVbzUWmMizJW8GKknec78hAPnX6PkLgu2NZ7xyixuG4
hnMERDT5C9OwhtAoAuJZsTMNs66ajDpcwSXC4fOLCuu8lOr+m6tjexl4L5TuQZcs0SRuO3sHRbiW
bcWJ4xevObA0nte/cjEmOGDSQ51/lzNtWbH0vOAT51U4F9U4qenJ+zxFpfv2JaPTC92OIkgIPSm5
T2WrQT5wX/05N2rSiiV/ahpN7vRn9VqxQ1eqpaK6aaJHU47S4FyYrvZTK0WY8HHb5+2ZkuGSiLHH
Wzy6oG5ujRerK/rW5nZ81r3r7cSXr0IK0QIpDPUTqXH9aZT81JfxjGXELsHT5rMwpWvrQhfSVGO2
tz3k4fl6b8rFitZ+6H6IqpJxX9e2td6f7h3bB0uqfqojBmce7AHfI9nr24Rjjf45WGbn4EyTM/ry
t1Gki+D2KNtvdtVXVWDvsL4mHBP632D3UakGb7xZHxzqG5N2jgaAXVr0Sxp7RvNL0WJ+5X+Yus14
i6BzMVoqJfsJ0dgfr65FZRhL5BXRiv5D3oS+HLC29nrYTC82QggAed0TwmALNtaxWJsxBRp5t3l/
KHBBlMtnB0KcQ8jY6XmodVjFwBSht3HQQ0Ha2RTobcEZhyfIHkOkh6cu43iQjzRLFx1FN+Mu6FGP
LoFlCewRVC2dt8G9WRDod9fvTy0uP6OCjGagUiXhHY3RY4FNr9jAzAcDuww7bKkqVvbFSeMsHpEh
1wSkBZoOcL9gU3JluT/2qOzMNhkZtLehuK07Z7BbozX/6iZwQu74uzfby2q12d/9Zg97COS5fWgH
isHSfNA1YOftoFx26Y+K8HCbk0nj2RiolWpUSRmrkhQvpiaru3xw2V7Tl+r7nXpR0B+le+Ky8z3o
8yTikrMxDhx0Zv0KFL0qwwUQAURpD16U/WIlOIhB0vuQjr1osALdrpDn1M3WilYh2bNDc1+rDDa0
1AsKreHR329YA00vFqFl2RO3FzWx3Gnhj/1up8aDiNKPqsayqYjp2yExis3APV11W8otNoktvp0F
9lsw2lqMD69O/rBEhGXKoKRgI2l4SiUZx0OfTNQXYFPJna8N8IjFTzO646YR+ms1USJM+jeY78Em
tlcIds6Y8kp0sta2sjTKzyUavI6ieeMxwMRWCJruB/PcvJ1q138KQ5HJqHdNr1KN/Thx/m/AcWPz
lmhMfrqb9Ph1kd0crVGdiZ3FNur7vaC8fffvZholjL0IPiKlosL8SLsPi6AWtF42ANEvPdR8mlbw
rfA6z/LHoVA8JStyCQADg5HWUSDaDKt+gAT1FZSrU13/cbwGtqWhkPeI3dXtxBeDRFHOq8FTD3Fd
I3p0lAXOG2T+EVEggUwDIPETeVMtM0rYUfdszabrQAA/sIitPb6QDoG0lhC5sXX4TIZeSNQJw3jY
8kCGtTvemyNjmp3RI/94ESsi+xjjWUnvMlVd/+E8d+M2xjEE8mDGrNcz22HwN4Agq4USyNIoEh3F
znqRKjFSeceZtt9j9CGdx2epQ5t3IKsasrA8TXPeWA4xal/ui28HpEAExux+UazzITB0++Dk9CY+
Yrj2DqiT2wQkKlbRtAj8XV4tAB7J14vGyE0S3jFFD14XUhVgZjn7/EiExE++5SfaWTVDVhTUMpBN
CStBbHvFZHhODvNJ05nnH7dXXCI8dBRnnMsLTMY3xfKGcA6EYQ0B7KduJhMYGZZ4NGU0xZKPefWL
QBs18aotykWspCuLghjEgoIFgraVg8bo8McTGNTXTvCZQA5KRdWawCo7YuKOL/LAuKZR1XixiqWM
oUPfIulybyVUe3YNCCNcnO00+KfJrfsLrbUlIQlYDTst4xb8w+RcfSvMeY1XAD10Ytxvut3S23gx
Ceix6DYZoQG/KmolCE3n8S552cUqtr6khvTIf1qC1MtrU1TQPTfOBTFiYXrKs75nwgHoxPVNC5U1
d+ODIePPURO1pQ6Se/Qvcw5yqhH4G7fb2rWuA/pcE86JqyElfWOwUPL14Lu7QYpd+Y5BBZCBo6bF
tsv64QtKmWovbYFoTOGEalmkxpalkKbVZPb6nOHZnveSlktC6fZT9PnGp4KTwwT2xa8n9lPbvV1q
AfGN/fMHtiMk4/4gAhcL6O70nduAjCGpVG1ipZ24hXg+u0N9XMTKPVuE45JcLiUlgkfvJ/lB4qnC
HyKRtoA1Xf+WzmbSc5Yi4t24S2urPo/e7QkkRcuj/gOq9Pgg9SKt9M1G+7iqn4MD15NYQa9a4Fxd
huVTE2aTRQDV+SwGqwzseM+fSm+GEWsy+Jl7ohkH2A0NLvNfC55jCfq7ctiJbiuLKi9W2PTVkdYF
PdqktxJDB8KSisd2XBw3Zg7kvA2iQT8g4R+yUixdFiV7Oy0FKFtUoYSMokF6A4gC+hfVb7vxg9ie
28tXX2btaE+jIjWS9W+hOCc60ItpC45SexxSRxTfhdZv/Mlec8aaVBC+zLrGkRSTHDn4jf+2mjgj
d76BePzcKYEoWcZHUmP6tnTn7NoHavn/lR+hXOPEyA6l8JhvyaZ8vzMzozCokJp09mI2EDo1iE+w
d6If+9c7NHS2dpDDPjbxOHumigs5g5PwAtuvoRmZDX/Ul8teXoDsjzfS7432MbSW53CIoFS9X7DR
WH+2sOhOlsRxBWgY78JL+Eq7wzpHD8ZLEA6FJyBbCSqk6uxBgN6R3s2AyZNQwLjouQGgSzXh8ph/
MSW0P7nZneA1wJpbmaM8uHjj/DowPWctLvGueMnxXy1c1sfKkMflJMER88eSH0M+CFXoB1J4mNeH
SkLURp5HcKXx4MYONiYXvLGxXF4EwkIMT5D/RXMPBnFKkU40ZmyqFT7cX7CDn6yTp9Ow0QsCmE+b
Cb3aC2j2dxG1yVOPUz0p5YVl7Zx+kJz4eEpJleR/CD3WDf/EIGu6lXZ8qOP99+ZV8N/0F9Mvtr5b
CcyUOG3z7TSKo9N+4L64VoCc18gtYjyDDKXrNEgq/EQeks5bKVsAVbhUSpK4MDJRlFRZZ/qragE0
9o+KJCtwHwWo+00C1DyX5yaeyQanB1IKGHtovPe2ZKepLXQE+5MLlvnSEuhw2RDPwqRz7BPW4CFv
5Ip7ZBZouwS8E3sXHR81pcbNGjfAwyS4TH65YiZi0Wpml5yUGnQ/JFbI6LapnYkB4ttzz1PGXIuR
oeHmFidrkFWLsl+8SZjDVSznOG0mg8rOc/hMkfsty19tb/kX+HussXcIPUrogeQ672G4grHFrQ3w
ezumQ7qvO14yGGorzfy4p/J3Ar0TmnSRZ1zfvAbsiyPnxUO+M5LWSAK3GFbEX4i01cO4XHWEwzJP
gBTFawkXtO/3+I+sxmw5OGbiDtXOlu8yaOzuLmhKem7vCixdHohJDKXrL585XWbh6lQowEEyrBgJ
8A1iKBbQ6NrppqasUzBefNk1h2tFHhFJ9j9JX2Tck3H4x9JRZo6tt/HN2Zy345OGL6CqJP4eYq0B
NzBB+q2xcz/52NaJoIFe9eg6BoXUzvnSQzfivsUrIA34Jt5d7Ia5BBcqwh02mUUZdlLWT5z8nMLm
ZXpBwxXxeB8g2ce3gzZ4LchYBa23mG9v4/+pwz777M9SkFcc5I7RSNEE+7Sf/ookghgQJ6Zj8Z9w
01aYIZHef+Bmt/pq225qvAdLGV+0X/Kk5hdH3qUm+Zv8Hjaz2Rrc07g2V0SC3ca7mczvWFltPS63
BUc1Jklaf7N0gxctaZFg3hUM+oLtgqK/aem6joLJQJf0wjxs//340OY9soXvow+JlzXd8+wEXDBE
Sucr9EA+gUJkJvUsPa9EfTCnVvxQsxWwYDzYewTGdx+1qLbPsXnpExJk0M44VM2WyhMK9TZyqib8
cHIXkXCpwPQqiEMxstLePjJLjlLEejutNSzPTeDRIFzcaeS3lnJCIxEBcglNVAxVOWjG8EhY9fMy
77RUQkHvO64214/oHk8WgxPVp7Q09xWeHpiXexaw9FI8srzTitWHstVrVfWW/WC9tyDkTxLmKBRk
YOaFUnbRKinVNpH7RYVN5DQRoOq+2TndRT7i8d4ntDsCyDGQc25VP2oEdQX4qVVOkUJeJrDjiqZU
XL/Wtp/Z+WLPg7g8FyEB3fGA+95BSJFGlRaQKpO9aoKrU3dG3itzsfrcSQKJ9OB1BH6xX+VslQBP
pd9CkKKEhfDWPUb20tmuKFBgrpY8P7VBcdbVO9RM+yRGjRcGbgj8VIBOPYk8z+P77SWd5MYfYSdh
eRoA75rsEoGsaqrLVyZJGKmMvBuDEvy4UzjHB+adw0pYOEJBaXGqG237fVrfqG2oeEhEEdj1t4BW
om8dn6OlwnvJztDjfQ/CXRGX74gLZP6lcmKz0CUG2kEKiyclemh26TaNqrt4v8OZDXvcYgEfIxeh
53NUY3KdCUSD1NHYj+wr/9ibkIcYVdnaU8R7fqVpIRPYbdxQOIKIuBC9aM/n6/OUooGsV9oKJjpr
Dp9Y2XxJ4a7F0y0xKEN7cfmZuc9ZoJ/b+Br6Sah6EML6Ipns00rFxaUGr7yl01j/c8A2Xhxj7GMC
39qSnQ84a7f+Ldqz9/hIvEpI4XnwB7R8iEd1VtHwxOqIyzI02xZiZU70jvB7pk69PNXpkGNIBbKb
Ojs8ch0kb2xzegwXdwxieADYLHJOFcx9q0C7vVvqMAzbYHKc99Jz5kbaIUXhs9CC7Uqx+M2oFgBC
Gj2ZEFsp0Kf/o4NbRAASlb0uPi4By2sk4WOaOv/O51vrngEsyYlaoIePpn1fQ6UyzTF0m5hfgUff
ZsQaBgbHHvioB25sCZvjya5B62jdsArZEXtc8F0ypndmkafwjZMbzbXEgUE1Jmx9xe1uUrosIquv
N+7xa7wdE5FoDy6us+G7CI5v6KfHBicpLDABFYBFYG2UlxvXnEOdDRO1a+2bEeoj2A5Z5uFLF4Jr
svVUPuOYdZubIc5JpdwiKYsYEFoOJHUXn+33NJ4FS3Sxz5g9i8yJ9DLASkbqyK73VFQAAVOJyHI8
vI/5YkJbt7FiM6+/AskkfFN+Okgh0DIIU4JanR7qYomPkjPNEUfxWece/tRVqJR85yPVJ6MLB2zb
dwHe6nZQCfvvV5EucBuO10kZd8P66MbYjEzlZCxowsy/CfkKzHOLI3fxufJihXIySu4g6LYTJaZg
diTx/L2DN8ZbR+1D7NZ17vyc5m1FWqxmUZU/QYnHWB7oGehvZm08+mbv2+Pws1ESRznIbfQpfmGB
mvwZiiRJc2k2OCoGV5UyL9cYgIGVn+mZKbZwjg9X6e31nwzFBvQwgsgjK/iWLiSjffoGK6ZJwfju
YKET2GXZmQ7pwa+7kBj/VcKUbzeca1YtzYX4qgLNju/ct9X9Mj9VpplNzUMbvuPiQg5n5Uw72zSv
51TPPj2IBLNAcsZawPOkRaCJr6ieQbJrbXAUV3mupvcbXE6VAwIszTCzOaE4X20Rj3N5jcvQ7/YH
6newsFcP9Q9An2AcNcNzhmi2dmScfFp/Db1W3g0/fD8sJVFi+tqhf95vVCVncWH/wwwlXCieAS3x
AoP/LcdLmbHZ+9qoADYelUTZTe5bPfK/CSzWWX75XnR+bFKIkyOKxxu86axdgiHrsAg2I08vt1eV
3QQiXU8PW7xbzEhf8pen83zMiCFiEP6ei/nrPN4kTgp1AGIKbbsMK7GphrhwMYiXVOZ0Ic6EmyzI
OlBwf5X2EE2Wvw80UKIfhOxyj55xOWHgpU0qaKz8+6FV//M8VyZuco2oOrky6/eAzb91H0ykZLpn
njnei32vRym5krksmOHLV2dAOXFQqbzWQYp1VkoMqvggKvcfgVGem5stw7MKapXJc9KXkf2CVr3R
DRFr42bJkbiaznhK//ISB55IKqoklDnhjCtqQkEtCeSGflw5tstDB3UYDmp/EfVl0WkdqK+wRHNu
Tmrtty5lKg2bYv8DJ8C0y1qe/L+twxN7oRGVkGhc8k0Td3RsT6SS7WVpUE8FmdC9tnINoVKe85Ro
LgHbY+146uSzqHId9EXPVyUjTOZFRuWVCv1HlFUXZj+Mnsk1pzf8RoBCBBsDuccXwPK2WUdvOmY2
+SwchjnRaRUOwGo4s3ZdQpi8hyIKtptj4Ap6VfUk4SmwZu7knaO/JCuk6G7mfe4a0+gQeK4BZ+pC
FJdwLv3ECwfQyNbaqYnnneqLuVQ53Q3dGQHL0PtQOpSOkgtzK12Z91JGYOpuMQ9skG6/16BZTyGi
nxtw8Nlo8rKAISSaJ566AOwQ1loqCgq1s36kwuFQzrCvCGm+KCVoUGm1r/Pju1E10ot2EEnqE079
gNAvcLfMy/QYtu3iJsNXK3JRZLRadXpGXK33OoEl6hwQmsX2rtCc6rhwzU+/BRcLfXQXsge0fV23
zPBTM3ouuO7gfdaQQoT60380NjkpzT3vUx1ZxBODsIHFDtgpljnWiKRxhZHbR3curR4Y4CRpa1wT
DqOjNDs/aaXKVFaQw1U9FAb65CxP0WKfERbdl+j6XLxJHERGse0LI5I02tjDVD6mn73VwVwQfa0G
rx1T70Bdb31JsuiRpWtPdUGroQKFISbS3SUzuPoLhvFq1c5xu1u7I9p4+jk5nauUmlOc0gjdoaDM
LL+/M4/PrwALhsQfWSCbq5QCGh2Bm3W8kMjzuHNjjmdTVpchEZBrDooNO/iwfeVSc4/cez4Vcm71
hza8ez5fjyYrWxx/nLy+IAGyv+VQyJEvYhwh0Da3eMCI8J5C0IR5jcwmquH6n3azHFHXGaGUHjgM
4mAvSEQnzJF7LEoZBz0EL6C/e93mkb4Depwp2lLwNWswz5YyeJHkQ9+/UsM1Qx2Sp/EE0E/nGWGw
A6CCOGQ5gDKSyCq2poLYKmiew+o37B+2mkqkDRUejjWgR6wTwVkBUR67SwwdAq/lTxwuq2ikhBnO
tshaGy19Jfdg/0y111UcoLg3676IYhuAjWOoxU4acULlhWNNfpr2VWuZRKb5U7PXSD+eTsovj4JF
AkQqfk4/moD20xz5+wyx7Me7YLJSKCXoX/3gozXfu0PlNBJcVVri3pHJVXNZyfmgp1eaD2qrKBEG
7di1bZjK4KVkpWGrJA2kuvn+3kWmaXphrHs+BklitHaxTJUaaG7fTLuP1ck7OluBsDJ27apo+BdC
v+sgm7L9TKoYlmwLNv+1dvRDvwNN8Dc0CHFt8D71VI2JXvOidCMdydLl/zkgs7sUwufhcP55apFn
UAL+LvFrSMnoXwMeILaupiplqkhXsVSw/HVBC6COq9YDppT1F1huEqYMLCI93TUfrUPzy1v7lRcU
5pFxTRxmpxIzzGloR7GfpczV5ypCnpM3GZXIeEUzx+IoCpVIRjwQ35o8Wom4ocKvU93pU+gReZlE
AwE4FPftpAYp5L79/FLKhyiEtFuqeqDfuxgw0RSFJ3vLumVA4rjuaiOMtde4b9G7vSaKvlkJlWUm
KsrGDRmYj7Ecq1l9oKzWzhyCrpy3mpOZm4THlkhAAlauE+98yXZXp09JX3xn1LiJ22qX/MNfklIH
kcQ60SJ4sKfu0lrnSN1e1b72rU/YHhF348SIPsPA0ca8nB0plFPG+rq+2gGB1fKvhQTzQDjzzTpE
1EL3QvT8/Wyb/62rcF6OcNUYdrzkEh/4PioeOr84lpWHJt60arw8oH2HRaVQHBgbJAu5aKWfH5Ok
PkTSY+ny7zRJzalrCXp51QPb2vVqADUyzMPzX3mCcAM75PP7kmawpz44ug/OeB1WigUtsZPXEJgu
cKbp8d9cDowOzG0yVVuZW9a/Ryqfq2PruwIGaFiSWVJ2nVjXOBnd866Ns62/7ahlNWfE/6jB8bHi
jfS1B5b7wgb23qQslbRgrNbRpIoTkwRm/qjB/FE9xfqSjN5G/44loeMg8eB/13B6ZPtxtFnhNXXf
t1ZuVe/Y5UXhUSaV9jNeHY9xNxzFR5f7fKMsReFb2LBP5F7w0goWOz7pGgRaCuTXW0jFbjyek772
QbcQ7PA02QmviZHtyxCWRBYlS9BdgZf3AjTzkGRiuLE2DZ8R3KY0sktWmeA8ck9lzI44DOZgA7Wt
5s/CZJjaCjHFUkPXjaCWC/DLxc1qZU9tbqF/zT1ff01SrsaKdfMhCoVaopz/igMWU6oo70aBHlra
0u9ADhOOxRLwifqxv7gwrUloxCt8u7SWsbqIZWqB0gt99nK0MU0yaTHwYOasFu6RCIPJ5wIuRWib
RKFBk/eNixKp7n7JyEkd8PaU8reu1JKDZcEHII74Lt+KXg0Mmt761MpAZXvNlFsk3zxjo+kfE1FN
nQsAXeC6RPVTEMnNgxqgP+PMgpAb4zs/Mjm8UyLkVKbwFl5q0IvMmGgnqu3Vv6+6zi43S6IzolQn
DDhBXymFvDxOibDGC4ddGKGHzgxj2pDRLC3Uh4pLCAG0rv9trnUXns+btwjxbDnX7p2mCE7bgAcv
jiHajgOQ6MYKO558RtlrmEY03IP/V5Yuk/rI8B4JdCsJXvNZfKSOlDaBlyFT7Q4FA1BNhLEZ7qLP
RmkWQT4XK2v30p6fey95kDV7pB90WQQnYUPzxYcYnP+ffy2Ygt4tzveLRDNkYfl/wkd6KSSLQ7cR
AiwbDGP2qd35ytKOuns+5KAgV1p1Bp3f6KdR0zbXhh+x2+Qosw4fYJHy9to5lQh02gRDBHrc8IAc
q6V8UDgrmi7VcSLOqve1QYDO9SXoyaFydJCAuGCcwEZ+9A3VrZ1tTTRyENh5TB5ILulEx6M1ht3C
T1yktGQGVLxVADFJ1sqsUI0kvx+bfPqW+aC291OeNwTlEOu/OdAC74BgwJ2NqgvbO/r/3NOf9kzI
92Kk+1qmGiNbfNK9FywXFHsVlcnrkQPMKl3ApCXe9R2iZn4WRHsv/BI1MOoNkjYq66NizUvRdyQM
YplyJJdO2dWgBNS/HU7XgoNQ+DArX5OtfGahi22cR3sv1HGm2ovONcSUIIf/qwUdNzpVWFO9i0tX
GyI8u5sJEuyr/St6QzSDAKsIt7I/3ivqolXLhHDOZeACuJaSl7KAehjeLAbKETNZIloGWIdURMfU
Jqjr3lbqt4E17MVT6qeoh/j0Ze0RWkv6YufvfAGde+4kZJj/pNSnjvKv36GREPJikfF9lwe2AiID
LjH2gvEd3xSEYmn7a8C9Ubdx8CxtHRULnkd7sH8ATOa3JHl4dPjkZYkO8akgc04IMrTveZ23fb6p
E9OACRRowC5AKzV1mK55BYiU0lsLvXp0XCgMmXEq65iO/QWNzBJzd3R8UyY+goQO/+ETT15nWpTY
BXcvkdPgAw7iNSwABYK9WeTYrzVRfE1Huu0ZV4m+DDaVc97oMEllJTb3cZxjlemPEpP1w06Mxiyo
r5lqe8bMWnm4BjeiVBIkAFnKcGaOpFGEl8ggxesSSpASmTskADqeqSY9/uxV7I4MFIceDEdrtRoJ
/wh6QjJool6RzmP2W4jiNFNRAiOlfG6Mzq7I5ovpdfqhOS+r6QGaAywA+6vVPWgq7OoIRPeW+bjF
M5rkuBkuq8/Vy42mxXSv2fejgYaxdWapGLPNF7rAwQW2Ve7pfPt4Gw6Dygctle8QAfmTzXCNOWVZ
puAyFFUkaGsOmoWXEleIDri3S3kPP/BlpTjy6C8r24VK8X7Fx7cnopkACNmwCvxC68KouNxsyKMp
7TLt6HIrN8UfhqMmh7VXOSaocwvva9taE/A20KnEyqoBp5r/80WrYwH1xKxu3L63t+5haCrdgebN
j+U0lJUFdTWziVego7nHHcOzpG0cUZXGjBX83lpCFKwJc+TUScevFBWpesIAolRpxq7Efd+kQg4w
v384bcQuZ8C5DacoeyYWzSOTAgLiU7SaOb8R86CwpO5z+ipmW0yRvpeEKMl3dgYbq9JOCptUGGt+
cOaRk+KE3U981uKpzFrTa0MvlDmQCY9t2M6zmSQHP4WBcoM2KWB7EA9UZy3VGGUXZ+enXynVZ0hh
wTOU5HYVQ+8G2VNkaa5K5yJ2Nf2cxkOV2Mxa60bISGdsPOBUq87Rs3GdnIHG5RQ9fXf773YOvXMn
tdceaVsBvnyrUK8uzcGqNc3qWT/aRYhqp7F9ctKtSiJmnzYbWHWmEqw/Fif0veswhi+cdwNAP3ml
3mcVHtnhoUOwRUiN4DrhvN4GV5WSquw1LGdQFd9XzWqM4WIqjB3tJTPO6lmgIkYkeuGsVfduFTo2
lp2VXCCeMBuCt6tETY2HQ7MX76NuUgCLxEsjIs6meCSzQG+PEwT1knN67dx6r9U/e9ibUCSjhqBY
TW5IVm2f8oFQCQVwfl2Eefdcab8y5dYCGfnJBeJGw2yHHqZNVHKjow/rgUDzv0SvrQKUiEQ88Ujk
1uqW3XISJ2t4Q3dZrlI2Gcd5zRuoiBvkXRDayF7g2FngcWq9oYXAH2FOCIZ49V4VqcmiU776/fcW
zec6h7fxDConnZpNNgOT+Lq/7gb4R9t8UhVbBygm1X0coulluIGOHWFlApFP1mosApFZ+VR3319D
oMREc3sBLvx29yag4wzoY+rUJ1WN9dg8EVSrwD1jg2EAKYtUDq2TJ+fnjd1YELd7Ajq/RYL1gK32
eQbdjMBNsJgYk5h7sn6mKPgQW2HYZhPE/PbX700PnaMcbQLgEOLmx1IPcU+1RbdbhK6GlxKToG4r
CQtOVQogp8ae8MYedUp9QlpuojFOMdQDU3yUKVKPEKB8vwQsWu1JespVAvDx6mMR1GNqw9Xehm8D
azay3D5E+ANULFRypcIxZ6UOOsH8Fdi7ixdFefZXDNRYP4TmMPb4CZNvM3MT+M+mLspTyyU3f5Y9
oUWZwySqvbfDijpHfFJJGIszmPAcZgWC7JphSnEI4jhjcyq3hGQWUR0KPAI9aAO+xdTksMIXXmZY
N3JTzwtkvjVSviW5/yDiH+Zbne2Sct6MBvQkv8blsEtSN228zGBRyccmFAXEB1d70NIfzLFX4722
PFKG58dZOug9KuNev0bXBzNfno1YrwL/oT5BUu1sWIXGmCu0cFr/GjRkDVg8uklvwXWD/Xe4bXQV
xQHiqlQtfb4wkMTFRHXRJOZhNoe41qLA/YMuw6D8IqpDpnJwm86RbnJCcqkwpdLKoqxDPjbvHfhg
DpnZmB/wVOkP+qLPp5sxoJm//YjJCfmCMLyXCtGufKSdCAh8agEtwSTTP53A1mx8VAHxkl03a0qh
xZrQv0X6U+uHCudxA1d/7/Ntm10QvCM8P6wm1ry87p0OZnaHyFnwLDzFyCm3J/XshepFe5kVbGZC
ybhX3qj5DT4OwAjGkLtr3ICvOxY7GpzUb0z2IJ82kiXctWSXX7MCevvaYiDwHdoIRgdUtElNNl3h
uefSuPBrcAGTNI6PnZ/uQGpkOMRyY7TGkPH2ZqTgjYTkkwVdpYWRLd4Boz4WZMdYJ21/3JJbjsZ5
U9pV1tjtTBTNvlMKvset/1slxGXDjQQQLXk4+eW7BINdkzomnQcwQp5VdP72nbpDpGfEPmzXq7ZA
e7a/Mc1IaWkFnmfMY6SQlfz2Wi3jL/5EBiWZGk4GMw41pp3nuv0nYYoTsAdj2G1umKhmC57yIpqC
2ulBHohv2AN0Dc2DzwjKUkQclOiONDWXlhAEBXJqCJKz7HhHnKq4CJAPRkiOhCmbIcIrXOLKjleE
djW89ilcE9HqFzpciCwu5HRefpwGB+YbWqb87FUgrb6AG9vS0+mYTWPinuQHwywcwfUNhhl8qNKQ
iqAyfVAykaAoiyfVLl9b+DA+4+LGwP7Y59KLB2hglBcwM6cLNVkIDWZdggqe7TZiuTlm5FLIHUwH
57nv55LS44nsB5eLkycefaZwcZEw9435rcl4R67CPUSowyuDz/2x/cHwEZ4xjmbTsYdm5Glo+UvI
ruf609mFFiUtxXfzb34fgbGOEg7qo2bSKf5NTJ0dePHn5B242f13V7abt3WDw4T9mpLbSN23GR2T
2gDvl1ehnlyVMenl29LGDuc2hNmF4VbALTVtL7NxIO0xsMIs3kXAma51n0EJzwLYNHaKUiZ6dQmX
uTmGSOUmc2nj7hHyG4SKoI+bSEA9T2eKDlt1uhS8kr/11DX0nsGkD2pis3WbBNAx/TWEgwdpJSU1
XHyd2QPvecL2Y8tN3/R8T1phqYfGtrT/aJgjq5EheNbIBJnVpihrULxsnUNOHeiAxG4lEcfaBrAJ
o5/7X/cnTAzfMciykouKwqz+IQjcSEjUhsbgBnh+8p0ADwekJTGvelQnQtpsIVQdl2kLuxu879UC
dufPLPIGTG50cw4/tHPMTLJLDhmu4J5883DTAzn6qFMVNvwao5wT2PPFjrq4V4u2c2mo+s6yHtY9
JmTi+ZZnXWuBUGzrhtRvr6GcYaJbNlZ2XLFIUq6AdG16AvNP09JaDyP2KHPJP2yMwc/UMCdN/a6J
NoWIcFYAyzCenufOJn4rS8R+YDxQKi/DdBE0w8m8zvkmbaLmQ5ZkYXW4qvkIZn7s6uf7L65Wfbx/
gXQZ8i3bZdJdQIJ1bg5T8bfjOYa5pyeUYi2zWphIUOVe4sbXa+4TxlC2RVMpZeFF+8MAZCB7bBGh
1VasVw+x3Dc5dn/lEGvOX1aPovVY2jxiZBrpX9cvNsir9CR2DLgG++Zswkz2sEIwjnseiPqNUjuV
UayPnHKY0HWXhewA1SDepE1cJAqaN8l2zdjdn2uml59UdoTFlcHlzsIndA0TWpP941kSl83x+iY7
nwmpR+fSbqOAdEsRVkxwpV7IDPVWga7TgXvIsq5xMkbEUhqyZyvcqINhpMkehcUzDYAp52Jixltk
9YVR7LNKxL50NwD7gZT1HsKVaW0qKU0jGl47VzOVJQwYtHVFuf9i44l/tKm4raPDZhmroZ2VeasB
sQIDEkM008URg8QOMLNQ+f1YgEQlaYWNhfn5bmkUMKyTWbl4NJ+qLDmqmIUmN14Ox46tdyPjwZpX
EZi4u1mQZSkTrryP/pGjHdeeqfrvCZHYLomYvTI9uRFd2UTlxXT7r+ErTjxcVVrB6XHIn2qV4QB4
cS29DJcwKhcWDTY8+9FwCi/jNBEyOCw5iGkdWhbL0W7duct7fpaQr+t3eNXVvENL8kHExJ5o2W5q
cEOUWNeYo0AOJH5KeUvLl/sPiLqdMY/CbENp/svEtjE+r6C7Ej85tc6BiBoN2qE11Ru3XTlZZ298
fP0dQ105quxFD1Ep4xLxoQAI4Ji6AzCGFJDGg8JRhP3zB90ukDU4KzAKYnOLctK4GWsV2bj7bMmZ
1sLkSJj9eE43jvqNygsG60EPTRed3k31DcafAMwpDv8XIM3KQn/yNIkJPZoBitf7vpzvSYOkGQdt
ChjJRzrznUHEayC/I7tdvOod0PUwQiMqYF9W/kyzPXyJEKdlXflKWSGWmzMX+lRBdXG+ISC48OgY
zH+UY+4fRSM91YnMcUGSv4xg9l07U7BO9suskRmZL+AYk1Fa9BMyI98nfa1CSQwbE1nAYKC7SBBR
FP8gG5LoO+elgSdAfHzHpcQJNn/47n1qqZCGgydcD18tR7HUSaFaBZbhcjITjriO5daXk8luNje4
b/256K8dH+pzP9qQNyx9a1ej5jam+Zhglp8C5jj7rbCnpNbMVvqrCasRZDoFW1xAEROMltejDGqt
D+d76Fix1TncfQWykNXsUdPO3Rj/0LqQEVKppaNEY3UYLNwyaJJ2Ex2fZqlxxYM+TiJRVSknnLuH
h6UhmMJMXKkkaUNHjKSuXxQMjHbSHbUp4P+QKt4ORTB8WGAJwsEWUd899P2k74A7/nXlMfGRezyW
hI62gr7OaFTFMbvFQJj/d+PFx8vE0IfPsV3bV+A7mVVPuXkA5qa6GXk90wlT1fO0FFjd26D2wBKD
hHtJUO+GCybeB9NyZhE3M2s0GIkRQ86RDzf63gV5kzx/liER51U7cjcQmM0lC1GaCgqBRSUKjpam
WCyl/MMdKFdG0zpull7oCQbF97GUnuFV4sYkiunDXU24TMwolkRb0/ya1QNR6kk17q5/p8TyTNd8
k1acNl330wo1Es1QRpFxuPPOOFRzZpCEw5rwBbCGT2Fu7Yg/NWasLdKNxyD0i8ahJYJb1Hp6oEqQ
68w8s1c1ZGlkX0wxZCKzD4kLHpRlH7Oxp6Xj0frdkJKJYrrHB72yrlMT8/aVOHBKGi0fLtdyfXm6
zQd1rh2AkHqvnPNim+d9OHn+RIp57ItFMnZsM9Jxw7Q8oqxjPt0hecgYtf79S7ZvAJ/JYNBMjNpW
C4+kToeQ0CXQKkJ2TZlTd+cg0itZr82WIX23MQc//BrQ51swvoWlmhnT9XfWO+sUz6TKI3TtBFSQ
qM0rEXf/crRi9B2aayX8FT2nQ5Q33ra8NVEK+52iC2f6Ki/KmTVfpGccPOTqjtCPM6P5VhNx+nkr
XUxf7wcci3Ck/gElSBvCUAqzs+HsEPHeTOXqxn8dOb1knnTmY4fMWjS1cjM/EWIXttfLS2Ll4m8v
wu9ZvsSLqtDxoq/sDeVE2q9FWRgMwSmyy3XcLxV1m1DK2THK/2VRq8R4DqEVFWjar5AHdgB+lb+/
jO0tyswP51+SJ5a1A7jwGbHtAixJoPIYhBw6AnWO00PBTtwlB21ns8NdZ9zxgsKkrj+Ob/M9QqZA
+mzNr3+6USQ/DTKk54zRIDmS5ZJNgTje50gfvA0JGUEiqxnlwAHTvNS5VYIJdQYeNHPT4bCv+ZPx
TOqZG2UeGGhdP39ohjrNk7UQIyema7lFTNUCh/dgDIkFHTZJfVYSlVUXs5UQPqoWgmzNA02S/p6N
uKEIDsDoD7GOehdeoUf031xn6Yya8mEbCN3Q1azmBX6Oq9pnYb+Yadyf4+hvOqBmYnSc+CVb0fuf
zfiXqwgH42bU3Ke5SR22odj0vrWJmCrlwcvRTmasXbynbTimUJ8W+YIJuVqk8EnRimd5Lbm88QW8
yPbucceaLx0+iZNOminIgOVwIdUI3IGo/Vr2KSWipeBvGW6cUA6sv8wa7NdmwfzzU4fhSc8iYPu1
jHISACnIrNO+mthy1b7ghSTGgBm1+1axRlsel04IsoHIAdFT1tI8rS+aL+pLyXt19eM4Qj7uSHJE
N/uB7KvE3WpNfmcfz63rBV87dmRN5LzzvBHlcFaPk1RlT49CMpcGv0jNQNtZEL9ByTgCTzDmqm6K
TtdkzzTfC4pg3CZg7VRlDHXQ+oiLq1eornZkMF2dp7ITbh5sPFupO7+JQOqugdjkaC0JaZGX27c/
3N1Cp391NogmI1GIemJ83B+OWJUOGviyCw7ScjHNh+Fxq/de9rDHzsJaqEIP3SgwXV99r1rWVpYR
HnABm1YHpMxZIV2KPXMcU73s4SlmvV35sC2+IZp4V1npyM76o8NYPlaMpw0Ztmkpn787wfWrWCDi
rqc+XkXSrwEb3XQ+j70PRGKoZD19b+RWM3w1BQP2k8tNIkzS3wbOjDt3n9H6ckiR4V5OwWSjj/y0
bzGkmj0YelzPJpydGuY1INB9iGgCKOnWAYQ54ihHcFD97Y6tWBjrkX1vos6orro2pDUK8BzB7nDn
J2LYvmQzltt763TEXaCNZuv58+lPwBHMMaMnxRXSrtMuS5qT4qW2EXzO+9YSRmaj7YYoUqyOXbIo
RrROlEjOB5EpIO6LOH7OuxkQvPPE/reN3AS/6j5JFDaAUeAAmwiPLpAv2oZ7MmE5/boPRPpMNYKX
V6N43fMaesVs6uHQNwwEqA+xACzzdOeEvPXobwO/Qtj6l7NY8PdG2iLDTXNDeTQppbGAfc9jy4H6
fWmG4GQe4mReKI8JlLRXMx747Ucgv/AWyoMMF6FqbBi8f9zYzrA2g01t8nzSsaADizAjFIqHkjH9
L5oa6YAvI/DkFSZSJtL4IfnB/NGl3L8kZbXBvQvTnjcFcEXhi1Kg9cIr/CAtHjbY8JuZWNJeX7mv
2YC8jDqfzN/SdcpjtrpWNEB8kiziLDwSl3+c2D/Xd1/XA77dXQHf5aGkifxMst8c+5WNnL+cpmIE
RockKUl75eAm3VAoqUGW3kfR7Htap7oUjiVVUp2mix/IjzrtKsN6jbCceWuguL8Cr3xOOlt7OtGJ
szvS2ZJWkafuHwb2ez7fd5B1oO4U2Fje9ssTFlIthf4RZJ7kOgKcexp5KD3Kz/DIb51j459uaws6
9uBI6RtNTCrKmcs4lF87MYjUEbm5clZRzXoXmtL22qHkjXOTEJlIdvrWdx8WCgWaTcNPx0EHn9r8
m/ZOcFacqQh4ZSLYIME3CzHjnXWgA1y/Hfg2zDTy/iIAUBUywUXT+qeWoLZcXgoFWtJMRMzBAMm0
Rkrp1GRfpkP901qzxYb1IPZVAWgWmqRrWxf3l8zKDyR32bta9WpomP9GSBVQIASWRcq9sqyVaZ3j
dJM6083EONVBBuKBTJRAxB5/Z8XB49zyG+AJ2CGRluYMJZ2D3oJemNjGAWUOoEH/UjIOySwfg71y
5o8VIxFQnf/WE+MQtVhTvXEOnK2pTpR+6/dYteP0G+F+LvH//D4GIQQ/J3Y/Qg1XSaCIRnGZYSq9
OygMS7hUAYM5zDtcMG8X30sjrKJ2EsdFI0rg/hm5GHmFhzGWjgn19aNy552OSBWUUr85OFtvqOjI
TCc0PeJzjs1lWAMdWhZord0+3/Nrhxp+sTmdhQv+RDCa1gf43gsejY7PaPt7LqR4aTLKc5doYnua
xIBazFiELKeqXQop/RTA6UyvgJCGfQwR1BApwPpLS5+z8UeYitoBMcSo+mhhKxXdPHM0RKlO8su6
V8IZ6cF2jxG040P3OB61/TgnEN+Ax6I8LzH+yUxQQNx1ZXrUpTNulu7fWKH4vBe36pP8AkfK7jlx
Cm3tRGLRSYw8SxXcC4oZP+LWUIIqA4n9hq3LT/tnQLtT8Ls6Wm8lKmC7z4O85LRvKpE8dltIInPD
ZKBZv+RjcHJUl97+uXo7zl7Yh1LFYwn7HT7DG+NoYbrFRDDDLRQubmGAR/MAOrgHPTrorFgMQL5x
NElSyru41Ay1wUg9M5QZC156P3/GA/NAXtyW4sBzZi8fqcRMpr/VbwAf8s5HFn/y7RBDxiYFcuCu
jEOmz0z5vx8q8C8c9bn7xaz64kDD16Eu5Sng7ImJ8jhkEYOa++1w+EBceKiFc8YxlKC+x0pOzvRK
VohwiaNlGA+UyQPlh1MqHKkY1++Jdqxt51aRuj8yDh3Sz50O69naqCmwfPfqfoQx3Iya7lHNel/9
YIsiLzu7MEAD/sGDxdbhqbHf9Ux64G9/zUlFNIRdXqAinIrGBT1JjVPGtu0KeeVp700A2HOJlWI5
GDMyGioLYfVu3dy2HUOwPYqZeSWOoBOJk1w5YGZypc04kVgoslt+KDMuB6GKBbF0DPl/w12WUQiY
zZYoqocpBafCcJ8QdJrInEbXZlF+7bhHHZxqIaKOTFzzbgbFLQAexA833yiCe897sDi47omOs+Ls
mJP8oBXXcrVMoslEZ1rt2ghjiygopBo6HoJzZoTnrr7NNUejkI4IRCRrqe72tqEmhQq2WZGy4GhD
0eMhAiM8jq2MSYUHbqVJSBkdZslvwXELmf/Ud096+Xm5J+i5bd8HZV8kj0ODmwlLyKUE+EBtWkBn
aNnueHnO7BZyysGjvFIsMAiXxv/jJcS0r2Ozb0R7YvYYnsDCfnW/4SALyLVeakUkBpHBPreHnp4i
4Mu17ZL4dRq6Dpe7pKsZoPnRcbdIivliQtpiLGh7vz2oL7wPl1DibvY+gzJ8rwsqRK809FlcKumO
c2S0+6dPoFk26L3IgC8GDdb6ds85hPW5jl750UZ9UwOdmAKLj7Fp2IBJRp6bMniCYreEauo4cPM/
HmAtblZfFsfTaZtalmuWDA2RHjGGnGPlIWMRqvbht202hylMvTphZKo85xLdKkcBSkmdjq5RoNPO
qgQe9io2+fPbWICPTstRjk47nPkg/dBln9pB9cCzD8bcFcbnQhsWioJRVUo7v2HzKg4SJ/IUMg+j
cDe+dHQeQXwS4F1BaNB/N78BDsu5hly4+km/7Vm0q8jARNRDTcbyIunuzKgD7pYFOxC2FTGJ7e7N
SYP0srwfps9GCXLCClflrdXnoQH3dnyhDQjuQzv+FHwzTM/zRj7BvfyDGUqSPsvO3R11kpiTmE7k
uGWbKkYWTMv8cruspPZLTuYtkTvpEc2FoRSbJ6bUbU1KsQHuo69hhkVOULWedjcIl+KV9ofllDGI
cqwzaX6F1iXST4RU7fznFX60E1l4kR5yVkBG+zth5QLfF6h96F+9gByHLPrUiEwGaL5D5l5B+r2d
wkKU2Fa39xNP9aSLOzSkqzeRh+T1Xg07KOXm+GiXu6sBYA26vU/YP6SkBQ9uwebwcyo8sz9JAY2L
FlDN8F2/FgnVvWBInMqIUPQg9nARhl1GcoESV7akCKJsu7+hT7W/kUYN9C6elwqyutHB7tyVlWP/
SYGw7Nr8Ui4d3cgsAXqfg+ps0P01bV+c4p2tB8UcUX+dvoSGjmrwEhUYrKMWImUaqNBs68/UeDHd
nr8T0SrxuxZiqgKTf4F/DoQBo5fD6lFInHXOdG12vygcKPWd1d/t/1zbFIZw0SONwDL6qNa65UGf
mlkEVu+mrQufzDaCoKgydcm67y2JEjhBIoi1WdPl86HNc7lXzuE0MvLAYM6AfhEDIna7mG80w2Z+
2I3PgfNGNiSNvkhYpg/pemXIMXuvFBewpqbV9hLlrREWVb0BMEoTKtcnwuaahLw5q6TEfXK8zx0h
qKTyM4mSiZU0NGyJ664bXDZYUNzcwSlNsQH/QY98ATLsNVgvJXLzPxNRIxXn3PpwIX8NlSHn4TbW
6VMpdhI+F2psYI6vUgMB4RXEPS/xSwz5cflB0S83biQYLi9Vd2nwlLKHR8ou0tiwjt02mWm07xLK
0wEbymZ8zel3M5tupZTeJbUFZCF6w6FoiVC74gMdAqLXna3ua8Ygf0xlAdc2flZhJA8O9CzK6ADN
2OMiWn6Fu060fSsP3mZlkltpMUpWu9PsUj1UQuBXsuvvhQwmZKdxH8/TNwDrK3P22PZGT43W1jIk
xNEC214RRiFTmnWmZEK6/+Fplczp8GHt8IoN7KYOwvO6nPNeiw3VAflOb6vZeOu7neFW+4fXPSAG
tJeL05I3kZ1pjgMJ1+hBG7aIOHJYojxNud+CcI5fK1DDX1znehh9jwkw/Pjy7V6TI3vl3skghWGo
iruZTLiZ+gnrtm4ol7Ia5wbaOHerhQL/H19CIujXn3N87NnELrFV/EsCHEXkjd1GtDt0HzQ/CSxc
FBd6G2ZPeea3rTSuy5uuejkArTOBzhEfTvvm92E1YfwQ0g4IdHyA41m1Qycq+/QyUZyenZK1wD9O
OA4KEbW2F+LNNozFvERsCmTrYgIjv6Hx+WhyNdTFOdhpnVWQKKCCkMnh9zV+AF/ZPLqsnvqXSVPT
g66gYEIbzDx4eliQh/rbtD2WQKzUvjfLMpNtEBBV2ON0UU04bmr/O6AH4tqzOnXLivsoiXc63dAM
URGN12cYPdVXY1bP90HiVoTmtYBx0aKb2t77yMUv8/aYqOfHfm+ZifoazMLdb8AYI90/qRtKrXjc
wOerTfHoPDWzXBSo97w7dYmXKLJzk2XmvyQm+mJi5NsEiMpDDSDMHv7YhOLiyj9MtdVcaLrVkU3e
6T9gNq8yl8IGjjPdlDmHoMTwFzd2K4j1L1SUfuouSCNLc96Slh2EoyF3Rmyiody5DL2pOA96P30y
UKpfb9R9z7EgyJpt4VO/pmnkY9xDWnRMIz8UA9gJbkxoecxgAeOvfGUOBHer8hBJvm0+9hI+orMv
Q3Oi+G4BWlNUzE+RpRJjw0wlv++VpodJ50zDXtiJ/i3MeVksbLTGzik2IB+uyF4bl20VBesBVLBp
uzL9HzUUcc075ioLNw6yrebi2rRVAHC0alvF/YEyIyc6CMIUC2qziC86mGcp8NzIMHm5MH+gWFTj
6uoi3oCkYUveVZZvJhs0vMBdFBYhr48xiK/tbfIgiwwwd+9vDCyFNbx89Ksdft1XZKTJgyLHz0hU
wEk7+qI+URR1ZMt+bJufMIWQxUi5BPOTurRTLCNfJy5zq3kG6mWK2wiCtjl4g7y8NskHfXEj9WIC
jZZI2GapFD+i5oNSTopgZsJpkk2zFt7D64j9ErecAk1KrAIB/M1DMHWfmVG7yVsbi8jabTpQ3cy3
0C9tg6JX4LWid33G+bLJ3yN1uIt9zERyvzHJKVHYuJzQyo76EoWvOA8op23ZtDX7s9YED8Xjz1sP
P1gk50P3JkXXNOTnt0JUDPIiBVFGFu+NlLWAvpwCEcnKXHakzOny7yYrkufLdChMXJMss9hhazn6
9Srq20cdojtVtKdDogHqC4u6o95G7MuLES26MLc5FKsOO2+lwEL6o5oXsyMATLCOYvZ8a1ka0Yj/
IxFwJYi0HC3V2NdIdEfvhhhbZZtLguXrWwzV3Fq8donzck0SoDRLMYZxgfvAp8CIty82Oqc/r9AE
Tw29snNMdn0ZyT4qve+GBDxvEfQHCoIpmOts6jaCdUG3SkOOArtQRryCxZRAog5ARHzjK9jUWQa1
oEQ++Zf9ozFEQqKaXDhuJDFacn2G/2rIDhY6ppjLWYxyB0SM+PeCBXwQm1nDp4EHINCjxDzNSMYX
7v7WUrjauammdyWMAtOFOfU9ABxiRoLEAOiVOuAP1NQDTMf8bAKlWG5U89cW0xBtZ9O2AvlxuiOS
zqcXMMWFslNM9G1qTMGOjmMm2Fv/IJKkpiH05+ur50A6fNSuxrScu7LinxpBnnHm1rIpZtcRu98Q
kXPTZkKZAFP4rwUhvTo2wF1kE/UfK0yKlTWQmHicsZYD2YikJ2y4b8Ho/nclwmK4HH6uc3ZrmeNV
zIIaz0aOctXir/IDRNKr5nUnjxjoBFyN0JNtGseZwuFSBd5u+WYq5OmNaYMsO9RhSZM8giyErgaI
3lyEsKU08lJeAJGwcIfyFjVBWySVoRPcUO3H3yd5wvWWr5HWfm58//H2X39cFTjBCMee/GYKC9Zj
WVGklCOYZ7m4rZQf2cPIg+1/2mVr/KvWM0p71+rBCkRbfk9of2vmzVYOoAR7V79H90ZkQUw5Bx2Y
YE1SKI1gJ4HTr21Mg76lZH2luMRy8kcPzrbtbairfTdvpEzG/UVkYEWflnJ0ya2ZUDy1ufyn7r16
ceCYAlosb/H+Zf+9SfXSHvYAJkyElUD7rbzlztFs3ZXOUJ8Y84GRxe1bDCMqzTc2NrQ3VzOTbxo/
MWt0kudKZRLyDqPG/i23mUUkUSStXWHnXnfOcE6OOTJNOjF+KE7LzAPu1vdWNWw3iIMTLUQNsPAo
KW32vGkkXIUpxRmA32slFqNEXxRIlpzFXNdqC06CD1j8G0cY+6DyUazkIfsOuNE65V+n0b+9LLEv
M3QjkFAK3pzW7djkuxlt8uD1Ifq8fBTM8Xobf0Q3gqc9Bz6BXBehX5DVqkAkS3e1RAba/1qE4JQf
7CzJKK/ayzNTOnOFdjrp37fB8LDMtmg8kHoviGrdMHTPQ/TwE1I8Ii8YJGTnaptUKPVV1ypj0gxo
nQZdoWiF9iBomtpIH2ihjElf2eEaeGfRA5CmvfcjEVJ2vETx/ztJzl5UtbQgubkYJGMhTFvUd777
UsLP+SzaVBijiJgTGmv0hsyBBGGKJ/llZy0IC5JoXOPXObLJeEhDzCzB9WdJmqrWrOPwXYo147Fd
GcgviS7cWksr4VuXnPK0puKpSYWEapBGOa6tTMhhMs69ILyinUCpwI+0JxvS8moTZmY5vdGIAp5W
dBv5dZQxFaKDdg6QwE6wNyyRKxBFPppGKmR31Lgw0Iw5eqo83qhRvRcRDw/R0xgjDR9jsvbVyWKw
nng28Y3HV0YvPanxNG8vUF9uD/ZVm5iQax5eSjSu9ayVII6eOUU1PnM9rE4G9TJ89cgNz4osKrx7
53KugdVzhtKdz71FnxaSXUbruasSFLTXQhCa4BCSW+BMf5/AaXr8Q2fIEfVfmo8XyluLEukm7cn7
fyzkvU6Lr4UeU8yj0bCfqCpQrvCWo3kwPaZUR6J+cK2JqYp/q/AbffaPC7Sd/Qhgl3hGSwNzEmeR
SbJIFlda2s9ptjb4nKePxYekrkrp6iNlW62vJHSPxGFSTlJ04C8ckSpOXU/4ACoecSKjQJRsZEVl
7FfnIltHX49QUdybf3BO3pHEsYathJwX+pQXQIpWPplVO/SV7f3X5idV1Mep7MFQzkyszPTud898
Quan1PEkoH91/Q9x2CI7RYV/85QU1Rrpman9Q2hIaLQQCYugqNscpdpEjB9VW/EyMI9N+p4yJyGG
5n8uGDQ+u18Fwelyn/jJze8f7cEUy8yHMMJY8OiTPZOTm86sAWsDDVaZhuHyNC2xvs5ZUMkI4hIp
p7xVmHmWwev8HBt78SEIrsTB1pX96wFNeTBMdiBoe4TFLpF3EG6n+7lv8Y4BVmPeaQC9jfD7QGlh
AQIwPzBv8DujWrk1b8a9Q8nCtxfDxtw1WopnW+jonwZByQKTq2qYnyTG+P5Bkq7daAlKEUzUPIlO
43FH4DlDbv3nvYWAxpfPqtwunkQ7NltPVA1m2bsJdTujKa/XctgjvlB0Dkwbf0UklBY8TFqY777Y
WUGJU5riPEVluFXbLY9vIw5L9/0q9hEd8Pk4hz+0rmWEWOTos8q+H4L6L7GiUqCmAUPUjHDJMl4L
41nuqtROyxGQYfemjKdeioV/0QuH3NplsZZ+SEYUBv1QKtMFcyErYWldW8fgBStX1n7Q2vLvI8+x
89Ej6BWhnLuyrQ1//YmoyRBE5Kcync8/2NuVvE0odyYKf1L4s7qb69pTYQXjif1qmcvZFbqIVYbd
IOLJvJbDhP10ViXvvlNwOYCkHdLl9ueHHnzeJjhXbKy2/f6P4xcklXTVFK5nE04As0pNYLNqUWLc
Dp1nSiN/cWoCpLlzSugNQekwQk/EC+Sj7CwK0k36mINU49htE+E2xyYpby4BX7haFnVNN6urAhYy
nAXMiktMUDoVk2DxEf8Gv4JR0QoFXB1c8S4W6WlE/akOVbcvu/kSe1euRbvm5CCxAVPumzBWnDWr
7c6KFUcY4I7ttGZXsbEDBm+YJN1hAHjuW/1yapKD6F9VpLFDwWnSEsdhZR1kgdVOkZMY9gdoBXXQ
76F1tcY7ye9B0oZjYBGqLgcIyraWaU+tg1/rZSWPQLgTo4XyUkzN380iZ4CV9tOeCT4nQ24bTx09
rk/mJFSDQ6BULfrz1MROiURV9CsfVrpWpljHAdBZNiEHOM/Blh+e0ah1rg7Cqv5GbZJUCAtpcydR
p/eSa5erWwUZ3MPwSPFzSRynEf1RwGdI6dvIRh4b1zr8q/GWcJ3WTNpmRQ4MjHZFPj6Stb42fUVh
od+Vb6cjl4+aQMC+TCYb9U0bg5AoakaurUwCHDPWWYiuKFDCsolb5LmhacuA/uIws2reLWQk4DoD
mwJvlkxoJ38buDSGbmRYOF4EPg5Bl+QgdTbinjWvL8X0boeV17eZ29cqY41u09ps74fJL5i0V+vy
4zhySD8Phy6n6trPPGubRRmjUtW/QgiXWDWNHliAzT/ieT2U8oO1upCQ/X1Alb852UyQk0YESS+F
pYeQIHqGOOIe9OnurRhrA8EVz+l/9148TL2qc3SVE+Bkp31HFH4fDQA1V3CaqvLwsGRCQZetRUKK
6Ec2ppJJko+jacngN2FPR9Y0oDrsI4y835xkqo6+vGa3+QtRR/xtpeLe2QyLXU7ZgK1OTFvsCCtg
XOt0iQ0Su5IYziaM+coeta/lFY0OZSZ4FVqqivzxvHYedFofnLnDNMtyVSgHzIS4T9E+knZpLiDH
pOXgqSdtNTI/hcy8C27iI1EyxbbBwWjxf3mV2oEKxLAUv23ZRl6XhDzFQXbT7Zv+RCAq/OJ/O8BM
tSYZH7e3zqK+TQzsb4wliLndRmmDPdHwaX2reRTvTfqFPjh4op2LDC7rMb5AFBxk9OMUg8bbIpSd
bodzDV1Cg3Cce8h3koK3WT0dBT3gTouoJ4jKSHSLJlwc1oOAno3RfJQP6CmMU63rER1R0AxMDv84
Wl2phCW5gbbTAmVPFRiUyfnYGkpaYNOjKpNVNezNfFSfmgXbWmR4QEdaFzdrBUhrevHuhKtZMYPv
6ipCS3Xz8Qt1NdOTwSyEe7V9VLHOunvm6MWFiKOXucxYY4P/XAk0vwsT49KawVcFS52sfGypgVPK
zsA2ASX4d0l/7OROxk8aoT2eMawEGLIbfUGSmKsHCtNJb89CepTTcj2iJDuWRro3otqa3MudaVKy
hnOEmXS3MwF70TW06suRTzBKvZ8QdKnv2qpB6DuJMVeqUB58jOHyNueuZhdu7DavvaTWT3eEXpsd
nzMRKwG3KCh6iFX1vfGOawSXcxkxvMpDGIbmMz6Yz/bSAZT6EODZcVI8GcfTcs2kkllRmjygR0GL
gJE0NrutSahK8u8j2doSxW3GEmOwgWckAXWioI3KBIdiQ14cIPgVnfYmVdB5kY1gLRXdc1963NJc
LdmDXES7CA3jGhyK4c9JaenVqtjNWrGogPUcj9Xmi9np0+O7Bisy/ftXVv4QKN/Sn0tdG/e2fmuu
uXlH4XOdSzunKX2sOl8NuDDIV4xc1GBO7W+Bz/qcJT9Q3aRYtwoL0djxU8Tnw1Ef1pV1dgNURPhu
LguXrmbYWoVwrCi3RxtchpUVRY7NBu1JueuSMNxg0V3qdQXra+DiUVcIKH2FLvRRg7uL+Orn2IOl
Ia8GCh26GqqexdCo/qSROP+09HS7fiwSiGFizFVY6vTyrvvy3Gj1YC0MpLHIuVRB8fVFqsqlCYSL
A5FeEx+iHeLMFeI/r31Hhy/WfI7Ut38X6Wy17LEKMjQJZQ/hnR8u0exPGZOrDTicB/XA6cNyCYZk
sVnrNnjWdeVTNfEgleVbPBpQid8Xkfx9q1mCN+ovCb/71wYrQOVFEZn+dU14mt+ZoffeOTNNZ/i5
+P4qhA5+X4d9WMX2sMY2cpK0juKoWhAB5iw3OItHmWgHAbx7JGkoRxjPGfNmRMhWKOoftcD3g2XX
pPDulaXeAFQGlIaOJoh0MMrf49lPuTdbzASW/IyW8jeYwRnGjRinCy2ewk7aJXVO/SVkq5AhwHMl
MeJBuWP7sCLwhV7o0xiJQ/+MeTZCs7TyR5E2Kr+44nS/zV+Mqqb/pPiHy1D7S9hupNc+KxEL+We/
EoVGuspEd10jjDrrp2P65D52JSS61vxMRxuR2kjm+OwM0A/87bKRUIue1gXTYxwxu9pVvYQpvPE4
pVFq4IIRrSPLZi/iT+fHYppoCSTSe0FeLEvmFkLeqaFX5kKrIMjx7Te1M9QODpAw8TP+/ubWvfxH
PlE9jqgvsgE0GJ/lJgqlmnTWGOfEovWgsefVQulra8ELSbtN1NS8TAW4G+TKOGVqimvrtLVPqbbh
XqBp/MnfXrd62WLl8xgDXhrw3nYtR/kLDWfyw09v+yXOA9B7T6O1vt2A128q0ipcUdjd0HiN7B4o
TtFxYlWxHL8pzqgVM089KcwvrnPhplDlMc8BgNZZ/nmFw27NX6rESX7In2AGERUgrWtQ5cSMKx6p
yJBEGV1vvDiLihjj3A/VuYEE0VjnTMHRalpDS/YHMP522yjGuNzGfwpBR5aj3oRdJZN1oaEusYNw
NaWjlEvmEPdakoiF8964QQDkjMOlvR/4ld4YixjkLa0ELF0aqm4+/KFSpzQwdoVsJK4X6Kv1KShj
fCQ0hNWGXut3+P7166QXNNv/PH//SAWLGqORFnLfN9coTrZ4Jzoao/Qx7vdX7cuEWvB0LVlPwMnT
eGMheZqvXH8J7IbLzP0qCzVjtHDSKYhzuA/JdDFAz1N0mxk/PYgg4Si2KHsz69inQVrp8YdPPh7I
AnYY8CIwAaP7lfod1qEQ2oTWj9p+s6ZrTwwRJ0NQ7tX+ctcblBA1bYGmOTABVdJ0PtcDApN6wllY
etLEOXBdqgWSZipncZAjkuBVMtSPOLCfx4H4T+1SGHZfKc7YNrb7AyFoItJDGLGJg3SE4/2UZeaw
UEdJk5M2LKoKcUSCwXKIGZZySYoWufPn6g+TukItTYWhsZUOK1Vr/0xTYhBEGzCgPULt45Gd5HaD
wiwCRG36uaMbwwlcukbcKcus1Dsu1vf3seYE6OM67riVQiVXScffNxQG5wtRNPOxD7M5BLaDxB3s
Qe2KhGAncIJM6KvShJiPCKtjt17UojacGYsNkah08n4paafEbo99U1S8ZqX+Ze8JPnUu/Gi8D9N1
KlOizHHk8p0uMaP+J2dfZqwBv7nAL8jqYPnmtvdpVmvTRk31CmKDzvTNwKVhmXs7hC7J1hdll8pL
qk+9hjElSbJB5TONufZIlbDCDDMZLYMDcM5PIfkX3P2/udHkYOZpjmAoZTdA/G1G7/Ng6kjZVqOM
aZHKxYvC+TrAoKLMOoelskhP8+IhFa1LrLHWnEeo5PrtOUB+sgjWbpGCumusS87pN/vjJae3Jh8d
7AglMUGcUgWx5gDDVOmXhSzT7LkZVtdBvWHHIn8of2jqmr7PhGRi+weoWEJ99icEmIKNhXsfU5zB
g1lRaezTLYbJ12cKdWpBhxEZ4cO8qecfxCPrnTlmO+xoWNjZGqBNdq3lsV8h9lST0zVNUVFSBfC/
7P3ovCDgKM57/wRNw0aGNdPOWxeP51V9oCRNqQxvNvU5WGDVOJFQBnTcMWGTCLpq+yzaYsLqmcsA
nYBrVUbgWwPSq4HoecjAn7MVRJHuLNN75fyRFgnN98TPaLkDNIHS3YYYunRRMi3K3jKhKtyu54Jg
lCMbw8rymUOAYjyA8WXd0ir0wFNJ/BtOOB8/k3zcKXHX0BDV9wFGPTd7mkQc1R4P3VUgRL2ww6ro
onw4rOiZ0/5kD8ioVUlKz9pevro9oTMJQv+8SL4+EuzadsFJWqCKmRhaz+JIbZ4usV/1pdo7uaKX
tuuzp+bkDZo0lIzh7Saf1MZwZ5lk9p0xr5OAiS2tyUvK3Mudr+gOU2ZadqxH5fuyC55+YvbPlGqp
zTuRlJ/BY08hs70UsrpG5QYCC2AewLqfQCc/QCYDBo8qRbVsKclQGNyZXzE/SB99QwdfaOqifKs4
JuOGrdBcDrO3DcwwNK/DubVBoc6gFUssftXCJC/akBDmlUYfFA/iyndz/XNA/vEVjw0287PZ4cou
P2rfCgh/OS8b9aIc3ygrurzuuaOocrRSfaeT0DIN+BykIjUlmoztFokITISiPqsAnMj4btW+JqRW
cRbpTtQ/xq51rBDgHEx3fJ5ClSCdlbv75Ksaer9Se3BE8Q/0PCM66RLnwIc8k8WgMUae1Rtp7UnB
3x1V8Q2d9jy3u5D/SZSohNJN+jqTlyvRsHccIm3XVy9qaixv2Bnpo/56+qgy8/D5UYvDAqZUHZrO
e8As+42N3Kh+m1IE8e6BKyRLMNg/4Coke7jC0m9GD0s5LU1R5gRnQ7XyIX4Rm+eVC9jqiUMGYALy
ddBEaSk41cnOMlBQJjgdlvXVWUuXooULcmDGYT0SUxxftyrG3ZmsUj4eK1v5fev5luH4H0B6JZ5Q
WeJzkAovyAVrRZz9tghltePi2l39J6130CumPMkxgN6buZynKSxnk6VMoxuLraFIW7NgYU5Mj56p
dsXVvAbP+9AXUquXD2NRYCygddeoi1blo9a2yhMzl4bgm3beTnsrAsjv8bDVyxaHZDWUr3A52Bo/
MxAB48H2lgdUyoc8q8FayNcVX/9exqf0C/l/AcwKFPBB6szYeH9ggX2CQEQIcLGkioTJlLzu2HjY
lMLz8/7Pyqnpr+yjwZ0BJ004sqMHTP+AmzNtRV19yggSfCSAVbbKOiH5HOelol/AzVEPI/SGL1UG
QrSU6eq0QPXZiW1P3BSXou9CndQfhwouB4EZ+1FtLDAdDciY2zU0oHK0+dLDkHAoQyG7b8YQMm9P
OrUMPz8QBYg0MHegK2BMH6kS3KBNxKGtWQSLRsuNPcoy7vVgPGmCSMm4IqHR2l+MUqjk+JdiD0ES
59/rsx0Tok+vnVQXWozrXRzdpRT/tjisZIy9L1UKOWPuPHDBvyhDDig4hMwihPZBRjlq7fCK/DUj
8lP4MgWr/0yVZcFuwG9VzFyGi0Mp25R1CwL8PxL6VaUnK3JhFfNEfOrmykf6rDbWYx2DN1EFFYNs
UHkgmmqOeYsj7/pcIDMrm7tiCl+YmcYduT1bfuT83UD2shikKdLLoxX34B0F5dinay2g/68Ibmd4
Rq5jz9Vw5aUp28p6/ktLw3k+uo0Hps36jSp30zSlcdTxI1QNapZtW+RR/geL6qJ0+6kh/vyGFX0G
9i7qT+LKkLFvf0pWvLTM6MhKU0gFKJXOKCM3P6OFYar3GmT3JVodhnBKSF41DFZnWs6UFfQUCSqz
ZTHYyzA8GF6oK0st5zfUmaPRTo74l5La9ul/bj3YVU5jA1StGthLIome8X8oPZisV3+AszbhaJfH
+H4xRGU/Tz45t5NfAZ7NRdbyhFQ8kt4qaXcjPCm31cT2QBuVaxoLmcz5+oAa/Ek+1KA3E43CjAAZ
cZYFtvbZ4gOYDi/7mDGJmmgqa9p3AxT0kfGc61ELLM0viDjcRmA9rLSMULfUZpfM5y9lXXXyhOOe
+yRzIpfp2fsJrD6KZ39R/AiJcObt2oRFX57oq3C6xgFAJHHAd5yNnBAD6Vy7NzGCXtf9ZkD3dSIX
yIxN13rgv4Gm4HPaHZzrcmSR6r+9QcGU5ORLGb0QWXStGF4S+HM07NVsYho2bmzo1yM+uT34KE3d
GxqMRgbRSqrSXzKA1cx2H9iV0AUYb1s3Dglb8rmeI0lz3DS+y/gEVtQBpiPvk6CrYYsIq3aV6tW6
IPt3W0sGBhHwI56ARlpQftezMAq9GJu8+e7+Bo/AHiZbXT/xb8qVoCVo2Qj6TWYnk9YZocGhePjr
pS+09DEEfqmyUPq36hEGAXRzDXT/50pE6guW/UdqiSgTaatj30sWlpsZiW/Av/GjliGwoQYZCDj1
jx+UBLcdUOzzJpHsXyITCl+GUFbERr1769C6ui00lwBUKzDdzpjQ6j+BIwa3o1IGKw02OSBZ3m/n
VzZXpc8PVcuny7v+L5Q9Tl39+t2aENqPEue1pUObww1Je6Fzma/7bLs910R1MzOPI+fzAA7t1/UQ
kJ8kYTfY2xREosr+13SN3z+kPGVH/HX5SIywiMw+QvWw6+XPfjbfhXDE78xpWgnIaOTijvuT868n
ckgLXudHZ6Lla+I7hbFhJr8fKICUoFYgEREqfxwC+umZLqbfHoeSbMd41fQncYAGROaVO9XAX8fr
tgrukHAe5Dj+qp1p484WfNc5rhFqOmLalZVb3CKorSV3aCJnEcanEvJAd88W+y9t/fgUU17wfl+Y
/fqXxCifoaFZ40wuARmDxen9i0aYztYVTgR9264pisgTJ9b06rGi6wJqeFsw0yEdWAYeVamJuOhq
QR+uhm7FY/9NEEXGml9Qck9zY2KABgdnVRtIiWDQOhaRESdcHJiIN0KFs4uDpNrN5q64RZ2dL9bk
GHP2bj9tAmT3BbxvCpm3hInzJ3LlbYRfcWuOSwaJ0lCVuth1Tb1KPyFZUzMo22CxPUf4pGXg3j6e
DAZkkXmePKXnmSs2yBGTHeuzivc2BWbt2hAIN+NeoOuh/zXSF+9c1AMboTrUEpwMJq2ovXzzhdPz
qWDkXdy+kXYX1oHXaECciDs4F1MjEf9t087iMjZdS+FptIkjlI8giyC3sNVf8doeLUu9fLBwQatu
EoJcI9hudJ3JGVJTYmgBSK6djpyjs5tYZuMCHqHEG9GTJAJN4LIQMzqQKGiAXbL5FtQvN9phIYBw
0/6imKXnIB5LJzZWhzmcNfKcDb5rzXWfE9FebTiMVMqcUzaW+hNDYbXWmYTEMOiB/pyDgFafqmMS
i+NaQP+abHkfShaBOPlCZ6vjz0JUWzQn7NAr81MseZzNOwi0DfuQKV7ESgyjh6UM2phtNznylV9/
e0r4iaKB5FWbJ74nyc42h045YD2HR15Ikv7IQqCqbgHqAanHRhJMYi2VmkCT7w08m38ieNXyBeeg
vGpVRWCVOf0WDok8vdQxPIIx7ui9ASgoY4L1AM6s4VLBQvIq5soY3bi2W/jiPZ4p4a92E7ObHNpI
mSpbYZ1Ioj8PtkNnc+ReJT80EX6P3utfhLOcek+JiOSe+HUzaBUpmooPH2J01nRvEaixaFeqIe5Q
mppgN+kqiU9JAz3O3+EjPSgHdCdeCiZuTAt+ZZgQNtb/UcgM9/f5nvCKvRa8EPY071+KIlQhiTPl
HghCZEtGi+2+oKn6LmAVbYIMkNaegT/hi6ZAv36jaM475HA+3KlQmLhxalYgtxplqwgiXJz2PiYe
aJfEKLqfFkxm2YB4vXnneRprSTRg5U9l6dhOckPoKISFJdoey2f0bEMhpT0E50Dma+yznK/6oSKX
GEbNONB6SZ+QfXRsVQFsSTWX5ErdpU49R4Kw/W+EpxLSkNfuBxV8Ds/QOw/ZUGj2mnXxhvRkonDg
ZNmXs+Eqs6s/cwa02aLcEwcp9GjLzRGJAcKU2LA4bc07562qx0Zr623D2drqMaeyFmFEnMZs22cY
pnqHn+4DMZPAtGnU4xdWmLfgNIgu7H40KwTMtm755J4FY5KjFb+KHi1lMwGBc4Nkz+RVU1dbaUHe
0hrWgnrz9KuZcM1fTi0r80NiOsXl7CA2f3Atw7yjt3AFwvJ1EGPrKSdZL8OGI8iI/jDd7FJZkEj4
Nv45msHWNi8PUAnrmAWsSUsVh6ry/eigHyk4oUC48zSiNq/Su3P9UzrVJSLC6YkwGU306NfadG59
3R4RGz8fatDjJooM5Wp9KC8MxONU7QACSj1a5YiCpLuVLQP7hRBnqLPgSqWjHm12bKe885aAlIIJ
0zmgUKQH/LlwHEpJCmPPdy54qKC58A41z0+A1AYY5XQjw/QIH86HcpIy3DLot11qkO7r2y0n9yDQ
lZG/y8A+2zwqtROJCMS0wfVUdwLM3pZJCKf4lQz+GsclqD4UBm1TQqinSp+K7VyA0+K3MtTfZg00
3WI6rGMmtIvVkinoDpvKm7/qB1O9ySR7BjDKAYo+z9krEv+54wCMQATjHauXH1xsrfa4AYw3gqDA
q9q8Q6agbqZmv+OoORzi7a3+LwWBYFgFUIICScHPP4fppI4+67pTPvW5p/k4XJFuZHLDm3tF5UIW
kUWkwzFi0t7K+Y8UDdq9ck8tqHw3rthVHDVciBRcJBlUAAK3wa4H0J7O+Cw8yftbyRye9iuNzU0+
NVgfFAG5a0x8/bYzCQGEp/gIzxHU96Phi74kJnh5oEkn2hIOXEYxiZ5t2DHGzhUsGIz/C8ZDMFp/
C/ZJZ5HfezLZcGKhu8T8yQgrCGiqzvaCQrwsFljidvvaTI7GgRtoj2OBM+Mnol1K0WoUo98mW4Q7
ifOeWz3PE0l+dg3CNPbGEXqCcHgDICx5QLYByC5xotuh5KP9RbJ2p+gf7LZ85UCzFdw3Mvd+kgiy
MD9dS2q1QKur8dNUJeA+finp3mfw/jkkPD1t3/qXcRhsZ9rv0ousBh1gtF0E2rM9WpSzW3pJuE0F
8WJoDv85Hcj/XqVrd+CIHMdNca4pOrpeue2A2GNkjD/CYMLy1VQ6nGH193k3po8+CQEGVk0C8+aW
f87DDgHz5FQ3mzutNnQHJE0kqtk8Fies4AyObZ1L2XYumgLNytVOXGdooQHSyK9w6Al7V7N7Ue2z
SU+ZVifk+50d4TSjmBYrWCWr9QcNI+k1R972GBY8rLZsKtXW5BIi6MmgyPFfqlrYVQViGkU2ql/T
TWd6EQ9Sa3Y60kzgEBnAuy/buBWFFvQWL/mxVeuUfq6R5CC2FKyi9cJNRh/Iy0z25qFVQbhWT/TA
VRgQzbMdZ2KYaaWhPruhwCf9MBNvMwuYR4Kia2DGWUscJUxxGF0A1x5CsdPybqczTFYBX2ADVFJp
Lhv9u68b6mnnhtYaxcNBu+6ZVtWmqa5BwxzWTqnUN/vlz4EadVvHX/kO0QpFcVVLP9XwjL+xtMDf
73eYF4zg1TpMYZVhs+X5W+JDRkqf8rMTR5o/YmUc1aJsvi1xsDQgd4kXw2E3Cds1lhKhDvcF4TWa
xWWWJ1vRj8WcwUvPtFy6EjUFrUOgcOGALR49p+pZilzgsfYiGgqV7bCht95cyKyo0JqGwREBLYHI
enxtBGDNrVOGKv7yf3dcYHpkUvFYjzhPkMuM6oJp7K6VO570zYmoVja2vt+/XZ7Z7cz1xV0ALRID
iFkkjhNYsZo5xZtJPALHf3ytKFSaeC/n2ydqH4MQ6pyxcSIRlgRdLzl/7yRgM2W6Lxlt/TexfBqH
RhBCHfuCAcKjpGSRZMvJoVs561ByturEdYxCRbLSszmPVJhm6yJcG/6YHeWTVt99SYHH9Uy679u+
/zV+2o3G1fDGJ+4UiUBOPuP4aCb1J3Xy3NzHgSNljcWTDNniL8//7nTyWkqQBUWvVN9ilzEEX512
AmZsYk5zSfmkJvTIgld0+0417CF/FKcOkBX0PMY9Y9awbHOUw9L1GsWMIbn+QZHvvWzFp+1MATWj
TJPWJmJanNefb+yu9PPp/GN+w1hUrjmzIGj/LhDMkEdFkl+9XjH37TuGbSjcUDBXajugN/sxdKOf
vYzRwh0wxCLihvophiCGpbRpjADGru6NQtqFVKP1W6KtB/bcOdCLyrGBMkh1Lsv8JRNvVtOMZdSH
1vaSklQ1H6v0e2U2oNCSnGELRdtBXL/PZ1BxadsHdJysC3Jle3BUI06c9ffnciMmBhkoTXUAxBOX
hsqGxzt1aXfuc6ZRILiOjFS3X1LFS24t8zlGjusdC1JWm0xVb8ERN0OzxnB+xNEysC+cviM1GSVL
WWkq03+nzhXXaLokJ67RvCVXavWgjEXmXNnp+jgV9uyugKEghnux8XGo65ZD5av9WqW6Of2l4Vko
UL0vxguUjLCccXTrv6rwZakXTztLbLVN0HHHmHzDXDsH2+cnsAfgqO9ipuN4iOCkMEueIveBrD/P
CeZtb+Y/HqFANUdKK2+HNO+s2T4jKGIsgxYE0GdNpSrl9F5pZ6pclkZ+0KszuU8WVCD1U+9rC6E/
AFMi0rXTELwCzH3dHB59L/ZWmguPb4UeneSLTGkyk5TVHkw9IFHAAiG3YH0bF9X0LXpev3BhXmCi
tczR77oKqh35jZwnOgeUoXzIEUap5c9Noebvr+k0dONZYCs4dEwiXpQ5oRhevRoRwawUIVYSFZUr
1ZdwCJAOBjE2yhwBRu/Z5l8eOlrM6GS07o7wpD63bFrXw1mF7yC90XcGgu5AIqdTRcyELuXMplxp
k2KVV52mGGGmHRg9Dr6Af9+EILH0SNUmmwiM1grrNwVlE7wGWCv7zH/gI4Xl9fw09DsGdRONiwuc
gOVo1Yu44DjshhkJ0o931K5OWFZqxXdfQOCzTDUYBhCLQsFT05HQ0Oyxhvd4wvao/rhQ8e0+MTe5
+YUMGH0XMhc2860LjhC4kQvuf5Tl3O7v1lld2kEYhr+BQKsmmGI2hfQT9F9YIrM9OvQfg+Vo7bjb
VAGgYWbec5Uc+UxVrk8mZuSxIChYJ/hX7+aJhPVnBIInJqScCnuS8YhglO9IzmGSMOli1BFK9PuV
WzpFTAJGkJYaUq30mH9naF0yTQqDfIEdls9c2dH3YLxfIhHegdb/rGGAhmpl6+HFKYe4PvDXePA+
37gyt9Dfb3W06jn63ZUoLBXOVrE8O2ZedHOM4HoQr1z49EZUxGsMhMTcqWRzEglpqA+BbvPVT2sZ
8DpyiLeNs5202Rzj3mB5a5dOx8Di5GU2tSZyE8JVS9lW0Wu2bj44Q8EE7tSzMpwNRbvij/7e9yZZ
OSzzeSynvm4thky5oindqxf/k3AY7xRZL4qQjninPTQ95uhNE7l2NcF5yqoj3Ly5Gl/jO/JWpc9P
3MsDVrN1txpC3phniqCatHNPtNIzIDzZxblwtBbKOmnHza9z0UsH50EgGZ3kI2QAjBj89RXWYNKG
z89TaOEOuuMx2o76eTbPz8UUb67+gGHMJpGly8YH7i/r1+YmP3/LwptnJJ838eYjxUgQwNBPTf/Z
fmFcdpcOboCuWBIWNoGn0s2p4mFsqzHqanwicTaTkFqdWPvxkCPZSybYpNn1gSrayy1gCsXgoz7T
ovQt/NOpcvasELz/rgpubGkfVP1k3Oe6MYnnp8SmADMxj9+/Cn61bIbWLtb5ufBtJaDtWKTWnzJ8
WoGVUb7BOKIENsA1wtvtXwVsAGUomzcsIBSRiq6PiuPfBA3//nIXx4f3s5r4ktjNPK78wsGi8nat
ou/foerNpjaoUYaWdrkJFmWKATb9ABEGihUzZrWZOcB4fUE6FAIzmiUoDpyhfgGb3ywustLUncHE
xn7EBGxGcRPodIiiVQIejbm2eqxwtRl7nn/cf4k+mJ36YHSoOpROsb5ha0zwn+XeA/bUrTx+yv5s
w7aqVrQCQyFOVlTaiTONsNf2r1f89jHVwOYUdsJhCqpX3LnEYQjBgC0EK/HzyMSuuP6/+FxrXVWv
QXGn4ZEGzJBj9DJROjoW9RmCyvV2ZRU5E4qGhr9hGjzX9Td0Nil5ZLhdl9XasYq1ltHf4EsZh1//
L9GB7Qt5O+M/YCE5Dbs+s7aXORugYaBy/CTHFfkosHlvM3I/CCjvCq5WiJEK8EW6G+ml7XSZpI73
FHs7xrSae7fEtRTNpJeRPZU0V9z5S2d33JWQZ0F+3uRk5jYNu2yHklKQ1ZgBD7aUBqsAd1t+CbmO
jxHxDHmPxd8kBHVYyMZYAWfihay0Kb1a/5XBIRrV5vfl/MUzuUVIP3VSSQT6+c6kkhYJACsjag6B
4bCIiK18MP2a6pUFifzrrRKB40W3ENEy3zUaeOsrdtS4C/ix5gOLUCeDmw/a60CfIHxipVIYUbAG
gYfe697tUMq5NpdaOoMLRBzdoBSj6OQ8ui8tyHUg8CqtDpDwycFO23MPJchnSZZNJyIeysr2aCcN
lXCFVmNzDHwtWsI8M6awJBQtpfwRyUEYlknV+PHaxZlJ2EKhcm+7+ePW+AjZT4Ze1dOUBSL21Cjk
ScFhZTMA1t2VLAFO8+ZAv1ecpqRtvey4OzesYNUop7ebzMTLnv8mFXIvpEAoFgYV/Y/06l+G0zaw
qd4h/CuHHDqkNAMVPPeTxcL6P7wCFca+24I47P3/gAbtybIhAkrdVzgmfWOmVAvZp1KWD+32SSiz
l04Z+sc+0t24Jt08u5yfVM9cI724wdMWkm4L11fhHEu2UDCPbI0pHlNCCmii8GF44r5ikuyvvdLa
jM3e7VXCWFviUPiSSKufDw3PNrL9lBmmsQIJjoEBpYTIDGblQSDR8+r6cbZBIjrUzlPTRnwyJJd/
fzz+UmVwY4YKGSJ6FrXqpOvfS4+zk08GAuu/WA7GGCiHf/9cq/kUvG0RIYj6OGf2V/OVfgjQcsON
PwU0VHPUs4XoWUNrVD/AjZtvr2xc3xClTZmnNhpEesAEyQ6HCJ1XoqI8h5Ie+UoTsyRO3JQ6/5uc
NnR68/63RXtpH+i1WJ9LZxLlrnZN01+Lry89iR5eWa0b7V+IWzeoRRvi+2FwicYYamPXIpSMhtw9
AQeL4Cuu9qies59V75PpWJFL/5mPAD2B3BVm9JHqHdBgL5PfcWQDZ6d/asug1KGCwV9ViVtv0Ms5
TWdly3Bqts5+OS1pH17iO1F9zopAEoJmuTjp0jnzQWc55KWYWerjNlBFp0hlQtw0LeeBadPEhXHf
ZfEYC3qI0AVUE/N5JFbyuDb9XcDmmXLimMFtYkAQJ8BgXj9CgS462NeeBK6YUdCUjhpXvAGzoDmz
gRcD3gTQAvk4J1fiDNBcM3fkJdCNzWIlxYuAJk54rvaVlO2IqrQ3lcg7nf0FN8jEiz2DsMmfVUmo
VNvOTHHkyFrLu1cmpPZPnZQ+ZIvr0IFxZcH8d6Yc2sCDNWEoRFLWD1YdyyJM0GHWcfeeBgOddRSM
Lq7UWq7Kr2jGvhN6x4EPxBiR32NfzVIjtsT3/67ZtSa8vbxBOd0Iso1RlXMVMybTDnZ6ZOAK4+s8
Vb/SYVdjPUnK2dVvGY6rbWC+W+7EQFMuRSk30S9cIMpGc8TTPJszWh3MxWoOH/Eue0BlxrOzY0V2
2b4pV0IQcKmi2Fhgx0rLeGXZBwsyE1v6yLfNK7+mTXhACn3zgtl6J7Zis+ROSzn0SdpC1M4mxKoo
Ll1fmpXXGpKgdVAs71qOv+0q1uP/oDwCu8GyyB+gvkQb1JL3aHIPkX52rVlvZKIMRuayxFYjZlOm
u7LhMDZkKgwRavNFS3udfmKLwYvkZlsmOCqS0t0oDzKTS3f+Malk6+7FjYDu+/rMLMmBbVvOfGf4
mQkU6dMaE/pyBr8zNCSq4xJ71LH5SFSOWHccpadjYJUmLG5j2u7n0iZJCRj8og7BoSLGeQh+lqNI
/eTiaVKKIJrb4Oe31wNUMJKw3hKwLhrSUNtgga1f3EPLL9ZcZdj3TH21A0JUonhO+pFW85H9VPj/
OVVtR9ge4hndoZgZ+AeG184Ome680MCdGMkkO/q6QkIJg9WHPDSUJmqGKT65WC9DIDM09GHIyj9B
6vtL4flf0Trlzvtcq/1CdaDeucCGhgEDAFVrbqyLdSVdT2SZovSp6cOvgXzJXjdBLue8CaIq3Bir
AAverAEMy/3mB7SivoEWfkeNii7MCC3+Nlt6kYJqBblJyvMfRp3y/O5PQM/4vSKBcM9m59zl4FMk
wzNK0jAZXaw2cr0xOc2+olbkVCsMPk1dGatgib3gfO5g40b0pANSCHxxKeHGsuen0gnu64FBWiv3
ZaUfLJHSidLRTirfOYidzHiYCMHlEOyf/Bs2HB4hFPqUkIz4/uMRWzHl7EfCQU5a/kFscjPyoeAU
QG3OlSyipUx1+Byjw0KfuBYv3zkwSx0lmaGY6jj2EUF1PuSenC+2sIMikchpaKDSV/TO3UzsKzlO
ldzyNQdCEzHpDJLOT0mybwsxHaOP6NwubN6jLyPG2GWAVxCafJ2y9yf25bu5Z34BtOgl4w2nXdkS
WEyixgfCOEPvc21HIWZW87d0ZIzT+tGT0phWY/YC/7CeZFme/g6qAk6jyCaEPu8BFJ5Cw5P7wFJJ
FKcKgvyNwLYpS11Ll0HjYyQXQEoKc39iZCiWU6s0JkqxctNMGaaw8ehPGEuO9DJlYd7oiPE5hcfF
b1kQOoOBCmDavqsdWsZZm8ktKeHb1/t3SWUXonCmSn2bAqWcFFcWBHuaBenr5Nj6tQhkrEB2/1g3
j0uMxp6neOMYHvIOJmjPVTEfSVlUqFm8hRrZ0ck23Gf8CH0kifOPWiyCK0mIccuPG6iPgp8SApNP
HakzbbJ9qQOI299o+XV7xEgohnD1tmT4nqm2Qr4JQxYcTSBO2HqTmyvAIq6fPBfRutdTzU7GHNOq
o9MU08/juwPyadmFwfstPOTMGBF/k1RkKyKHBSaKlFww6XPM7HehUX4QXr+MgAhUy9Nl01XHAnTJ
IKbMPE1tj2PJ6ZtSeIklKic0EWoHq+L9tweyBnX4TQ1tXHsKuzRJaaHBrn7S9BH2iGc61my1H9K/
xfSL1tjFlvnLP7pxLQusg63vyLHMIrbN/lxdtIdj4/wufXVCIg5Vgr8Cywq6h9vySP5Y65gzK/wh
ZAGQrqOEL6M6Jjab/CIfSRZCr5h5Ed/lW4EaQEkxovlAGoo2a655CYPYyc8gY6ftRO5I6XKb6PzL
iDrbBfp6+zuSjv/xsz6zxWPzfx7veKfgX186eMFangYyw9BI1ibhGIIumvFtqHi44x+PM5VLfvD4
26z/aJqz9bSA10fxBPIjV3FM6gQ97ruCIwS6J8lE1iyKGDguQn1deHdLl5Odd5zJ+4FDQ7sTCR4b
zVWyDHJPTJgDGnLOanQ4yyrrvI4HsNPA/Sn9ySbpEcavjNfvUNdCZ0vVb1qiSS4Tqusb0pH7bkuE
Oes5enJto/G68BlrcpJjOHlbWbB7D4URCRMFgG7ZYLYlYT/r5rTUE/meDYnhJXXCew8WxQahNJBh
kmX/PzZ5Zl2ekwHdCnns+gcDrC2Kc7iax1NJHmTzwPQuWOT0tkJCUzR6f8QgvvjUjZ13LYD7XECZ
gUF3Gdw3ALtJSVXwI1Vgvz5kI2HlDqwxMS0e4YlzVE3VCsu1rnT0G2QJYH63v+y+Gt/KRbwt7X32
FZNACW6A2qZ9kUoBuy9S7pIF/DdnMWJ5i+nQ3nhiuydTasN67wLBOxFxYpWJxWEPbptBkgziXU4u
DhWO8rH80BeHcwFj1zEMu53E8LYWf8r6Db5raRBBkJ4mHBpuGckKkyzLzuJHj4ndli2TwLLlDg6M
cWfLQuiN7dyah5tSyA5Yi+RPrUKgkY+do01rCEAqKnUFYtz61EepYn5N/4Ke5u0DxyDxW/TeeOzD
qOWmFLrNdSw9iVK/H2g6li6A7CMZvwzUxQJt0h/oadG64gB1WS48Vy8O8IU8CR79BWedLeoffp1H
m/FkE4xNxAopm1VrbRWoJXCUr+Ygj9vYR1OcR146U5sQ6NI8+jrgaKjUWJUQfqMwdN55eWS8ylZ2
F0dpO7ziB/NvkRKHUxgfxbjQ9glJ+uKHrCWF1rd1WfYJvni6/5IrHxp5rdP3dokF4xPSowVB9gHK
OSTpsnLR81zmxIvpigQJAmgz35qeI3fgBg+MQGoxLUZZLdZv83LpexShJFj6ed+cO5CzsLHXeYxU
qdRBDLRW/r0/g2K5+OFdlAZcLCPTNunw7M2RaDk7vUuVVQCnVevNrLK2nRzDWbDaERdgdcyMKoA0
gXgpLf/Imw/bNlFE08yYg88zcvPbl8Pt+BBG8MoeuPv6oYu9F1W2ACW8r2kWKdM2zIYtaSwmtMMQ
SKiZ0VH2kqS50K78Q9oxh7VLKJck1K9iWoj21ulYIJv8nQDQh5UTaxzsi9/7FtkYJTlgeOtygwcU
U5oUGAU4zx7gXLHSkHQOTIP47H4H7KuLBU0O07lsDV1DfB4WQeE3b4Qlr57GxAx/xQsFU6fnFwSd
daB43Gle8u8M7xdQ4Ul6uPuVM1gSqUwn3zxfu7amyNpZVYqypC9VNMotjmfO4zepLnA4vFBlau/O
tUUdKSjJ8PV0y1GOTHMbGuMa1RdhEvhCrFD/Maa3G6noZbXInzh385DjZ9L5AKyi7vdpTCxdSfbj
AS9qX86vznLPzbvPYlAbqpWdoVqkq6/2iUFVnRuyt32wsLT+0o/+vkQFzmnJmHVGOqp6dw45OZ2g
0SfNQU6dEww8d2rX6shRxG7uuFV6ivhTg8Zhz/tpbtrWtguGyzhIu77a/JmC6cx0/ZXjgz9lWNOD
BF2XPqgr0g9l8hahkuKdLaFZcXO5SvBAVHQ+QDqY4VfDKoGjN82ahaYKk/Gfmk6jTYAgewMVZUWA
soJtBV2t364O0FC3RgQcFfdjCMLOlTki+ImjWrZgBt++C/zaBD/N12RipEXRJLLpOCfg0yqzSi56
oO0H/h3DLmzy7epy4ekIOj48Szfs0jFYL3HGY0HCaD2nxxFDHTzuGnJjjuDDsQWQf1yxPt2ApB3d
jl34ka6hkHqS395Xxo5HgIo1DNTckgQT7PADjd1kgEP3//0Mzd887sgcWVme4r1lxcLqUgkqbH5U
hAz178yWGkSAR/R3ddTDUvaRwsuyI+biqDaVjqxuwHUuWkoAlsZZ1kR9QHxiWPcY4HwLuJR29gAK
o3DHKQy3btEG0NwH0+4Cw6E2KO3rzRcpI0+/z3tpXJjWES0MSXaPyWRaNLdNifS64jClhxGSg8Iy
bWhcxxbyodBxxNc7n3RJgj1SNLmBLJBFoif7a5cOscwLkFtccxkTs6F3p5vRmIbzYtQdZX69Z52N
o3DlKrZ2Vv8bRQ2ohonWEQCyJZzdHW39R6+/tgl61tYG1J1YHkPHwUzf72tmbu5EK+kJYaHcGiwU
eatAn5K6ubDU2tI1Gz1X9I8M0CgijiFwZaHkvONFRnPzElKbdZyNQ+dski4zBwW3U/zr9amznQnd
chkypefDU7/KAw9gXADCxFua/TGQraqB+ERXL2Q1jRz9+89f6RrIc1/SCbfTrhGFWA8DITs8Y7N3
d3tvPmxOFiFLnB9ob6TzWU8XhbrLEkk0+nq05sY+4qOe2EGHZkze6oMUj4tQYH2bNZwKSQATS2vk
I5PD5hLLjKE/uozrI8l8DRTZ1zPQMswJYtcY3Kc8UoDfRntuA0ZcAb+PzB6T818j4UPdMCLRzKr8
/+fOPxxxAZxA2exFeP/5qJ2KNA1JpqE6gvVLKEUSOAjrP6XOsdPprVtdXVw4ZAayaHyhOLP0oEJ2
79Y1yk78nq+0lNEbAApiJ3JC05UbxmMhQsAB5YJ/RXABWEfHJCq3OQdj0X70HNemq2IkPrKUIWM4
VetXN7MknCXLKAc0rrW28kOwEc17k0zF22f6OYd/NCoT9ytRKQD1s4//L+V9BAopUcYilkpKzXBb
aE9DD/G7+LbWOFF6rw/mCU7nk/Bg+vxFUfyBH0mVO1u46x31pCYSJP1xIX/UBe0lLug/TfLIkEYu
pU3/PuqjK1C6hagiWyGqrm2GmTtKPyy5TjZBV4X0kezHe9rFj/KkIjVGZWvWAPHJ+Irw5CkPGnO8
kP2UD77AKHGP59RJ1O7s79sZvaPFolnHd5AF/f4+THgu3MZYCQyEVlVnaVGXjFhHVY3JLDAjdGbn
JnPWv9IBcJjDzByEBtWdsqbRSEaEsRQcp5jZcmGIxvu4vCmwoxUqwevKWrtNt4AGax8NYOy7ztbL
f4/kPloKELgNAcjoI7pa8OY+hYJwg+GbssrObYrZ8/05EGDpYKilhccRP+kX1tzoKN1qenu+EoT4
LofAnwzwGLa0MwoG6D1GD/txOmDYsXXgF/dakSmqojwzIu1QksSZnj2Kdo0hS6HM8+IBvE67+aro
3mrV5Q3EdIa4Nghj+pBjBDjlwHOaaRMP9dOV17XVvwr5thNdWrXVYFzBS7DSCQULX0ws+MdXMy0I
bxcOEr7lSKjL/szX5/XeLknV+nnMXYREzjsQKY2RA0ce4+3ocDKg7S3Q7bUCbfZTR5O+j5yEZYz3
FaSZ1MwqHtVST6FrjuD0pdTI9OLGLYskSf53RLGukHWldFr3Y/oTbJvUQ+WaAqHPUqs4UvvyMddM
eTsPq7xdxk45LHnYQ+moDEbNiH02jaylXrw1EsjJztZck7N+y0yJRpIP08dU0+1VOYPJEM+qn4va
Q4nDfJqvEwAD9Kd8j90+UjFOMIv3TY8bpgIaX6aX3d6IosrQxhHYo7QieMRDivApkBPEtkDm/PKq
ox7s/hjVkjGK98aCcNSltltqMM/3sjoDqbypw30Hx3Rgk8u0LpDVlhcKWIcny7cyIS/h0nvNsZ/T
FBX1p8jvd5eOFvW52VNanL7iLLIZJtbpNS2VfmI9EdEkNMBHMQLmTV+cBLWBATpVDJpAiuylRvI6
TWIsQMitLrPeUMTH3TmTddfSMnLyDaH2lO6P+c+Ckkp2CkGcXZGp9f4KwTda+Z31aNR5cdxyYm2w
QBGTrKV1r81I8zgfO+hiu6TYQ8zFcuz08oSUonHrSyQz5Th4DI3QXAQC+P/4r2yqDYfIF6KzP1/d
5C78kbirMU4buP0hhQ1BCRjiKWxHbK0qbqfeIGy5Chao4jNvfPgnJZpoLU6C9PoQDwm3G+e4mzhy
3VIq1RXffvwFh/iaSgzPNwTUH5af5Q5viEOavCOR3n519v57KYxUw6oNmx2WxBb2nNBzKhzgRrYQ
WiL4ifN9kvYrMEF0a6XfjfXlVQ6//08pkxed+JDx3Zmf3FRXEXK2LFTCVAPJvE/wSG0/Ko0qMhsT
GbPNFhdfOF2owqpfvIFx4e7YepaqOrf81pkqUwcGOu7JWbUl1zCG3m206Ry63TgJhFcac9uis9tu
l2I1rHqAP934B+ECvg6hqF4nW90TvY4C9gY5E4PJINoFyXQHXysyE7I9Xwxy0itb2N7PlhDmRUL/
JH8cPDinw9UYL1OzrUUqXyiue+wgsUXuA3fNiJ3/upVy4rMuzbO3oNq8J0d5b8Azypjp03mhxQgc
rxf9iwcHDp5fTvIuUVwlWK6l2tz6H5V2OZerpB16tWnjx+OQJ/MagbyRuG4E8jda9CKGolONtp0S
gZt1yruwStpOgexsKwH7FdaXmFCQ3xPUD3LMzoak76bQ469yK4fHDqsLy4QOC+oaTKGdI2fDjs2P
Tr0KjvBIgedZSe/JUAtrlaDGsurcJRnYTb84auwfjyFL8fn6rFplMxOYXUOL3akTA3FSzof4mf+H
+u3dZhIBc1KP2mcVkLhePYJtFtC+5R4PUm9l+wGYdjcnMhms7D1RRskq4azCdaeGmIoVJwhZ7x9l
csoW/tI4VX/tRYBg0K0NMuQDehk9jcLYE5suLtpSDubrJUFhfexPzVdjmX/3ce6Qvv8uM1s5Hkvn
wV+0lA8DSww4+LvqYLOblDIUHaCPv302yowo0waakpY5Z6Td3OEPZ9eBCCwcHUX1ZTuXoB1uBkTG
WrNqi5SrsxUrI6apKPqDAuJWYc97+RKdIf+VXDfhF+W7c+ZukSMAeG/clkReFTDxkUdWF4hZrI5F
+/VPVtU/0NC2ASRIRZhjRy4VcDyge/uXA2vbJKtapP2jOnXbIMNW1lDbDYAAOmUR+3VZe6CQp8L0
n8G8dqz5GkDHQBQ9yzbYY4A6TZGVPZDddxjjB06Q1UJ4K5uyj2vRURa8KB5Ybh4t+x6qgwVVfxYP
adkq0Gn0AKH2AkK0TazXvhxmdZXkgXOCxo3k6NAWexNk++zgC0quIVTR9thWGntDVHB6xYYLVONX
xUG8iaAcuWrNsRcEjdyNzJqqiulGsY32/f2lYXc1v/LM8gJ2RtUNb+PFDv0WBC6prYuiGi0SMyjr
uAbR3FX+lWtcsQLAEND6Vxqg/LR+P/rcP1JCvTluU6sxXsjprV0IhmU0O6yojClLxw1ywJIbM99u
DS7UodSXQaHjRs0TJYVkA5CDbCkTrXt3xRu9IFmVTE4nvYgPmCZQAMU9eFAjCdosR/JYzDlYeLzB
UrbdN7Nyuqz7ZJjiM7mDvk1JIAS+A6Pc7KyOHGX/qA2CeoSG2msrJRhhLvbsWu8D/6E5pdXJcg4e
WfnFShgCbRl/CxBE95xlp6UVUS4L3RrCA/A3rwYvpTU+nY6SEczcPv63NaBjKiidaZkU29lzC617
rPsC14YUZgNW6ARnco5LEklKgKrJoBv0ocFoVjHJlNOnIakRZT2ErNxszV3Q8uY3b3JGco10noPJ
sFo0dc7wlVWJVxUry7FZ+6zhvXmEfBcgAJ444yu1w9L/6SX7vaNnK+6OwT+Ug5QAQlxL/jNPFCdA
WVuU4Xe22hJpOoGQ7wX3A3Lkhh6wrTs8zqJSeTFuhJ7pOgLLSTTA3WnSDmiMJtJtBRwp/R2KVIVq
ifbidTRcJabwRneYKPBH1ok3AyHxeSvRDkEngOR9s+YL4pt8UdzLGpeeHjjDUfbd5/JHzWwPfC4z
Z0Wvl05wXEe5oEOtChICLysweVRDpO5uLjzHw8OMXNdDHvboHv0R9C3BsHPwyrFPZGc4QlWhdVhw
yH6VB9Dt+P3y24sMaNklPFAWncKwSqMgi5wFrWc3IB4zllxCW56BHniEE5iFLA/wBR/nxwXa6SxQ
ZZNlc0XZxHgLuZGOhAjM/eRJGG+hhYKC/N7Rhbw4mCfqu5V3TpFlafrVZD2XkMk6C6apKTOs6asA
tTaTgP3cxzDlIroHsEivqWO4sMvZu2T+kPmsKxVdj6UEH86S1gtySKCUMg9Ne5mwyRq45MUcVYSy
/Uw3PSmZpby7Sv+gxusNGguTJfB3Wn85++zB75ZBprJlB22zJRpYM0yfufFVuzyuM4WxRY0q5eR/
MzMFq0dEZL1BIQ8fOyZ0mXwntT+Xu87zGHExgu2kOEzOslndbjxIhLwvxC1s6YLIMAo456QBEpB/
QG4Fj6fclyThIE8ZrlSVjuFOfNvbf+TYx8PupttfAT3kxETxVAW9nIs+SVauviyll0cj58ru4vGN
m3iamTRyM9T9pSM0fK28z9ZER8bvQu6k7a03a/gSqE/TSgQpJnCWp9VmCWqV3/A+176AKfKFX8di
mGBlDOiY9X1pQFakzomvAeP01ezcN/EHCjpiFNg2rLTB6IyQLkH0qHYn1nPX0qXpeJs4VazVt26a
9bxMN+I7tDeY58pkKijPFjfv4QvwB7aZao8D2aibqy1MFwkA7hKe2+0XaIZ0WVe0qcACcD2k+4FU
abftrsmw2SLicGqyZFyJ8TfwQE1vsgT23MOmq+YHWC1ubAu/WmqK7osqD2B7RWtbpkX8NECT0yD5
KEBIaqMXPjiSlIdav7JtosLGDWu45uAxyqfhfyNZy2DOIAFHg4GizOcjvfVxQxbt1KO/d0X2X9sw
rP0hri/Rd0yQUxUYJ6TgXiO6IKv4FM6c2ihEk6JDw0Ekh0JQ1qtf5Nlk0hML2+vmyVMA0fY9gnk7
ay2Y1Q2PQRAEF6U6aOxL+p9/T7pqy8mSzdhuZkhetDMvJ5QQhf/MLugKEu8BeX0hyqzN0/udlain
1aXbSh+Ot4Lg7jnXoBJ8NxYbUC2L7el5UeR9R88MzlH8vhuUWfZA1rycvVBkAmqnCyReNdOGL9si
J91sWyvrcSyX7AKW/pn4v3bslqPmVvywKUy8ORg5lqXu2u99HGPUq7y0pfOe3N3GCD48eHB/aBoC
3iRJtV5saXzDp12Ho+H0iVS+ZuOVSvNogbf7ewwChgi5TKip/2djACJZ2k2OGx0OAiVYLzm8iJcW
eHtkzUgncNURW9MIwlJEyrK6Pa6aXW5jSbWedVLYgTq1PcddVbwbnMsTtBVO37a/x8Z4YPRrHB7b
9QxEsqKakONh2b3QuWpzWqWeWZxCQKcg0/P7miSSIgpAwMF74vouwdQoQ4k1CGJX+wzu1B0VllAR
Nw0oAmO6g+ROlwP8/uX88JgEqjtxcLB7DFx9dpNfs/EP8ai0Puk8HDK3sTLeDLdFA36vDfI/L4e/
aPvDdUqlREb0O60o6bgvs6reBH/L1KZsKGWHhBhvR/ghmnWyjG59f17Pyq1G8fYVIMdHEtCAYxdV
7fiGo6KVg6jlZTH78nnp/rRg5f8PqnShmxcTBs8C2gEix2IuzQkjdrvKs37QxFAp4b39sPKF/+Vk
iaXFLzMDGvPx5jsedwgayR6tojpjzo/8tVMUfcC/jKkCyGPbVaYSz8Lm/NKymufBU5RwZGP7thn4
QpHAriMiglKCb5DJIamJctGbUeP9k3hXYQza64Tq0qIY0vwMKPTN5Vw7Gcah72aNzGptoaBRs8Aj
cOl/sweu24v1OoG/rmlzxHbLGnyrF+0fEo39DpuLXSb4CpP+XLHhSJWrty05W36b+xIaglZEtBlG
mtrDmtbYHZ1Q/AqQV0mInGswjaeobS9+tVfPhMQsc1Jphr4tKqCjIsQxQlUcxtSFAu9Ogahp3xfD
xObbVdNL6IEXJ/4qFMXz0XNv28w/NW11xmt7U91Ge9YuOCvTzefavy2UUhYCOJ8r9Ziqxr175/Dt
YeGuREfLBwQmp15aA4L3NVqd5AYsKBO0Q2OaFPzkZH5N5ztQg88/Ob7uEaDwk9A3Xii9cBvLcbNg
p3HNLSb5Y03+EKzKyaKACAl6cKjOjZqtHa+scp1o9ng9HNyd/ypcryvTTcEYt6rWENEhMsEwMKm8
CRoytmZ/BWkqa7rOdhT6ZawY7gXmHOIhNV3V16RSQJcFrzb0QU0Q+4WWswTVrgHOHfQHH5MT1k84
Ny2YBpsi+InGZTiy+VIxzTkwHnbkFE4/l3sGU1/B6ibLuS5ckuKmEU+U4QWtX0H+3rIR8H/4ygVF
AV3lnazk+S5NOIjws6oy1KZHCwP8QIL+0SSVMUmtuioGXqabKYiQQXNDHWhmX/iOIptb8uhOLw7l
oDZ5Mr6+3h7gXsEQ2kmtKf1cjdjy1dWHJKlaZECq40vMwx/Wc4dZik0EYD6LgifZHQnP3KesRW+4
tDyQGMnla/s9t6b9Mtj36S2srxdzWuW9AtR1SLN305r7/vT8SWLZcoPkkRk0iZu4ESBc7Wo8AvdX
ZYNwc/T7VsLIrLzozL8bVEoqubU3ZhUKYAZViNEAvrUx1QKnq75uqnuiKWcex29KuLhYjHGHwv/0
g+czvHzr4xeC/uud24qZq/z1L0pb/SjQVo+ePoej4bRqJ9ToaJT/JuDstjCPUEMe726KWjN/3cZU
WCrD4eMuonEKJz7hwVXilu+jQFhR0gIyyb7gOP8Dphu1o/5LxSnWnpJzM+BAaZmh5cKaVC7JybLd
Nngzf5nDDJFstYg999vVLjjC//ggGYm1nATaLM1q7kOD1rd3kdQzBp4uGdBfew2PeINaBOXFGv03
ZnbDjDurxdGRgC3eXqUZYO84OWIdlRwzBP+0OA2Xz4aFksPljJOum0Pkmu9sdpgqNCqq7whN7SDW
i33qtJa4YvkSXJSJ1/p5Nl6GXBKvnzZTAbuAS9iGeXkPXl8hGKDpDRSKAsyukMhzPhHvrzwKahFO
fnO4PnBQDfA4tJF4hBJDM6JG6VXDHvANJfomNJ6XXgE4dHOWQIjpjBPMFdXZ81aLYLFJEN/NrUSD
vVG1Mi76CX8U75GfL3od5yGfXcGjEfEUdPNm2IeQavXczT7uduQFN9IYNwteqAOnBiKow2boTabg
OrPLrK1K0PTvWSLyGUHRzW7J/ojlzV/HPL0pGi9sO6L9AM0uL6VSIpjERdUg+udHAFTVYcmBXLL9
/azBu9NS1NUEHcJjSsLLjCLI/ny0Wv7RTtDV8tN4nWdfpDv35LFsN8h86PgONp7eWgaZpEDKekbd
qHSP1Jo0JWJBHjccPIHMTx6CsTuD/oTrDVlb/Ew7hTWuAYvUTZqb6iHp7S/N9aPjxa4RlEW5AJh4
BccW27eAq6iYqYuwD1ggf+e3bb8ajfLHSMh+RjPZy+jT3AjASS6/6pNWkiQ6TMcI2AhOgNdHjQbd
NbH0soQMPJodR41TATWZqBg/qksDwq5rm5vrPFqO0oo+IztzsoP93T5MpT0m1SvcjHZ8Q/Q/q/vC
YOV8LOWSp52b4+QSVTlNdIPzN30xK18iyCeMOjr/RlJwH315fRY3JnjiSNcNowraG6/UASnNLJaj
8hhMOBx44I7pw07FkikpyqkZBUX5TyNi+LuYy8oIvPKKmRAoZxqM2faUq6AkzUK4Xv8RAMPI38bO
+zTlgbJwUeoegSOm/SY85uwKr1hwroLZSdkYoT+Z+BU8qLw6+/rO/9P4c+Hzz/vBdtPCRnCE8v3g
zAmdqNUUcll6UJVjIqPQWwZUXcB0U6lGHa69YpqG1W2ou0II3FICeIuiSmGReS5VFJ6muO80wX15
7dl5Y3Pei+ITf22IaRrxv4YN8BjfIoXbscqP0vSVINw/TXlkjrUYNkowFS5WZenMLG4DCO0ahEL5
2XYfbax0NNpqy9SwEGVMaKUtDnRHSixt0jwaGhm+Qh5+TU0LMJKKHwb4GAs74pjSfMDh94FpyuFv
sDY8dt14TNrXPJZcNyD6h1787OnRG/qqIsLXMmbDguIKFjVOfZm43qD0XjD09ITT+KXazOuE6DzR
Xo7IBE1k0rdMVDLW+lN0JjRaEkgyDWz35WfXEuzx3ua6gD9Vxy7qUkI4CYLIbpgYMFKySl/hGm8Y
L3oUdVvXO0W9EN1sQE8QALcl5H0ZvZbwdXUbQkIbJl4e2teD96N5ImsAx+JGW/unO33+OzJx8Zei
UnTfLNANhfTatY5OuzWqcZW2q4l3bTnVrgIkNphPwhLpzIMV3osNAYMFFDZcPVsHa77wH8fVu+lw
Fm8/A+Lk4JCNN098WSLM9L62ojXl3wISYJOJ8kttFQEVGvNfhGtZvAfIUtKXhdHgW0ErOBVM7MIF
Mm1J09JuJYIwOh63RSOdUWuej6DOP1UG1xirPh03NpsrEfVeRbGl8ie7lo+fNQJUow5pQnT3a7QU
YihhPspQBNFog800xfwej81murHnUnBWwM/y5VRsCS6vC8Z776vOtUVP7VEpYYlFMUlaG3K18qss
+cjUnElxB4ZaLn447VWc14HZ1zL0ss0IfjFjC7AGvI0QueHRmpC6DghTBL9FJaUo0YAh7IUAU2cz
N9khD22pmZt016evOMF6k/FHgp/lD8QziG1Gw3eFS8emScfpLX+L4vMOXwa5j4+1knDMxxdVnmC7
AIQ/OsYKQOJWOesxHDkjdIjgBbg/beX8YM/K+ysk9XaY+u04jczzBoyTpaZqbzqCAAScL78rSB5i
V4wFHnM2yussRLupKzgNLRVTu5x3ZO5Tmknu5iFvQS6wKOmsuZMdNZOCIB808MQEB+QWoUGj13r3
EtKOCbt32RRTlqRtaoTxp0n8piJa1zr7OdvnEPViyq1fBQrUKE/Z7AhbcoPuO5y5T4iAj3D3qPFb
5/ohvFy42WxutOZqDjG85zgrcJ5suhXnDHaj6e+JRG5AY8NkSjEawnWTZAxrkPaD1zgOHe33Z390
IieVoLJhy+z11N40ANFCRFho6yQxAosfpb9xocknOOLi2KHXbyTUHWc8xMpfNYGFLRFEnyOCYM/c
CujRDfd98iwOOYDxPpNEWkqKKu7kGxCcIblOUUoOycW2rF5eO/31noOD9nfnNzP93Lzz27P19rmn
C1xJ+jhV0JjNnd1z3YBdSgPwsxqhx3GfspJuBJugbSta8zAJk+UX6bfOXpdm0rDKD6RoGqGc9D6j
w0GPHgrOW4W8hDe+MO2RQ8xSynmHkodzR++IlwEnHbtsPjhNjJDgakrVNADdAIGZs4tsXZEq/5Yv
+CuowyVqqXzlvU1popUNSQtA6ygqA0Cy1R/FgsaCtxD4F94i7nhZ/ZAUfNxl1md0/e1v2S2fgIgV
xp2o5kbrySiVI4v+9uEQJEPosHe31k5OeKJqKntTK7d1lWsFQaEzRcXZe4nRBTHhU5+KX10uGeNl
6GETmIz5qoQAzCKuGSvSqvMZcBoyvZF0RcZYgL+XlZjKoYUFH3CaPRsuU+Gq39/HWWcv15q4zlws
80Md7cqlWwftz90AZAPoqqM9Fm7926ak5J2Dx0yRP/41qNsb7tdpWbEPQTyo4p73qlpDWQo3864h
PoUbU4B/O3HNK2gU3ut/Oq60e0RTbm/FyN+YyoSQbEk4LV8sa+c6zc2ZGlhELZ2GxfI4rHXj++0C
xgcf1UnS3nUX3ceV8DOa/vwp4CTUzt7um+b4+2SBcwc3Rgp96lnhxXL9YPALHq6nR75jSAmgiDYw
m5FxcEV0dxeiwlbrZNcwq3098mQWndXNk6En8Xe0y3c7x+ozjfdSzvzDr7mO7d4H9H2Qq5lHzqkd
iClFUidtq0FFZlD8IvO5Ik4iANZG3qK/2EkrrTNr+ST7KMx/+ikM573HNIFzsQXX3srIk+iHQqu/
0uW0X+PCXnMCT2xRCvqPdsqxADvwymqFVyPQOvaNWxve+erHxF+7Ji9SsXSrSLrFpbd5IQxXUXnQ
VqGj/bJFmubqox476DON4rwepYCCpIa9XfVUidKyq31JdW2iCqW8Dk0UO/cl1cvWZdkFeW+mCz+X
PkJEpjYFrOLkeo+7Hh3VJt5yyeo+Gl93BAcW2lRGWFKjv3xGBTGHOs/nUvReetyVmtsQOiw5do5n
qAgkEunyGFO/mH8NgLD8AltN+nclN10BI6xaNWKTJmEZ1LRmqgb6TBTctfMoZ7rClG6EfETxPq5M
/ahVYUy+PkxcfAlREdxViZ9QKXgUlLaIFU/06QWsIBEb6zhngFwunUXbQHRxhEWrysfnlvCYouEF
C1ygNIzbc8oH90SEGrL1xIX+yDU0kycoj3wj+sLx42VQr9bpQBqb5IwDHQclJx6jbLm4t2hnfxkW
BI1l1ZqL46UMufByYOkpyjqGBdUxAx2WchefHSvVzY9ap6+6dVE0c2xuHAUpc268KyV1DFFkzTB9
qk9tm19Sq+skE3b/HrS+bODH8msKSlkTwaVNixK6sa5bjIkOVtaM/zv+6Bh7Ie/lyb4u6Ag4+mJ9
Hwu8DT9OFIf366ruMdxa8fUS9k+tmoCZ7btlt+ih9UspnDs3LI8UkoAPWC6QRk6DBO+zoSAU3y4w
KsEo/c25MhRHhgmfHXhiG08fahjIxp4yEbs88BPj6/TEDiq5bC4haukB4Ogp7DMJ7tH2g5UzSHi3
vSp8sOm8aFPkeln5kPhTkR12D8PYBue2uhYq0DmH6gsgxMtzfCbT3VzJdIsgP+B9PyN5k8M/gJ7y
mFZbZVZgr2z6CqHOoclKfxPgPyxHsmhIC1d4F9IaS2OCaJTkog0qeyo6/DhBsUxaa+y0Y9896eNH
NhTuF0DbEZgU1FA8mj1sqTX96t4v4PXyzY5tNC1rU1QGBEXaEtN5wW9NflQrbfnqMT2Bhjc+F/r0
wn+wSNvp+kXSay8yR25oWlIjGnMxbDU2OYumDcCg2V4+8+wpuh0b9hx726jtFSqs1juCqjPlI55a
kwPj72oR+kBnm12wB2KCmw1B6UexUv/e0ARRhxUhWgLu8MjybuXZhEzct1jYouBO+Bpyc5UHtYV+
TebJb4wr9JzWHJGohW5PBtRDARGGqXM3eY713Rr5+nBAPw4ugBl+mkqpqn8u4QrCrWaPdQQKrp6h
FuJ0srgpqYYI8OLDGZP9UB9DnH1wmEcHNQMwkdXZCUspIzOXAEE7RJDU+eKwmgNFUpOLSyTeFqjV
OFILRdLaoZMU/3Zujw3wK0KgQJVF1U7vCpRZhxZQJJm3pAxqlWLgu4fR/q4ZBoQ2Cp56cuU/s21+
IUnh0alNDdVUyUqtkv7W5/BiAZ26sSRFjylD5LA5mK9RUPgrxqq/PVDSGdmb9Sr1FdC5i5DW2SSy
kmKgvXRNcUx9DvISUBsTjw5F4vw9vtk+PAUHsYwRmzCDOBM8Dt26Zq7hLkSvfOYZBcmyW57YDznb
i3oyIvj2UQ/AOd/40Uzj8Jv2pIRPhOt/VzG0F4ZXe0+KpOZNRcyjZb98oMQ9menbOEDi54t8wfXK
aPbKwO4MhxVv5KfZwKUYrQRloKMImtHOnqW4JObjhXV4Ntg6UC02bTaQJTAIECm3SOp/7Pt55oII
w0AtbZDGVEzui6RV8wUp2TfhhF0htOb7NLaOpdOEf2Hilxj6oPPQ9czVRJgCMGLc1jAL9Pi3JmKh
bojk9ktZhoiJjkiEjAHa+7tykZhwgp9CyiJL1+M/Yb+5Zzbiis2e8SF3y0Vz3tCnW1mnla9hhQti
ZySaPBW7+CAvKaGESuyH7aiZJ5rk9w2MvZsUFAyw31FAp+9XF57lWgEpVCCotbPObUYIXOmjj3c6
RJWwmnK5ASYQSdbvC24KixN0fCc9G1+OqrRNqEx+JiBqOsNbp4AuUL7FiWHPN11NWQxKMrGnVX3X
7hOZ9ZA8KBI8uNyCPHnqqddNveLqEsbunETEnyOaFLSYAGMeGI2AYMjAJozQPt+NfDIrqWDLPMmO
RdqaL6G1bxF8muAzYIdufHD12rYrrqY9yFuD9Fq4jo/Gd4kS41W2nU5UzEYh5Q94GRWO6rZvrzFh
vT8ZLIbXjQoKf0Pg6qOgjF2si0AicsJoPbCiJI7mt2RuS8OzP7Wfx4WZexprCTdawV2Rwwly3TKu
9EJ2aizVUMfIGDVs2FSXuPPtc6aF4grSktPZbRI1YMKnVntHNpWXRkc7n8ReQFHSFs+2g3MdpQJv
s31XXWk61jograOrrSERFvuhMlqNDDF39KW//Pkt7CdlZ565msL/haGEEB0onmSD4CPXQ6Cy2XEy
pa4X2gXWtH05bmvh9uX2UlueMHp3Lo4afvikhN8fZ5r5jQvicvkAubALgoQ3y3ESaLj3d7GTiMzH
hRYy+hfFVgJtTitahAo1PEek1Lzv12Y1IyQOcGyOlsvQ/cQ66y4iA+nm7/+oHeqqn050Xy8l4qRS
Q313Ns9EO82lTKqdqPduupiGWSMPkN/+8iJLBKI1KI+mksh0rAM7yXxLEPC7ongVEvuoM8yTp/DK
qZovCtcNlIxgDQcC5SO1sVGTgM9iqAUIJt9y/DY2qcnFTB/IjIAfUnm9oQKSDxzAfAAgwNZEbSlT
fq9Uw2Rx0lD5p0+6NmDftlAgSmumRUxxcTYAH5zZ9n1pbH3ZqNpaezbM9rrGTKn0TAvBcRFs/QM9
ZQqNihgkUCZg3jOY1vKfVUQVyxwbCB0kcFCHTwCaHOILKvJFhC3kwQ7m/srSPKTUPO+iHIITtxGJ
fMVLYA7IMhU0tSWJYRg1a739Co4ubLdRFJEla+247pn6tIukgg9auWjdKSO5e3/z2smcz7jOIt5j
f4a9eve6vAokJP6L5ANA+1vjdvGWs492jsJ/K8gzb/gBSfaPt0FvMRqY49BOTuJpEMxZqYwJH8nt
68o0+nvIWZi2WelEmt4GRkx177hzE9+KRuMrnvvdCZYBwsumryndc7Fi2f3BL2/fy9J7AIyxLDl2
kl+dCP6M879Fo8/rqErzlNwZEx635qgJotRCRhe01g6eZbSTM2pl69mqAEFhGnQ8AKXUNco+AkUq
zOavV/fgaHWO6xTiB5sPhMnbN7MSXAm3WV2cFB8hwPH7Zw3onYr99dO2827GMzWitiYVyi3Wo58s
D6gd2MGkcn+IF8U/2/YLxu5kbqGx3bgVgz+pu7owwl98XGzbqv8lI05y8YkqICFZXD+EHaudkcQh
pJIT6tUozDaMuro6eoasQhKPpM7Ef0i5O4aakF/083NAX/yfY5n7dVeiRHY3JMs8clConMfbsLW/
su58b2xa2GwAuqxTc9J6CbEPINCnzIShg88NeiJigj6ABcvaA8jebCEWDHcGVOYjYq++xc+4QMox
mQ7VN5Dei1rHKrKsO1Nu6CJ4CXRqZpBQXUSj3VxbI8/egLvDiddBohmOdoQfC9wPwuc2t8e0B7Wd
oHmqdMj5QXOcB1Bd8LNFJC4+qAgRWURdBRhk8dEc8GnuCSDEjCZhCHQn3+RtYe1ljVFGvcn1M/Dq
oJsGjrEp2KuAK8VZz3tZ3rVB5HIMJPs1TdpH6GUEdGsEY7uk6BrQxDQHkVICkZVdsTrxbNN9Bp+Z
/6P6Xm9hazMwBV7XiGK7oxadXRiaqek0y8Cm5s8cbsI0ueXkyn1unI32ndGQVyJT6vYjOqMLihvY
LrlTmwEcG4BkkqzpY8O+P16CcU+1pjFH4CG+Wf3262olBn31B46aJGny39ZmFqNLFZTFGxDEVlq+
r9swvLAQzobDNSDcN3VIlqGsSi9caZ/TcpzV15EGBDdf8rMszaj11Jlg590HqKTAcP86VIClDvct
j6yCSQ5vWzKTLuGLpDtH78T7eVYOw+pDawyuDbJUAuo5u+JbmY1T1dn0XEgUHqg3F+4iUqK17VCM
1tVZAEJjRCbweaCCOHxiG8+r3P9+WQHFduRxvFXswod2wPDlEf1iOg2KaemngKsWbUEWPH2RnMrc
L0z5QvzqMpY+BKKb8Imbj5wkdOcFpm+DM1OsspPXYEcPCSqnd+lbWXf/doPhUJbvC01Ky5i/2Uz+
7p6aWzcEV98k11ayZEEaOVP9Oz+SwVmToAgZ+4/j+X/gu9oyUOe5WJkBm5+5e0PANIPQ2NR9Cvem
dYgFg0pBNcYJU8i51MQohD48YfZGVXSSu4b6+F2jRXzJglrD/RD73IXpf47CjUNa7a5qOdxts6Nw
pSd+YbhLr8nT17O9bnUhsUCcqJUbjOQFpWiuEn7/vaNBckAV2uoqVLH5wDfQ9vwRyiR5o+iAO3CK
77FYAr7U5ARzMiV3SlCgrLkZZYsP/Acd+1F8coKkGuAnlyb5YlfwPl8fQZxbkmJroETUmJBVtBEC
61S4W15IJlegrCFbTLctUREftPkgbnFHqNFqByQAnSxVUJUX6Q6xITJFuqZl5KkVjID2dRmxUYoU
d+CKDDqqWaa1C9iR2fX9cDURtgVwgSveLyqW2OjIlmfC0jd0FpwKVo8/70c1/ZUff+Eh8g75m69r
Cy8P++XfBczv2zsIcJH98crvrEpFdgytOdOCqGvh0gYZ1HyFjP0TOCJUdPUTQO97Mc+mdihodvKp
LpuAoWn3M+OwYK/GQh/qYcwFZutAAibXJ64GfYfqM+3j+ZrqNaGQ2Tkt06eUw0DHPFwphJUcJ+EM
FRteygEd3NE41St1dOv1V6EoGgfThpYHVGlPQMf7+9KUQZruT0W/3gLVmTzzjle4vZfFDvPNaP83
q1t8ORkBAaH3bSekmO6BYU64u8Fsn8SVD13ExE+kxzgCOLd+IdTbxWkwVD2mcvZG7wnHaEHdQRr4
C5qlFVxnMjX1UDX2INXlH98Y0TvFXRtK7V/y0JEgvcQP9IDnZ7e2bIZFlsjwhUsq4KeAQX+wMiCN
JWPQxQTszxQtHycNcn52b8eBEAlAPmqbuoIopp4qjArzhjJZi3oVZ8FEHEPSfjAFnlYuiA6dEcEC
rwkHKjl8t3tb36t3CkzI//SJzZiB5Nl8s/ty1Akd+Rd4YatiDjUwlPbXRJuue++qH4OjsfuIAQPk
Aycd69Ti6n4Vg+gtYwjGC8AnNVBmgzCJR5LBsho4S+BDEstW7Y7l7GQg4d6JE/ZugZU6UNCs8H90
ceHRqlKZmL7Bodh+fK74XoBvpwN/KiVvQNdVGRyTTZqoUC6bIsPLOvc5k/yOdkXbyfVkvb3J0KKv
kGu9eU/+NgP/Q4p9MpmStVb4F6rdW/TVN/wS/bwXGVcxdB0TZJQrnwc3k1SQLk8aHZe9MVZ4bO3w
4yEqh/n23h3B4j8lHOVdnE4Mca2bvDP+0Ogd8taKqzfc+5gpLDwX0qnrslE53D87kajzJANey3w9
EGZ5cAsQqaIEBh9RdyX2A7gxxCrAeFi4TohpizBHy2d2/awNQrYxFMqIvuEznU0yNXIY9PiyFynD
IaxFUaRJyJrlw3InQ6cPODPepveFJSWdXBRj7P/QWsk2WsmCPjUArji1DifS8uUm/ES7PbJCk7l3
8RWuJk4s6/1EG78LaLrx6YNX0u7sKMr/56vsHqf13qoBrAzSDHS6tOTOQ2S0dlmOnIftEgEhcKS1
jNU6tBRNG3j78r9RQcFD4PjT/1l4ePbxCajFn18ty6k8K3zhn8X4vir0GLnfnKgzETLgPcxWSwzi
o+k1qyJbHEGDTo5o+NO00Xdtxtp4hE4IN7O7Dgl5FVcHmXQeYFcLtA4yNKx1deEfNCsqCOMn4nMb
Pi0mOrFbICOZwTeka8AclwtiYVZd0XO24muHWT5kHO3uvWL3jHZEnSMNxR/4ybcuVPOUzrMYfNby
QUbECNsTqpUbtSp+w/NPPkYw1deqFZau8uA/mIPMQcF0pr6fOHkpdwDn7JkBodzbhsxilkRuZpQE
7XM1FBES6s0X2eklfVaTNqQsrw1h1NRT6M8TGnE6WLV8GD4qznV6qZkyrA4jKC1EF/fSf9JfK8sD
gLi8yWl/9mrnVoBgMx4N80IKweK3DgyXghsjuhafRgr3vy3UaseWCYCvetb9hXTDCFqzFaC73nI+
CFNqQpbhfxDXhqi1mrjgIXj3+iYCEkWfPHk/i6uZPTkvPZE9tHWsogXO1SvyMURaun+GMAcTsp0K
a644mM7IkcMGIeJtLl1/XDKX2i5j28oQmmPZrpc/ECCQfycFts8I9FAvrJEEn4A+2Aa/bgizA/wH
9Gg/ehxdSzU4M3yJkv4QFSuMawCelLmAR3rtJyXVRfFmaV5n/iushajplU6HIuExWhywPeAtmZ/r
K7H45CUB+cQsJSFjCmjj+R3CGnLyoDeWT9hHWk6VFNqLWM3VaFbDmif1yUKy4SSjCSq4QESVrvti
drsuK7L+aZiFAUj2U5SLu+ENUPGPcW9gMBBfJZcAcYvIcxEEVYtU5P3Ho3sB8Mu8h0uOlSYtqp0c
SjE1eqDtSnEaIw++XVN7G86yLHQjxP4tEzK5N4PN8dRlsEmzM2HoqwnWGZbEA4Nf89IvfSE0ku1R
jE1EYzS0tj7eVyXFedyHfhGNoRw2m1L3RjE+aTUuwYYxWdl4DkkxiwmyheKOQsk/o9ZAGZeAViai
LDWClKR2VxiO5m9QQzOkj/8MYLxJGOCIPBoNE7Q/q024zaquNC930eTsaClq68YPmQG84ZXs5mgh
iZsV/2V9PXXoGEeNqdJHtfUQeP0+vrPpb1yp0Ag8VzME51YD1ArDnlW7FjJviTAaHUGgPv4f2Fny
Ywya5bMuhzrsVJeC7MvXm0NspAvXy/qE0OKxQIc3sRdl5d8JgGDb369z7xM+uIhHfXmv4rJxa/BE
IarxqwHIZlL7aG/x7OV+eDR4gXdQ8Hlzn4pS0qCovhzKasqxpRJDF5YueukM5A86BccHlIMAJWXs
C33waUVGGJZ8zleQQy2giwUgNdn42q77pZoE3LfsJnAwKBrKFd4MVPQ5LJGZBatZQcodxh2iGITS
METp6dZ8SRKSQLi3BHTlLUkPfKIhl/OcBlbtyowRyXjoZ3R+wOkUfKBNLRxZ2Gj+5HR/aUPXtHzG
nOjX077DYcnz6qzRmMF/vpF+VpuS96JfigfUbcDeTVSJ5iWXoo9Bsv8DoNI/upr/u0YpeuK6VGwh
pjuAdss0hoN0/SS1dDZAdtm9qKDPt/JgiujNtTdDqPn4w9cIQhTPyrVTIBvd2yVOR0fvmCHuYgux
Yy4FVV8awLawJtolU7YrtBv6+yO2lbjN70bx/6u03yum9A9DIAyW8gqVANBxBZ68VqOe/VTHCNHE
paWD34PlnmxhE4E+1UwOy01mxGOOH1WmRtZO3hy9AIopl9C/eDNoIbGLg1+CuWK7xLM9sV3kRV2q
F7fRqHTvaxQN2Lmr5WN8ef160zWmf1oxQDUP5YLVy7JKifGgYA1qD69vTUhr9XwjB+g6acGoPfXS
1tWRCcZnjWJNfV19bTC9nF8P/C5ej4fsdzd+0biLX0VFoPKFkgoxFxCD8+NefUPGhaJSVdF7qRgn
F2AHOTjAMNstrhJiDmtSh5zs1z1CrX2Mo8IABxdsPiWXwzrf9270r/0Jwx5/Ll3LYcAYNPqvbmo/
Fyu49zOu35rZJSxFtn00NB4TkKWsUrqAg0gSHUqJDK++I57UxOAD5v5H9WENA0ngbiIj9K238fVC
17KItTlYEh2nvB6pls0FyWwlEyT+WgbHg8korjtIun9STSTTs/UmQWsi5J/TC94vcDDqtBtjfzvK
IJj0Jw7QZPtZEHTZWzexXK1jm5ZGjB9pHBNjrEB1wFDbmWQoMN8YKCuX6YH+YQdagJggJWIDJZeF
R5J98VLTa+B9F2+reV3Ct6yZQT+Mg5YsIGW8nXzebIZIDZdnOMyovIXCPddk7EuX9c3057t8imyG
z2B+kk2q7Fp8l0uvR1DPRgoBPq87RqxQ+SrSXjBTlFjwcgVeBlR5Bg9AiSNz8qW62x6qHOuuASaZ
cO0JWLU4aVvyggqRw8owlDiRT4PplolBVn4NVEhjk9drp9/MuQVcN6k+VA5BJwXj7ei4SIXn4+JF
IAo7TEggXXm50w93wSEgq/POI8y6oBTmR7koaNoEdSabjqqKrDWOsekTUJr+UUc8H0sisQ+m8BkH
1XQgKefm6RnPvi6P128IA3WPWanw+hM4aHewyyhc/rVmW5x3ajqve1DmCegof7c/TyRGcjVWmUfo
P9HKuanmsitsWZ1GC8AIMyvAUCqsvd33RW/e5Rl5fnxt0Gx8RZ1LribCEgXdDtZ68JqNtkBvgW3V
pKN/EwcHfDKTgmQ4MqHMP9uFfpGLdm/lOMLzXVum1Exsfyqk+pW6f6ukWlMuYRElicSvE1Oee6DG
IyW9a6dLMaqZo+PXXU7csuGHOMqDWcbs43IPOtVfmiPpiXbkMncrbu3+X5oS/y3KtE01Xzak6PSN
CBI+b86c7SuWtvHzzyrletoRJYVIO1VUIx3QW1F1wETgA2u0BcHTJkISIXSN1zYChLR+4Myf6KCY
2GWOnEzBXkhb+6uFm4SQLhkje9Npbo6/ibB+QOPi9Zxu4qiYG414N4/eaZifv61oSBu1+Ue/LriA
bB8+8HFvfgQQNBYFA+o2TWe7jDhsnq3QFSa5McX+iG9h68Bh6FgHb4T8WjQ44c/c+tpieA/rE3My
T43GwpNOm1528nRf3wxhPs3cZhwmn1rC5N5x4eclgkfvWRaNzuS3C+ZViRNBqghzxMRGtRiQgkZb
BlelYvdplg5vz4/d76muRTWJU5000MHAQNp+1eTQjyFWRsU8n+1+PgOGb5XuFPoWEyomI7z3qeiT
M67BDzxJ5URT3LXw4Jpe8V1y6Rerk3DMGQOLc6c3VcVi1H1iMOtl6eKcJgLHPRLnjQoH7s6NFns9
VTWutEk37LmyCN98YL6rVbr5Y54w2KLv9hD1axgd2/yNGBwuyw/uNbeBmg7jH/X54ZzOQ+2AnYnz
bOJ5wLGhSCJCQCfrba/54BcIFNccVb8kC30UPYVKiMg+gj+KcBSXZFCVACGA5N7U/quQi2jypXLe
B9EwMUC3g9jOxsHhAtbFbqJ6XkVch6pOTaaThFb3LY87LddJagj4caxcPheuJizjgUNK5xVepceJ
yb3xoMklPGzLAmmf1hnWidVD0tlCuAXs0Z5oZvkUzCjOSJW4x1nafzmp40sciKMVvOHzT8rC8LN9
53OZspmYqgE6kiV/Bceo/q1+r8YCA11dO++1zNsmZp/A3ZoV6mqNSzADGnGY/W/R9hYdH7xddoxg
pAY7uvaW95tQVIXHMJEBWe5IEnhXEbTuFyfYNMPg2rmZMzNjQ4QjwQ5bOOCf/Ks0VzUJD3trx4G4
Nn7+kt+qx7NIbxb4xb/cP9N86kmfE2mKxfTUHHWRe17k0HDCdI/iyCFycdi6FCeieXGLmoi0pG3D
lCDU68lyDNpVU7ilHVpXmWPyXnd36YOqNW75YJjR0EjhXf7mC1gBhlLLDt0suPBk1kOOEM0OK9ud
PvUhE8+TJ5o5gMo/w9zc7mAJwsHKopeOk+aCHywe7uY8DIXD4AkJpne39WiQw8ZbzgjBAILa6fs8
eFyASO3dfuG0q1Pdck9qXPE+qCc3RxXxBB+/yDDH24wbHxaylru2pA9o92TQ4nWUgVJaQq0U3T9g
U6kz004GqAfQx5gpe8uWqR41wyyrjyaGdyugvbi0W7Z+MUwDRgK7zYPa7+YwNbC8Rw9gYvm+mkwz
h/HvP0BPt90IMUkLgmCUOh9W9hoKPRy+3MagZoRCkPgO6WwXklAlOAJAvKlsISOt2b/s9dtjvHmm
DnalUEw7NvyOxTXXe6kuGlmZOjG+ZW5f5aofsJd/pqv1lbj34AR+qsQV7ZIKZH3OGjFfZLOR//fp
XYNHGyvlHYCh4L590ppbxhVs9VTLdXdMz2DSsKBsgHUoPxZHL+GGxCpnG+Oo2isW/NrVN1OZyER8
yWIbfdwcWDyzr0arMHr1BeODdYVOGn3K92qi1WKOKvpyzmgSW/NXwNKpGL6xchzDqKHOcJPThsGP
nvg1z6HHzTFAoe5Bwcbo+d8yh6k2rUi92vqWm/cQ8BCo9y3ESI6InOjjWIiPQoIiUYYH0qq/y1H7
7OF3CcaDz4NmmBT3/x2twoqrdyFdeYqzUIeTC3KUC2hE4WAFaY1ByCcPwpzIZRuDaLoFD33OG0WL
h/XzGenwfDGLx3m+PK+JBUvgEehAOjrE+QGxgIBT6Mr0D/PPp5DMuQb/0iq1ek0IqdgZTYHU2ira
XZAB0Lgw6e5khNqLnS6jM3KMNE0jvi+0Zd572mnPEEzTWJTkAKMncKM6zDUg7gTZWV3gpBq8XS8Y
R0kB53Mqc070srL3p0jvHyOiSPJfgy/3NE65w8ASOWnvLpn1Ja5+r8xnvGdDeiwpiXlfRXkCIJPt
YgUvH/AACT+ApqNXpPuP+5s8KgJTCx8xLG1B9JLUUF4N+EQffx3CQjLkjif5wbqUoDZeqU3V19I8
cjjKC7qxVodiNXHaGHwCMKREueF8/k/kdEzbiYcG1sw4d0G9IwQxUO0pMzfnNzFyfD6nhmXmrsks
t3pkJ2AKdgOOFGKhSitbsTDKZ7FZn8PnIAOZzUdJHbgquZhrd9GR9JZfiPCqPXyE3M74auBV41aS
KHDxjh2zJs3Ph+Izs/Rjz1LjSCAxJMzfLMqeL2eSEGSws8UUvDfPsIbvBTihjcA3sIrND7/VdXEn
3VGF0vcSmMtCnXdmCb27dGS1czQ/JGh/rfpow2W5GTTs0YngDxRyH51Jkb7NghgCH3WYhbNjcp2L
9HwzZ/JENUE3kzu2F/efQHNWfnOF3L15wPlvAf+gJz0FSJp8lf8CzrKmTi3v6XgLhQ57piOCKKVI
FNpw9V1ns21L7/kDP+ZNWwjpybOuRxk2f0SduO96ElNb6PQadc/Vm/FpN9pPZwbvscn7Z8yFiqLF
CXe0DauqWLjTZ7Cg5xf4H/epAYJJ6BklTcOfAUYPYOAeiLuhyPvuh3E4jv8Xf4DpEiF1iEJODtO6
0YMy8AHmUduPS9K3K92zQuhDVIO6PcwvC6aDZSQFeLtSjN0lT4zliEsNKFC9AywyY+wtW2ABV6ju
aouNFsDCCekm6oo2HYePuWwEp/g9D8BtKwtPas7mFlZ4JUVCbAtb7tR21KM7MDo5zS6R0dGUNc5K
JHYKs7+tKXdwTm6YrfWnIfA6PDXlovYo62AvzCDy6KO+FIVsLCy+XPzxAw0RP2g4iWyklJ6o/5rs
c4Up7Dz7UNAKjqouJYM2Gbi9W+TNoMEw+U+R2znA7BFCZVHcOqdrXq8Yvim6mH0Df1PYHIiFz2H0
JjZ1tg4ihvWE+581OLSuvfdUagG6T12xMf2SZ82q8mljnf+rTHs1CMZ/fgwNmpUpGTn8fj3Dv3W1
jyDVOuZMyRwc81pUhEWlJOMKMzIjPPIamHqMDQ3m8Rtg1vgWxnxakgARGHHJc+JEyFQWRcqgmwf2
QQvxgJNWyNuVdqLSFiILzX/ZQuBlLHt2DYWsoffPTDvrIC37BFcSB/xGTONc8GghzTLToU7vgpkO
mGfp1tuPsfqmh2XdebqgtOdWtDkbJc6BzVQqeav0czb4tOQa56EDk/xSnS8G0Nu8gycO6oQ9Xl11
UoErjJiSM5BIgIJ1MkEGJBWVDKaWbUDDEJTlchZa9sjvy38GI41No7p28A/Kt/aPI5JMV4RYujvR
5lqNq/sFqFIk4KJXs2h6bOhEGWjJjhPFP3nrWW1sPK8zLJdCUX5jXVE6R3a9Ve27a1+WbObKEahN
xFzq+AWk8rNUgQBeaPKNG+2yjXphoI/ZWvkCJLmB9LndA+OdbWXnn/KnJF3m502v02a5b7WMJAXu
EWx6PYuRtUd3muW828SK0EeOFeoVNVD80Y4FJzWDkalcI9cRH/+pgxTE+rO/Vg9rn7ojAw33oFvW
Jj3BUykkCcKHbNDcLepnwxLL9U+by4b5UgTC5U9lhiay5irWKQnUar8G9xxvPCLRzhqQ92PyarXl
x/mwFxo0yD/w1RnPCa/+siO1hUJLd8of/xS9e2P8mTCkNUU7qHJe9htjhA49eRJAp44HdXmPi1Ng
IRz+0kvKCIrxjNJ88E75PvL4hfJDhcrJ5msVWzZexTzuUMcguq8pI7m/IbFATGUSnQwvEa3r4vw+
2H0GRvlm35l4wA61VdpfrixyUfAO/TTf6YXeE0Fj4MN5EkBSWI5xuG3HRkgt4LDIAYRN8Oe20z1n
g8q6mWiJheAbExNHWzzdZp5xffs563V1BiGoUejIXOXD+o7o25AcEFXPjKGitAxT2zdUxdJ3tvQL
Iumn+mG0PmzGv3gPY6v5Yg2xKRudtiMb4Q/UkRqEGUwzflDUdMsyFwfLQGPjyk7FLBOctLrcf42T
G91Um7Jtl4kK6h1bYkqJR4zusvo5ZGWeb6G79rF+iBqQjQuoLGeqEiMqDedLFvW7OIKMhXoRdiNA
ojJonPPUTnYxSSoDleTwbxWhViMV9zYdoRi9cvtcOijo2IVWuKV9ZTNEXa6A/vJXFq3qVw/41snz
h5IausiVxmx+A5iWvgM44aIodpqHkSa8fe7/BBITkOqOr09D2cJcSIbGX+DksZeZtcBmHw7hyun6
+XEPVocwX+d9RjFfiL1ECMmBZ8dKU9dK40q5W1sP0k3tgl6HnkoCAZ0hHSqjrTDD9hPrtGILmWvv
omxHVdPdkgSQWNCv139GwpVX9NIpoiKH3cbGz8WVH9gkQkDYtniY7V3i2yp8lcp3x6W5CPoqa2r5
K/Sgo1iGKi8HumPqKECNuao/Bjg/iFkZ4lVdI+3jptWUpZMEVBV5oPIxuPnZbT0gKvaUF/wbXexG
mJ+oltF8BBqZqDoinSm7As/ik8Lx9bM3xdvlqtzHcSMX/9rr4/fd/RBHKPUz6eLRKy/0X3UVx5fa
7IAFN7V26VLO3iZcDdOvDsq75/TkqD5XCmiMZpoHIIAeRrpJZf6Z04GaxUYmfhf89syU+sf7kTh7
9sMgCFO0kCZ3lykhYs/UYlHUGesWkXmGD1sOBc8Jyk/OBnlIOQVapEzj7ds24Qw/7gbEOr+8LES4
IVpl6ZK9GSrXb6tZx1uiFhbIhqUyluXpW/SNFvBYv7RFzNGv0cMN86dR08XJllMho1/WE7s3/MDe
2fGa6A2qQ9ng+KxuLJv3+CFMuFu5Bs10aWnkA4fBqYNJN1z2Mrhm8nbOWzmGxf0mq5ot32zERJIE
ARCoLDxySuu6ETcXfFFvpy1BbADDSyAY2vBu2vtEVKBrWSxq8aOdXHGIegNw/wMhocPacylAd1fQ
/nZF6ivtqDHbdDQ90Lb4bVQmlD1+FoSwl6Zmpancp8KiR6KU4Ze+IkRM/uDf1X8I1iWgg16Nq51A
E0dv2qDp92KvHcn2EGzc+AYQZETQUTEmdHl7bHg45USdPGYOsMScIRkfCUxJtF1ylFquw9TJ6jIx
sUpU2vsNE8z3Hg3gSytrIHczE5VheqBFRu99fwt8wL/e3N5ZkyFi/tNCizNBO77iW6v6vAP6qs+5
FlflBeAnPPl3Q/RTbhkHJO6Vn8M5E9trZnzBZbJ/S6YGhTAQG6MQluwUtnrExYMqRH1rQyjBAA7H
itsTxgqTYJRES4v3o7uFX6pVy1UlcDvzftEzaNLbWiK7RjVnhxV0dUbX/E8OhNUtHEfsUVr7x91k
1X1O8+E2bv1Gahtk28WV5Mc/C2DtXSXH6cR2nKejkVuq3kpsOgVRrBSkPGYrXKFSZWx9EjEVZW9x
ak2Xrzps5041gpTtwBdUTdAybXAFwEX3sOG9gilo21TsShUI+EUE+PjMQlyLl5KtzLiIsc8gUudi
peOz8zHPkPtWC6cTdh9mBij+r8PV0k+3Q9HF8u4/41zCAuEDSbbcZsk1YktflbcDI35WfoctahO2
0ZtO3+l94J2X4XuZYusj80CdMW9uVUHZE0DTe5PyCYyXdrOvtaVpCw0Zkr5flM3ZmDUVdJUYA9Oz
v0J8jaHE6TlKfimNjXSkVudzFH9fZQauUga0VthFzjMBmn6ytF1itDksv3FjHQvZH3UuIUJ5Ywfg
p5WmTBNzuIwfBUJvM5ey4LIWt5LJoMgFGWPGlwOQhHCWU33GR5GD6REirE+umm0KdooGot3BqICn
+kaK8IHcjEdNOHEUmk2BoVNNSmBkMh/tBbdQdavEjX86WAUUSo/wNTwSmY66vXNwJL7Xar5unSiW
JwDsQWuXNW0R87UP3B6/UcdPh/lrL6Wr0AsqD+c2aiGR438i9vonJwPH7ol52DmpAKW60hiCiYE2
gs0d/+/L01JyUmM9cRwPPaDgASgYSvtPxLJSBsZSLI+2LhL3UqxBntCG0oBwYWqd7zVA2VACWVbL
PNlRD+a7e6DIv75W6IJ82SZxxbPRmY4mkEhY2AgxXGe8ux1NNdrk/ouxhPzhZ6xQzUK5gz5p6mwI
u2SCoq7Fz7HgjMBYF52/CLgdHFuTygaPTHK3oIsbmoHiQYHyk8k25IAGbqgMYfZ8O8Jar9CFX8mC
El1EOdx0DJkBX/8Td9L2N8AT7Rf2ud6zjt9hEZmLdGh+u+RfTnJrVw3BUutJtGpSzX9LpNHB27TN
tWCBc41NlvEjBasDR/H13arx4LoGU6vnVTUCmYujHUGK7xJsV9eIMalMp4evsc/cgkjm/axQ7gvI
Ek6szhVfkg+/4dRcoPIObw3COJxGUHZtrvPIz6i2784aJXzDTzKOwRMgg6VIZBQQEdjkMgDJd+lw
bJY82vbuDwW3nAJg36YGt8+du4wq8jN4ET7OuLSt5aG5aP3QQr8BrzbLnvOW/y6mIsvh9xxnrvfH
hJTKirOPa42IJ/P+cFHhe2+oXrFTPoA2ElN4/56tdBH1uregmoVGjc1oQjdzHQVwNIjE26jZsBH9
FXsCDmgIn6iicjrrOr2nhx213eR3Q2XIM8J6BALB2wFXNg2AtW1oCHDomxJO882UB64k1TEV9YBK
WSCtPHS18lfe9XR5X+xsS4/kguLiTQSxQ9fOmyhRBD4DA7pml6LGOfHCv+UU2MeM+lkmyk+97ZQV
RksKOkDQRy5tyXN0Xl7lXB+8Ro0waTXv1H5rZvjj9Pw0bx9QJEJvwFpYwI9rF4yiBMxypK2fhZhw
u0U4781YVFtbCu8R2q/vZIR3RdwjTCI58DMGsSDQfMWFcB6uXtKM/tQFKF+lz9K4ADuGUg9sdHQH
KBRG0P0BcyP1QmELda4c7UxTXxil39skBWsRYTWjI+jM4zUN1xzxs1dW4+Vj8dJh01yU/ttlFd0Y
fleYZllPu6DbyrJSM2MFx3sqj8il7KFDAFi+9Z0Hhj+noDsyR2ql/gBID/mIR3opmKv4cZiTBUpm
a6QvWo1v3WjK5zsR++3b/UVuxVlLdUm8WriAcESOwujBzQ33yOwVAidzdSc5ZPK1bjDTxp+HfjcB
leq7uOiK7AorMSUhQl0pCZH6hJETWWmxSBkOT7adGdNoYQIUYM6eadbv2g+jw12e8a2J0Z/f7vnH
EXS2tTMyqcSh5HU2wXjZuuptNfiPhrHW1GYb12UOq6EmEXaxFuYnYG4FVB10diFXwkU5ekrvkcAj
jPgic01LUdkxFZgfP02QcxmqTRJKCLqDSLyCxQeDuBCTBigCy/cX7iKN1Suz5HvIZ4NfTXpBZGc5
aczHMj2YADXROGdqXwgUBA3Yh2hqyYdQQOIxwrqsK6GplShJfwsIDHerFu2J2wSeLu7ygmaNK1ip
xCZwozjszFNIT47BJkBz8L8fn2w5/1wpX9zRFZx+MzN3Xj4izBEwTZ6O+NpUKdekNoYklFt8ayTq
nc8aYj32/32+ALAV90UjbEpQBmC2c+fOuC30xtAzIxtzYpviSUouk6HftjQz6L+hgSA2QNLRe3am
Vhe38GqbbqK+lvjnHsVCLw6jheIf9PHIPCC4UelczkZQ48Dvufzx67XLW3YqcZCNX/DAXMTxTqzW
s5cH1ugwtbdfh+GjaBTBI80HSEYIQKhXzBOqR94NWfHSQeZpHz2ZFZ3i7QBCsOF+0og1o9qNvXEs
jR0d4P7ayloTYCCztS4UicjI/wCStm4BO2JM7CxRBYegb6gG6hT4RHtqf0Ww2ldgqz2LCUgbSF8C
HMhRM3oRjTRlar54Mbojxb1xikiJvKoCJ9j81UZvkbK4y8nE0GhatXsSnT6Fb2AHSA6d2cGOZiWp
h3BQO6CNdTT0r0Y1gZNOVTz7trwpbXRds0+mhWUXoH2nqqJmv3qNMiE74WtP6p+fl7YLxSgrW7NS
A4JMVYrvEJXWuoTCc2NtCNsu1CxrAgZraRtOE1/zq//JvaWApoJyYyIIazYcPkXnz3FxAztMHJdb
leztvIQs2EUFZNYZ+zziGyMnyKUl+esHKhHqTjijqU2txYyUTMfsnpONxrUlROvc/nKqXGtlscFe
2X485oSxrEZbLOJcEAsSPcD9bFc38jWvmPur5lzb8k9aRTIn0Gaf1RuTef74CJqiu6rR29MHu3S+
AdthcCJhHiYCm3MbTenaGVRQoXTlOkj6acFxEKZb68ZMdstukaHKZ7J6dDAJe4vBDd/wW0es7Sz4
C0Hb8IO3p6nk9s2DNZINXY4lB5oZ3Hjuv0hCx8eo4YPLDTZA92qD2HZY91ooJoCQY27qItWHApPZ
W86uE34UrSuZCsH3AkHLQJ5Db+DvNXJBVp7Oblb+qWdwZ0Zw3wOrMRAoJi2ABx+ztE7TOkuVQuXX
EbkRvFIf5eo5crfeG5X51+dzsMRPQhvmvW8IDH/5wBykmdlSCGsdKY/yY9vqcwttbuY8Vsh6Zf3H
ryrXREmBKp5Bb9P3Xn2PnyRPxYfmJ8UKfOkoBaSN9+E3STFMtb9KvA1jp26nOLWN1LPMAbTOs5QM
QrM0h4h3fdlyZSs06js7vtRFKyb4f4Ni67bNJkMm+YoPpkfrk+pUfbY8DRf3aBq0wAZgWDJ0b1sU
6dbwOPUV4P6VObAd/k8WAxl2C/UcmKRA50NQG0pcy9dT92zJ3h2KrgAC0dz1li6V88wwK9idkr/6
IWGeUNuXFTgZNvLLFfKFm/MEXhk+c6hxL4dStCfc2U0D+hkvuytiE6bqDM03X4UGUC8lMGHWoxRe
fXlk+b4FU2EGeMVbBq0Nqkq7oi9FLz+D/NK86+SNg9T3QSBPhfG+yFLnqdvDlvgiMAOt0lDw6UFy
i1Gm5EcyACpZZ1CGjUY28W1MwoUIk4EpuNcgBu8dQ0sKwkGWOiOvCEvSXP9+CA+F5scqlIUkWXmo
ffxxAtzy+2zdOLNQwlgX4CtRE2hyVtlf89uDnAwMyW3xY5VYcnK+EVR79PVrPVZWAS+OFXycCxRP
0ICG/PzYrICZUMg137+CJ2PB17hd9guFeN96QsuRurv118EFp378sraHIIdCG4Qj6gwHPzKZHtwT
mCjAX56qzqJjT4oyQhz/7tAYAy7xCoOcfsTUIZECbRMqEkQ5FhwBgbvFmwM6zMR08aQpaeJqU7HB
siVnD9cNPwgHzV884+ubJv6/t8FiIXxOCZ/isgDHMEGlf2riioWzqerF82EJD8Xlyyb/5JDYX4cE
EP7UoGtgRVfscfFGdTiAJR6sOKEqE7y5Cy7TUQA2iaCKodbg/pyqb5R+aywapMpSXGqKUbM2ugGg
rMo2cvFzC9JGXXbDC+8JuFJWaj3HOZeG5yt89yfWqjY6iLQGKIc3hQQsrV2mXTvL2JmV6xPEkrmd
fWImFN28LIamvRwmXvCHb1zTmbZSoJ/UDiqxt3SEfg4ljfkzb/FtBcOMjYZThgFPiqAwLQXBRi43
N+F70d4/qOhd0tKfX8uDwgquo5hbyYwmPLyFihQxpKuZnM14YpYvv85PztecJ91sArkelaJd6p1l
Y7EojD9bZABgV+vlumh4pOn2mQXTKW4F/6Xz0/I2pHQN1jPQjKERkl+UUltS1sbL6TbNJtgL38St
qFtpAomhcCo0bz6Q5hFQ6QA/y4o10DWys6X6IH16K4QkgIWwDZ2BNGS4jhq968XN6zIXH4QaVSUR
wVpL/Vay6UFeaZa6kYmv8KWXar86OWhor1ugFApAbiFrCt4E61PNmih4XxDubAT48+oq7mmkpLzr
t0Apj2/8jcgfyAwgYPjNp/rhCwXQ8Z/myTCwp79EJdvI08nf2OFOCiQQ7V/y9FQYLC68rZHsDM4m
zjO2/VGjwHtsj3NKU2uFwswX6gjRKYZWCbJkPL80BT63FDx6XpZd05zEyWQ2hP6EPw4i8euKe2Zg
C/uKl/paaBaL4lgdUUAJUXZtWWpwHWBYYw38ZaB6I7GftAujnHsziAV3PjP9EjNLzYxVGMu7jDu8
oMfdS1iC2mghvFDHa1TfKlu19QJYeYO/f8/vUia0VyELtNcl99oyyggFRFOrp7Pl8NDJpSj6rCNt
vfZfE+w0J1Z+VZV4xwPXSsliz57iTKJY174dBeepMaK5iC6L76Zix6PYcyfkMPkZoZZGGqcZQMk/
6DqWLk4MvcSvOGhNzOU7oHzpppuedsoAXF7jFc7wWDLKLj+Ji9ulLnqTKM1n/IikMt4YIvHfp6f0
Sl3K9Q+GyRO7fjJaAbnGOMzxWKpgd733itjfSzPNKUo1SVgIEJ49LZXk1UHk6qrb9AvPs/enqMkw
QcYplyCZuQnGKitcxMQJhx7FJwTGScos3EqLVdcFiDWzwSixEs6Q99fGLOaZh/fS8lBD9M4LbsBL
Et0aAr/qmILo4aX5aY8/c2/mlC9AvVzp1hqNb1nFIk45a+zwjVjNqkTESf5Ht9HQ50h5GYdUZj22
Jw5eZX8OdtggW4DrerWx6YDwQEGXfLqYzw9h6vyN5CDxlWaPxQiiwJAoie6BKHQ7xkPD3+WQTax2
tsDqMj/BJrlr2zjyZcdG+rnDM2f1wu/AMNLwU6O7dRxrf2BHwiokW5pmfGAE8DYs8P2VZeVS1UVO
51OVkSOYvY2eczzNdBVD1gCSbZUTSp2PnP5jSJNIUAujczZIG0t0xD2QPEScUh00ndi5zkR6MBo+
t01sfezFv2tuAW+XinumyXgOBFSVARJwKuvG3o+3uj+6/oGqqNe77StZwjeUxm/MolBSOjwjWP8x
xmWS80qNdoJPKmT/qRxFtC+y9QDpzVkdD0SpNo73Bxg+siBSVeQWkmlD9/2jMqxH8hZOWXF6oknf
MzVyFwGx4NNQzMpiKMuEwdpTJ4dhn3ap0dECqKg9PkTsOC4fM7Ufsf0xjpRlyTUS2uncnwXx449D
gesu58jOFmYpYvvIBu61I8akewBl7Cpqlv2g1GEpVwdCVmlYtJT7eYdui1dYepeGr2pi9bFWDi6s
6C74wVZNJchU4U9g/HesRuXtPOiYnX4lS5VJXXG3FF1tQ+wMpkUncNBYpe66vkl008nZ3vjD9NIP
/nrdaYVzIRKL2P4Z9zIbWw7AnUMA5BjqUaQUblqYUV/e2NqGi5CxNUOSxMB+vZNGh9sZDo3JUmJ9
zSBhODgKV/AFrHC2LGUyrCsRiU3kqQZt1M9aTWiqLZZovXzSsWbefUC2GlIq7SiYle7v6X3rFXEb
nYL+Sat9DhHfqiuIYctbyI7XtMOeNEtJhhkqleP08EVVKd81k+1verk3eqjgraQjDYqnKVs9zyR+
dcIpz0O/M0LZX99ZfeQfQ7UxZtdB+s3+/uku27sdXnAX6TakGTuZhKdS3ZDMbpEyhqCVnaEdSSGz
dnXmE0TGW7zvculqMxUbJVuRR0PnPNv9M+u9wgXIvlDPNP9wd8RJo/HGjTKnNp362RpOL7tYyI13
7i0M2uPeKHYymvMgn/RJtH+WJDqV0qnMYkkJhcOKtKCa9shz6RS0DtYYHuKDdIw3DztpR+GCqSsY
L6GmLB4BkAEzIe2AZ6oV0qwwSEltyoxrdrMK9cvH0iU5eHQLFgCDjY14hSDVTkpbZoIYIDTvhkAw
kT1KNP8OvYRTqBggR1G4t/splB6q+Ro+s6ZYlZdNNi79BHo2lt/VvR9ogriFtSFn7PckEwPcqgmr
iwez2nPc0nv6BA3IoH7wLiaKXg9z9iT1mJUMuPqSzrHsjKGIaDJv8OfLJ789pq4yZkChKWUtWcVp
Egq+pfIXIqSjclvm56GA5yqNdxI25uQMyeDuWsMd+RPnlhoWzRYdgFImP3jy7IAiU3KqvgmcwDnp
4UyyRh6O0KGqrpSQ8XOvtMamMVov6tS6AYx0Sz1dnnPbHNPbBWUYlyClrt0Bj67bpFSshvNaViQ6
7SA5kIXcGN3225ieL57RxqANyOIbm3PMv5Apgv30PGV1nPl0MGBWQp3t335WQ3eJg2rG1InTnrW1
PYVD2QnKWpgu9uyg0t5ywB2bHNWD9XFIlky+vKZiwhXJwyHwFAEoA+bfTINmCuSEmmj67K00zqFB
Co8TczwO+0M3QT+kjuMCXo9CJJDErYyP0+mA4qLI77Bs2W98xwM+EbPVhVlaGR9taXn1xylQMunl
dYPrzfyHn3WPLK9T4YK9iYVPHc8MntzyR6wjP9WjUCf5NZgwIf9sEZ/h/6TpFauYWhBXzQBb/rwK
P4UbdEcsZQ5ikGuZtnqe5/GvyULn6LQRLs7wRFLGIb1lxdUU4SRfPK73cm/vwPyuzAwRYG02/T1c
eKJKPK6FmEalhboY0QCmwsMgaZ6QVhmypL2h27O8F2o1GcWBWaR+NMg/JIExYxYNoYcb4NyYVXik
1QpTabrtvMWUb5fzM71TpFL60anz80R8/3k9J+N6TjbGjwDrZj5NJ4B8PUCGizNHFuwRorJN7d6W
JG0R3j6e3licJ9jm0VL4qIwDNDh0j6W1EqOPuom2gRJew0VGazbML0XtqyNuN4rVkh8jkwoIYnXB
OechT/adYTPtDFkmbgZfVAW8tRSkKWOTA0PJw3RXVhSKcPnIL2G4ay3G1/HLINqWm47LGQsjSBnj
G3gfeFrYJdOVOPUBe626PYRjr4wfcWn7fmH4fopPd3fJRNkx5uSmPWk5pGNRqXMbKcAE9XaroXL/
JVS3ZmofyFWhpj1ybQnwVENiqr0U8zAUDETOmX2GZvyUTBkCLcmDZ7cSNpnaQq4PTNrSm1qIU1f2
ZWOLRXufKyOpK+onmUt8Qf6lzd/871Dou4H2XbcZLjaAxk4Agc6nMd+AR8B11qD/QphrqLpOQCol
axnmySVcCnK7tRkSmP3KcgG9a/GguXc9TuOSvj9wExr+w1ThYO6HESK9IzCiQPDislSC7wI4lYLS
mU+SqgvlT+1dvHM4CD1YUKJe/RJtdcCfG2kHDjgWgzx7imAr45Gz+ALOExErlp6zfXpi+neregyY
4fs0Ro/ba1wlwKArGrgXC4copS9OZfIuGEzKz3SbqtOQ34rda9eSyZblk/ze+sT9m9B4jnl5pz43
oh1G265dMH/2SvfIlV9fRFRpL49cHyqmV96Ads0yVQA2YzMLgQCS8w0gKaDBqeXOCgon4ppqiUNJ
66nepto7+aRi24QgyvPBJxoBXA2NWIvs5qLGXOj0rRx3W6CzD/rcedYHTjbmXtVUuOTCwPbzfR1B
+AyJoE9uIBHFYwMc2w0Fca4f80FuhdZI0EW8b5GOlM98AFfF+AZgAjV1IXC1DQeBIsi7poe1p7TC
SdKtZDgWRTMWSbXhf1FDTQYp04bBfJE0RegsmywYlL51v4tiaNWf2VRVdo11Zj3l1Rb3W4cVDW/4
weWkP9T2soFSnO7pO6jcXXOmJSyuA0q6IRcHamwo+P5JYV3lzPf01ej73OE1jZAckYRWJLcpINt5
RIaCnl9p5lGpMKmQZKvjU25Ej3AQzlyOBKdvyt2qwd9nL3SW2auGqa8HsfqzowmzSFMgXxEyQRFc
c7Yvzmi3tKpXkpsOGW8b1xljuvlwPJu8Z3QbR3lCdtTs0X+qQOkUfWCHQVOvKBGHeTezE9XRvDbY
2eubWJbRhrJ2pVFHb0kzA+ifnJWY2/Kj2z2aDUF85h3ac3pUDIjKTTtj1e1ybnCRqMlhHRikUWlc
H6AhQ25Dno3PCTB6TDpCIUq+7j98PgDJ2h69/EDe6wWsrnkMCKxu8qY6cDcThFernfzepWhPP8Av
iSm8z+VJAWailV2dJyca6qXAN9I6mjhkzAv5YsLvIGL6OfKZ47oKRGccT++FUr2Q3+IQ8ibYPOVS
QSkxMFhWJhhx9LPZpf3d/+KrAZ9HkSyW/tgdyDT0QXh5KN1+hwzP2gxT7IBEG2AjVMP2nJFHJBZK
urNax8fuZxlznCGS6HaihZOmejenKMaYolUrG7EOcJJ9vNkqLplWDq6qfW18NiE5ZLIj4lNYJFOq
JuuL5dCX9a4M2jLOOBoF9Ap23L3EvMlmyD/r41PrRwHup6OZRhMV/OS6N9t0XsB1QSI3YTU07zEX
pfGNFzYZq58s8N+UgR4T6PUEvHYZ7GEuO+FGv4pkU6pAqQisOqBA6njzzGHQBTXOGHIe1Er+FsHk
DOs8OO72ZZeQEqHRhsvSwPP/4wsz9a2gNDEQb3jLQqPWdEUE3DjfsRP/9Ya/2vTnwFrhe91CvWTX
nhn38CElgD9aq38VS/GGH2Ebhu7j0qSBWj1HD24LIJ9Oyno0xApQzgtxkspbt04lgeSSZRsk6a+a
NNZWrJbPV2+7PGoCjkuK1+DOa1RZsQXK07WeyGzZ9PCIJ/fCf5Vd0Bo9nqtmblGGtvm8a7W04znU
cmXPa++u0yWePkl7b9VwS6O4sFq/8nPBqtK2TMB4UVvw37Qcz16FesTVJ5BMwddk8kKJBv2F88J2
P+RKU1irKttvRcaW9XLMy80xeGYeVqchMNQZuhG5qMMno62R6q71YiljwtUzxSS2kV0qHZKydkwg
NCTi0xbOMf0cu915LKamgECRrPdEfz8wOSsLP3gGF34TjyOphFR9DmhHCIGAuQ0Sw/BI/hXYBmCK
S1pqtg1jvsp5cUDXRZNCmpHzXYZSlZrUM0bWF2N4OcZQB/1dgMes5V6fvOuetcY8tSIM4+3dVljr
QjE6DJXsBNka0MGVdLi7LRBXPUNp2Z7p/upBGkE8Q/DKJlWQqmvKGk/kPDHrysH8N0k/+6bAoLgZ
VBMcYV3tyu+I5t/tF3oRA/ZB8E0UVgDwd3pZKxlaCbICCETmyVe8bY5E4OqCJi3Fvrtb6jU00iWU
VWYTPRWIr1w40YFshRWjo959RWlBZt66QLBZyfb9aJ5lOD2vOjkZ8eiuGvuSjESlEP/7AS1caxJU
Wm4svIRZmV0y021C0EHZlCMNF8xlWt2CGvUr7G+Z6nfmip9uFnlMhNk7eMwAz6Pj/01YKvLjPLBV
k4Q6CqUZKG/Z5O76roJpdyjzR8gA6VX6Sl36sh2xL/KVNnYCc35qI/Bd1tv3dz0WzdvQtc0p3Mp2
QTn760WpA2E+QlCHyg3RgOKhbsWoUoBSPhCMB/ReOWmv6HW+rblIz22LWtpZbHymKFQGpORKXUnB
g2klixD4TzfTBt/wIVcw4iObHWtr1OmwGTvfHA4WWPweUjPSazMWkDEplcqxy9wyMYQj3AwZ6Vqv
H0nrIUwRZ/dD8JhmH1KnheARc9NMhfXFx4QwKYh6J0q/O0zQbigk6/KqluMYKRF6K26+lkucbK0a
MlPLZ/sSOMQBgWRLHYLch0rHUNB645vB2szogSNyYoh+ER95D8w0I6gbVIxXQZczjHTi0nyMkjiJ
r13YWDcUtvhigsp/rLb+H5Ntk9z94ogLGt/oT3FXLYx/DNO1wYia+QFhhaNpR2Sq5eQ1S+rajIge
leH1pdFdyMI/bsFrfe+haq+CWYb3OVQslHePeHNmYf9pgTzSf2wU7mEJzDeoxUWKUlTgdmJvKl8G
QoNPfTlOE85wy5e+EN0iyG6oYOp/4K3TBnH8EhqbBX22U/youHVBN12jEj4M/J4dStAYolPvyURs
hGbs1gGraIbEdz52CGhhSdISlAVTRYS7UO8eOWrfErkIlTGMoc0mE9KJS7wlj8+bQoUNvsvsEUrx
Plq3mDuTyaImWgsG2+h+3/QKDB28GnEnvQJ3mFfbFWJygw1ZAvp/BkBAom/NG2Z3Nkl8X7adhpns
nua6arDMBAI/CBVwknG4Ley5qpM5Srd1QXWOLaVdMKcvW0qTKbT9rEh1CPP1/+uzm5RNHqLAHkcT
qdHXz5pWMi0xXsBtqKm2OKyFNI7MWWYCtWl2gzzc60mrkcmwtcRXHmtNZDGtlLtX+Ax+9214f88P
4SZKkgTmzmWf4QLX3prEWKOjn6AcF8FWxxi4+3UjFoQSEU8ezUqqQ4oFJElLuIlPgIv01J9Y/xhe
vsT9KAOcFN3EakM7463QF9XFfv1+ZxzFBPla28Jcgk+EhFJLXn94suBLKmUt/JXA31wxhf/mbdaO
Sl1aLWk77yxSs1HqyUhaNQrsm14/6P02WhhEcnMSAVfJcPAeMY7TLfdg77uVmJNm/TX4uI3P92tK
s8hS5UMR8mSJW5GkyP49BoLi+gDrQaJEEWL/1/73uz3hVItLLeRHIHTKJnDtBlzitzRxp65Jr46j
14H/qVdpEXneElXgfK7qvpCfyomozENuN25p3r9A2kiIGoMRP2CYV1XPClfDBJXi4EdWJcD1e+7q
egm6by5+jRZeL2ZqWVCoq3TUJrSr7pFTvlWqaBVJL520Ej5JnerxeMwLF+Z7tTlR5qEs/46SVf2n
rfR0MmwIYQVxyQTN3XLibiJiporGcrWa5kQtEEYBUdFl7mX/fK0dmfyirDM7jmiqxbGPpHpYmvw3
EZcCnzgBcxNkv6SOMM9pyWVlSNqKagu6N80sJuXS2rH0pVH9vtPfQJXLbRiuODKHT3zvSDnouzR+
XiAxzjbL1dN0XEfPYJBSjVVSiWf6j6nUEvvErCSJ0Ggz6YQ2zspAZ35mhbtLjkzUW3ZoNoIg8Jra
+5qh+jMbNQzlHqFo73HiZd1cuPuf9pjgSug5qotxbHMc6SSp4uhj3jtrU3hxOMuD2LmhQiL4BUk7
HXEJtzzxvhYaMc1H76nsP0gUnlmFqUWu4yRGmt3YxJZoNFjohcevnk9K5ACfCcSgIQz7+rFrkGkA
fEjht3gqkWKcyyVvkiaRiXNg6E6zfeOTq3IoA8pBQ+rdkslQlgR0gAgRvVpmBA0iwSpD7IoHii+J
B4n5JqUbQ63qVMhZsjfHORonIR5SLZ6v9gKH2XEg6zb4jTrJOHP98tXatkXlxc1VB+DWW2dWXd2U
PWzxnwoP3p0MPs4AljGePkMYdEOxGEC2EsHS5WKf5SEPO9bqYsiG439dpeyeeW4HjQk5U92uzP7U
mkj3d8xc4W4GzJOB66TSFn4dn7NKhvxTPedrw19uHXAUwgInZjhOOXT2EvbmH1E2l2qdopohm/QZ
8fKKURaZt0V95SKS6iUXYEMiHEstZrFmg9yC+3mhwSkkIa5Av8UOrvI7DvNdB2nT3NjpYNO5aKHd
i/l8yjHSIebDvzQrTQtWn0aulnze3UuVcrOGYoUpHOmG4kVQzGag15rVYwHIIbxRO+1Vz3JabW8j
Xf2a0MACV0+eo1BeTBbPyRF9Iy/XQ77wIWsIn95m6b7tQId9zg2uMzCMQNY9zV1mm7jqtXiWPCGU
ay2ZkYLkiitS2cKj9O5Z/Ssz2M5fMA1XXFFL7iP9vI3S0WjmzBQqFziUU6jWrjClVJdfCoqbhXmu
ZUOyfTLYKQY1SZcKdJ6KoRCthRNE8hITfMM8mOriK+Dw7he1Xef3VQSx/b7lBPrS0oXu4QxYWQUR
/9ZupdrCycTZS4eHmFSuoCdufmU7lw8tBbS3PkB4giy7QFCNBU97VgePf1wty43v9iAn9CzeTWgu
2p1JoKAXpC0Y8lD4sp8Wp/0tm6FoPAIGOYPo+dr3vcQ5omy1/ute5ruAftRW2rWReC+Vb6pvNKkh
9F4cxSJDQixno6v2nBoRC6J/0TfUsoIKCoD1HkrZy8UBiMGzgw/KZquVDF7BHp54yh2k2a5mqrYx
exzBCtnU+Zaa5vObORvihJD87l1Q3fMNmlp4DtIsDdTQrsYBKJM/OcCNhve1PmnkcEuVJjJ/zFuf
tWYi7FNSemVP8jX4ydChz/keB2xsIPRtKet+LWYz+7WwNF7JN37FDbype9fqh+w+9EZxtntR36LF
3iJ7OEyt4gbnGzKEcTVryYF/chptwIn4TRfJvnGRWoMt6tuisc7cQR7dUBzAftLuBn/+1TMaBQuW
RIEFsYm2f2G3v3xw08Llp6bc/Fhqi2yOzaGz/8seD6GfLAGqWRfDhi4OFGyLVB3NGu3PtfcqsK98
lAeyGtYXNW+psUMIgldGTbZoMvSS40DWiSfb7+y8mVSrCIl6vIQfJ//rHOPj1lMRxNFzAmtJxyh7
DpEyc/qEDaxVOXE8aU3NACk4RQ3yvoah2ExT0J2AWEFNIOH/5huEBd9iLeXQO5Z87KvxpFe7+lkg
zC4lEr3QveMIXUuXev1HifeSusIxA/dyawIRWKZEBzNLt/775jWi/zX6NofgYYdaMh/9NAqTyvPc
dxLqurcA90Kq3as8lvyDehKqsQzBNE53gKJarS913CxNFP8nAIUQX8O8zra4r9zaezqd8xhrRgYK
qw7Spbte4pb9OPKfUcL/UIS3nXO0Cg0/o87UV3PtTEwHrY4Pm3U4YWXM2rHY+RTg42tY71ryfxhV
QHxde7PAuXkL6PQENcwDGk3JhUdi87o1T84mol7jh5qsjlw/Fvoz6lBQW7YHORTeq8rtxOCNFQYF
3CwAHr1WjBjFxQWNbi8cwBtnKjYZSm2I98yE7QIhpfxcsIVSm4l2dUtLs+V2nHqrs6NQjs/0C/69
Hy6L2YTRhw15+LFeUaVllipxHw7IW4JmTvlZwLlXCYPaPvSCZcL3es7OQqVQYfavDD4IYiojp+mo
W7SIGtiub3z3WraXsSEgeU0FF8FLvmXZdAbCsPEgg8QNw6G1evgPPFxc54FUkhegHxqoig+VnyiQ
EQbt7UfbqcZE56q9sR+y/fJ2fnM2Mq20C7GmeVyLTEmxxXowoZiCfp24BK/kt5MLWMh4+G4QTev/
joICsAImAsXqoRqJmEWIQB4ZYJuhPPQEmQ/wVaPj2RL8jGUXsK9sZizWeVl3cGPsl4nVRRvbM5UX
iMzGf6I72yRaa+FQb163x8wU7NOxutymYeGNc2eMH+nLMN4mlR3aMDgqsolX9XkpuWNFU+tWX11y
che7FbNfZ/oUDtCS+57fPHapp6FBGyvVcluzXCd+wTATN22i/oiicQXU23pRfKnxyT06pACs5Yqj
VX5vFXvYuYzNfFVj+eNKGegZ+QV7mmsfg8DPztHg3Jf/TvLRKG8UHBI2I6r5tsKbHrKM9MwjdWqk
7qa6SSUfBtLk4dRPxMsazqzdgW84Wg/Vica1h1vk+EzL0RKfpxtDjoKH/TOMsRL2uQGiWNYGkQWY
DUfNDjE9c1OFdvkkS6sWk1L6ONFuJkvddRzH1O4bwDbkKZEBtnMr2eEX6rmY9/Bo42uEeNcIDTMc
qnrmoL7QqUeNOJmlrYV0LcpKwZN2fcJgIDZMgNhX7qjjdM2A7c+Q4W10Sc/AblpuHsEwsQp4J5bd
znT/JquAiSnIUeYYGwIVYnUKQZmitEVwpnky+P8ir8USxPfIfzLG8ULaHmvZrWznt52snqRWmu4p
y4Ul5+wO8d9uyyofF2osuXr2Awwr+QtVf19MoLAMJtTjWyjh7QCAkfDOKPgah7VYYUjMT1pUqlGc
GBUNw+2OxuYx2N96Mvioh7FZORubIMUb8sslmtC6MhWEqhkBExVqMpCrPZIJe9dT0PHTe+4NzG8p
lfT1tSypSsh77aElqQ0mt/LEsiy+nsAURZGBAvMJ07JqFubtp5AtOLVC0/g0K/dHBOFoXW3jd5vA
dGzqOkVSDEULjTX+wcZJ5csUPt+uCTDlT5jpqtfVJ/UoXaWdQjW6REKkDTaHHcwJAmSuyJolTpDl
mgTRTOFVh7Jjg7gxjsEKUAB9YuExMdofdfZ85K6mjJoEhMnIaiSbVcIYp9BX5ekEQfMsjT6tUS7w
Kz9RgqpOqbziLRj/ies1wrAjcM9DI9oW3fxurx3Pi4e9PRvIBZvnsAXGc9Qk9TjqqiJrv4zWGKpR
SuVw6i/wE0qux7JveG1tdIZZK3zpUWPetmDD8jujASRTZVw9npRPb9kSE95QvLYuy9yaIyqIummu
eXB9lID2aByrYcl7bG7hreFCdEGgbmHio3AwpPxGUl8wiN9tF/4NdF67zevA/oWMfiXCQCj2dN7O
v7nScf+SiugxYT941pG5kEKVXGUVaD9VsRPBloShioiv07r2HemBZsP406A9xrZWVkOtKdgR9JZ9
LwAfP334mhg4roF4/HPdKG/j5ngrxbOnHt9wtAKeNWyTyidUpQnwus/BGMSObzx3FgEgfRuVYgsO
lo+u4JsfEg4syATl3enDtegN8eiRUniUSdvtXATxo3GYMs9a+f491M+F6vAahaAMuzM9cDhlq3ug
Q3ice+IjQiIr2kr/6lXI6cAIx8Mf0uW6aX4gFUkEe+qG6vPFcZVfaVmLTZxwQ4AI2E97JKqLdTaq
w4BUI8tHY+fR4IL1fcF6LKqvituXDxU4ergG4omLJBeTU4ZhU2Fb+bph4c8T8sNiSBqR+bR0hSws
s29ZSBM4uGM5YMrFjP9zEmkb3OOajzbDOgO5VHsbtD/uZNzeaMu2p8NrC6Sd5FijCEcV/ILz+0Th
L0p6BWNWSZLS6/e8cIil6kz1NepK+9PsJcBN3N9ioxjxEBo+qEaiNgzlhgekJzqc56PjIMgJXvwj
nlAV6FZ+c0TBnzH83jZwu8tFYbGWNwJD6E1/u/EQoDfYttZxfVVrMj/OVd0PuGwP/4uh7MUBzjBF
xjyTzH2UC8fio4kGlvAAIZLxNYmb+a89eXycdAA2w+WlLqufpGH37IQzalvu1WLkbLpjXcSBQqs1
ATLOfXuoGQpTh4n4ALy4DZkOqG5PnVKcMNiFkhFBuPWapagGU7loUj8Kk4VHTPiT/qCvOId8HO8e
ybpgIdE4qPt7EIcuRg8wEh1tEY/4eaZVzlgao6OcC/Z66VvuLlG986x+kjWGTeyIWZjklPk/Jj5i
/mZX92YtfyMOFgh2sUyluRPx3Dvneu4TkrTu+ay4SD6EVJB8sPvWmz839gi/2UYwq65Itgv/5l2x
xKGg5XmzCExnwJk7vaVMWIVSa8pvOl8vg90w02VMJjNpuWplO0ebJK/0qWkqCKUgtsy4XN7Ns6jx
4lBR1ltKEbm61uidfs2KjLhKrUHkumAJsPiAm4Ak1RfKj/GS4cYE00qkDankV9SfZ+Kb01vCjnIo
PxAltU8P67X0zE17b6wjwOcASHXDDpB8CFk7tQCZcsV9dAj5Oablz8dtBbEd24rbnOZ0r0TaIucf
beGjtstUSQyXmNgr8fE3MQU88n/WCav4c9VCf+XUaFazupdfqCA6NM/T+088k8gfOHD19Hyw2VMS
awglpIx09rXjPWWrFdRsIP92wgtWEnw62aHvKQ2X5H8TJlLUFVYMSC024WFt7BE9XxmV/prMsstk
6m5IKaz4jarwqwXGpEuprs6eHmWgURe7hExhcoT7HHDxsixyvIQg7xoQTwuYnX7A+AkGE/ER7y6X
+MyTtfYVHupfoXTUI1JlhSSfGtsTq1PUru+3WNt74ShiDGhmLBbogBInmCog0E/3RGr3//r7zCzx
3P9fBct+qFKnLl+4zFkk/gDGm52rTV8pjPcgN6wq/lLuECGJm6FY8ZGi1uFap18CH8m1zl67tA9d
JIPX2w5qMIeUobsrrPcu2FEahn8pU0BNYR5Sv9dSYPxT6flGTcID1w7WxUXrQ0oFC4JsDjctvPdH
aWxGnQhLHK0eN3j1cF8h+dP9lYRZEG9d2vln8TQkgVQqaQcBo3A2SX5SYqTNoX5rAt0PT4LWyf8G
JDAmgpWmRdfxVNuMo5rEkL30n9aYL136JTf7GNeclQG2TzIV5U3/Id15fIcZfwyEYDGztzIlX/CV
lAWjTLcHCHXD1rmYuvVeUNnpxTjMlaeenTrCmvPNNB4uKAElmKZKqfbDtEifB7zZaAX2XVM2rxxn
1+ekzHMpq8aiKcUsUe7C0hNBhdc1XpXZ7UNqtvY88o0H/YzqWz08HJV8rNdFqzTMrlghnF3wAqTL
VpLJMujLV3UZt8jsaMIaqU3G9RvN+7UwCOiXgDm9cXqQSuMyjyABMw2QSdFm19T7/3nKWVar5MuN
WVBWyf53ZOG/pxSMAncLg5HC+0UdDfsei3ixn5f1rF7Uz+CDpxjNnKJhfqc28kKJ9L9NDfb9tA1G
rNffvlRJSc952UDoLZiSHf1R935zaPc+DdCOVd8bFPwELZSlRAlshHywqEb5NSKpz4j+EngF0Hhm
EW9wBBfSML/UIjAaPfNtbjcBnsLI9Bw+6Q7iV4HkPDWNZTXzsrd77dSuwq0cinHGGNval9XRdEJ2
XpNsP2ApWzCuvh2graEg2mS1VYgxplQR0YTLDLGAZHZQJa7D1TkPczcc3xW1G0+8dz+8cOzFEO1/
afYJ1P4nbjFz9r66TrZyaOAtEaL9n1gwMtcu+KWK8SXpKa6L8xdS3I8nnAik7a9ThCnpWSH3wYjk
JiOdOrbM9li+If0Ltf/yAr8rGO548fWbgDRn5fUboCyURTUYSlg8FVg6p9DHOLIMaUSg8Z9Txf+2
u9yC/6yVHYu2otuhWRRXhnIsgHh6hGG2e7EVrS81ui21pIL8pyPuTfZ+psrTaRi/5fdSGjdNJ2s1
StuLTC00nTVZ3v1NQvCePN7GIFuUDhQTBtmVVGoNWWpxE9f1MsI3Ereg0CUrr7LvbhPC5WAVCpjA
RydnMxz8bP9ANYPN0cpD+1Eyu53VlMUAmFRHASBaHUTFwCFV81s01j5qYFQJG4914I9NC3wTRlUn
W3xp5uOoAT+c4DBOx0YPNm33Cp9v4oMhJrtOzeSlkkkqN7o8J9uQii5i7wKLiE7CGm7avzOXSeSw
EmW684iKXUFt+Xo46IChxrferDkxrJpDf2URGNcgFd4lOtA6eFfBgfJLUQP+Lu0EWjJgtkQZ4oRW
INcyJR4UQQBYlxi+lbhKFViuEANh8F83B6AB02IUUIpp2PMfwq9E28tQIQTIr0nuonT9W3TmIcHG
NvDqnkqkTH+8mh8O1aLzEJGmZaxNF4OxgLXi8z7sEqNL9LbsP/SBUTUf4S4QazlR9ClAp63SeHPD
j0Y6Tg9T5BBG5QeHyV0VRSVndD0nG55qJ3ftK0txK3EaWjspCBwVA0j/FckaG9Md7pFEFqsA7kb0
YzLvArNvjdlUBbeB3hGOU+GjW0mopRh/FJJwCSTTy60f3tOftq38c36fpP6wSzc9876jJ06En+BK
phx1pXSpqCqnopoqKmKOLy1Y3Kd1+D3gQmDfYcU+0BXD0n2B4+JM+poAaDHokzwcfUy7dl4tJcBL
Q4aG/MslzXXziHhn8LKjmzIpbzxvDhx6PhVcQtvSvtR8ZTAYY0a5UWbP6DdjBET+mYF97PJ6SO6P
ncq79nUb2l2WzN0jd6SixaNx9rs+A1JvRUJSQYU7jYgrMlDzqDSXhwEcF6nlwbRb/3XAgSfTUfnJ
sfr/E7/zq2agOKpYWPfwa2jDI9x9jT2jNvU67UEwCTy381u+ox/IwsvshAUbSzQEuqjeTYVx8nlq
NPs/JpB6635McdJwrfuvizK/TLTilzX926ggqG5pih3l3tKgZQsy9xF8km1iQHeB5fiD1WUPsGZu
xcrJxJ4NrWP4vQY9/+//aTe8v4NkeK5ReDPZiPgFjAKrWPOttmw8VurhH4PzyX0LtCflHSj8C+vY
Eu1J5HmXP1S6mTKOSrFEuascNCGBmfcY8zeT4E98ZOAP3+1oktLqdUEcWXz52tDusM+IvGqpjXvB
4JYWd+C2Utn6CtIXT3XrA+kO7hkOyeflYhiy40mJmEVWAivG7UPoFEmq3+3JWRcnm71BSVriMIyi
qU+MNg/58xH8wWq9+cJPdrnKXoVEv7h3h043WNqgQYeJNt8rli+MggYCktXG/uwReJ1K+rNK+/H7
n2MMYPm2LBrM7AmhEE0lUno4LFyvfYAvPr2ZF5GiOSZJxqedpGAuS1KgJgFRfhv/jrYObW0DsXeQ
QsvQdiml/A9QA++g6M+XMKdEUDv8LijRqVQxsTmhkepa/QEBcOs2yrG8t7tVYzXfbIns76fEHkcI
dEXsAcY1vMgsVYqPuqyNj8DJbgs3Ld0pw3gR2xhaphXvFi0LXQat8slBB5ky/SL1eKqMEixA5lRE
zD7cf1za4C6ZiwxWB0RcqJ6G6QKvctB2KeTzB110eDbvWBfJ8XHVmZjyZF/gu2EeihTyN8jnJWPO
BdRdd+Uiitd0GHljeA96wZ3rip4q7E0lOkrdSuMXSoWNl2MEf4Vs6F8+1rk8FtTa0OcuhxXJ9RU6
innr758rajtP7CrVMqzyIGYYxU+Z7k3twxrhNvulaI0LqqetlFPk54IpVhgWr+ADIXL1bXmzzUca
BCUjo15Ly05BOCnbHSy494kCCWlRcxVwkhWiUskoVmUljVJMZDiZZJd0WJoJNTjI3JHDldxSPcy4
w32X/75nZc9vevFz6V85DYWu6sxjOqOqEkTeAjJjly35CjadcavEhjf9SnmS6Gic+m3bLXH7bGTe
Wo7Xm7Dd3GUxg2Y0BN/vecZ7Lwuer6J46LSiL8WULaJa/3PAyyaQnjfXTOIyCnH4ky6AjhSKrDiP
+RQ+dbSb6SNGJQvx3QTyitvcq+5uAK1BEJMsMlB3M4ICCrOu4obD8mfMTUNGUYKK6ox51ppcocUe
l6w4rBI5fH9HF/8fWww035FBeK0EjlYrRN0XvSteRSvR+77u3Oo2TrI1IFHCcMfHddB0XAlqkzHG
GMmY/pjO5hptfd4ix9Ql5N/bv34ImwnrU2IP+UXi/u4l9CLl3IPNTyRLgZ/fGKHMhBuB5D72jWWL
GhSJoZg4/kJ/mf0oXaSTvDy82nYkHgWwoLkFIw76tXDEqAR+u4uje9APS44ccPljFWmEk9OVO9Ql
kGDY7oPvK4FNzGM/Jbp1PXn16q5hDX1+a3NBKMREXnsKGOel84zAkTO4270Abr185xF6a+1G+Ejt
5HcY3Y7VEQDSMj24vsOiiMR5gsFrL2wNlViU1nRMxaArZJjTGuTH6Eyz0TiYSZb1js9fju+1tIFn
fttFAH/2cqvi91y/nUvOtZi3px9fBq7OFLaayYi6Lqhbs9Yz3So4hUGM8E0n2sI23NhevpXfyQRq
pVpTk/clJfro8rFhHTPtjC5N0C3HdnoRjkx3V2QL5IdVJBGpD3sruIE51VeeA9evsSRlZXknhs/0
ScpVpHyHRoROF+c78Ry7TmrzdYVf5vIutB5tptxtQ7lsHGOSb1p2l0mNs4Px7FhztyqmxFe29HGL
J65/7icneZtahKU06Dr92xXDcg5TDxFTf6o2QA7ac0y89sl72ILMUiw7l7IgT8CO7ntdPtCkKfy5
y7zm2Y4K4Azzaoa7ejvqw6Ox/xBtH9qomq9UUpUtn0lQYnSOPzc0aCvoxhBLzowG8I2UDNH6nSGF
aKDo73HJIz4z83IaHFAp7e5ufWLqXwtzJNoDdRkwlsAkSdlF1vPOqzSY6R9ffNDOSG8y+YC5qzRK
nhtdErelAsKspjgUW8C+65ud25pDqCcDGINBknb0RXuTyCbiWFHaSQEX7vU+8+W/XXjJs/dXdxtp
WRoRhm6zAGkn4vdAF5B27W24KuhsxdAdUVi7FmC4GMDclhN6rKz7mg9nTLFtgm8HG7exM3uUG5E5
WM+G3AtH0M/4nFhLcHKVpVVCxu9gcoXrCW8bdIYSmQKKuJcFXoxfENll+SP3Y2nBlSRwmQQhGXKr
Ww0f7GLz7uDo8OxGQEYLDC/jDGshu46YN7edNgKgoVk6TGLazAWesh15ZxIEQyTyR0qJFenqKLua
/9pnhpRxsSYHvDRmvz6sDZxGdIr06vk6Vk1BsYLG6dxigjRApf8zROi5FKrs2W5808FtKx/rzOwt
HFDS8tChAQ/W66HifjF7cx1vNUctaPGY4SjZkUaFdpJxaQBMB0n2zVYOq9yXR0PF1Pvi9DXnRgrI
9YplGcCJS6oIouQ1xNdnMQwJfZrYDq/NPSsjJEnv19boZteAbh4Wh9ozhwaWg6qdOKfFj8Cjeio7
O9VQsGQf8cMIXtqnyss7zWBhTq36jWz/h/8hJ/+rYv1zbLAEyIm9e2RMA3+/Pw3/ezGy7mMf4Joq
EETSaxuIs0zzvo7/qoNTPNT2/vsXtzPe5g+q4ws8dybN2gvjoLq0Eu9Y7EOfABySpY2MPS580Iom
k16TCvjHCZ3kDYTqM/uNWDIdOB/f2ugWjS1iakOM6lx46uK/YvimU7ca8jaiioEK8wWw+pWBX0nS
CsArMHYXh5q2H3vRKFpo/v/AORl5MG2+0TLIZhfwqL9anyBnCSvYvEo7dZI4HPsE0okid6SCMVNK
ZPmoLKSx3DKjefGxl9yC8jJmmcCCs/DY77D+V6vLdmZseauf4w2daSQ+1/CS1NJxGzhw6XTCcION
JOM1PF3x+UMfndVSyUbM87dLncvTsEOcVSCQqynarf4+9Xfdx9eEhMhVY/4QwmKyFoILzjEIqZat
HriQ5iGvb9X4uhXIqUFRETndnRhdbO/WxrDraYruDxc/1biIAj2bi/4d5/YqGI04mN5WS4F/rPm9
5yCKCGEFhzim0aro++jSNMH1XgzAaH+MpdWk05mdJrT0TzC3DSSBGEqWJudmEfDoRSLC6pwPE/7J
0wAMGGg5T3hbYzfPsMsBpiS/b27n/XX12FbKvR6FwMlWtotHxzNe7b79CiaHf4rKzSDEYctCBLzZ
RZEvUdCFrC7FZ6tELklijNSSw5weCT04YaT/InhvOSpaLtb2l5MIiBmVgdEjhrrvnzHhZv1zGlN/
vxdtp1bE4wpuJG7LI3gh1N9SlknjjG8cycqBGB51qhRL47Dp0E/loPJzzqi+/bUIJPZyLdbw9oU/
jZkehslboa+0TPz7F38LWWMVE7SxQywPLdsJdP1hc1ItG7VqAegp2LrQ9pIZjLSdrp1aGE+HFjjD
MJdTIJ1wyzJAQjOtgw/CEikxEWy+ZVh3le89ea9xAHNm0L88o20B7O6CFWGWFGCdGQdtLxt4wFWy
b0ufCgAp0QnSLzhpUmvl2RQDSHxNLS+DpycsCA6A2UhWBOft5gppC+BHxX2HZJ4K4L/gAtAJLcjw
NhP0MYgN6qta9Anf8Vn7I8dfPU+mW2rMMyreH3R1TxDWUx2FMj55c81yhecmTypMVfj5tWH+UK8X
HWGMAYYr23tyRHDrJ9r808Mnocvd0V6mmpLNjQaSBTljPxHq76MzXYjcRrbbXh44IS6HI1lbjIam
5WLOIjTyBLfcfFWrVp4DCjDVb89jv57XIxgbDu89vUUCUw5t+XHdSK64MsaL9MUY4uRRBo2BNq0K
GDFZGKRJBgH0ST4Jz3NLM3izK/pMRIW9fzgMj0YYe2XpghL7ZqJPtAWyWiKRgjGDEUpN4bomz1mi
UyGA57M5RVRqbb+d2TVrCtSy0jdszpxuTBsBrNphNuJufpRECohnYwCJSg7kNINKJxrZ0eLKGNf9
gPDT5zOIfXDRhrgseilHUGlwUxr4aFtAVM68Omt0CXwFgv/Wm1vZMXAXyMxDCKtq4QrIq3VXna+Q
yXmXX+BmOcKklssn/cNjDF2uGp7ZyXTzZfk70YXl1ULoB1YLU5MZa7eKZ8lwlIFQS7qk0q/jbJj/
iwmk228/+hG9m5vUVRPYT1pCXZXcUctRfQC/GITwg+C/2vpmt3XGOaOzxGzt8NqVh9rRVpfiRyAo
hdp0bS6+gSV0Q6TqQumnWItjZOb4I9Av5ODKn4aTmhwkstEkWqvzQAn9bqBOcLpJupdbXSAy48OP
0tZlf3Lwy0d2gntEAJwtMQg9dD34W7SOK76CuKUGwCpvnYDDnvznGBXHxlWL63a1ssuxstBDQA3i
NWlPvbzlnAU0Bi8SUZ/obk0g3M9Aqa7ND6/caxEL/cMaZOVlFJmXoelfb2Z2NbhcIIMSNcpz+hrQ
Yfj980f502o+pT6tR1ZrDAcRJBDp13LixwBWQSQNM5UNgu1AaPTJwTXXaZrGKqPjt9pPbN0y8LKY
fYrMe+vLjo5h04qpnzsJuyzxqeexwA6PBlz4mgW7RV8q0t7/JwGdSt1Y+yQsN0OuTK1Vz3AlWunp
uDrQg9lpX5P+T7y6N2U7kqikuh36mBJMjox276OFZaUfBu1u2C7Di5Fjxq1wErVOTm4EYMInC+hl
D9GyA+4vrgG0Wrev9Cr8HdEzoZVtIyz0alZMwfmXOb9llIrxYIaiOPgneFlwNaS6y4hO9mcR50O5
9ZKY1M+fZ5Ms9oYicvvAudITAwNQUKqXtbYhXENI4v3j9I5VKPcD4MXSYLjW1chp/4u1ucKQqVKl
lbtzIQUYXFtP2/y3xWhMF7AZK9QEfsGjTlN9909iVnNcaXNwfbUoxN/3/WWyHn8qaNgQQAJX+qdQ
b76rUtuGRTy1Q0im2UIT9fbLLOKLG0nYFm35FfC3DLjzmFs/jL5y1SuPZ1EIeR+LhP/26BNb5Or2
8okA5QxoSZPPueRsQmlicM7X7pdQ7utnrnAJ5vyu+f4Lc3FtjFTSYvvooP5uTC8Sa3aV6ZtwQ/T8
ZAEEYrTvvrKnoxt8kNvPOvasmhsfcsgy1taY/Is2u/+WPnhjvsGeQPtpvZrIh09ayGhVMfIuz9SW
9XJkUpcyP9njT4zLXcZ1EYNN/cvtbUUmG8V4m3KZaHH2WyZ4DlM3UtQlRTTR0p3U6KFyBrTyC2lS
DkH5M8u+fXcxNkaBPwjR9ZY0fKCf6jvFCnfm5rAIXKl6Ky3BuAFWIGhuO9E1I9hAWXP8PJvzIK2w
tip8Vd4yAD08Wurzwdfgw1oeKwWWRwG2C8eJefWRdKBCqLugwV6hUWw2xsQ3iKAGPXcOBak56Sif
c6FXqYehFsgw2ZqanWUnGwx5hSW3ee50mI9FRaz0kI62gWCZEk3ndXceokdifCDUk/f2OjfTVYwm
PSelxmiJAXBn9FI5JD8nkw2x/rpMzzt2VecdG2ZJF9yjxf1gTqDDAsAQxb1xu2PHUFcpENMBl7I3
AjzeR45J21anMh9ERGXWJCGi+UZ6rsFfxyZN+0NdOdcYbbHkPE0CQivvHQDjCfz42NSczhsC3KJk
ANnJIlCPzsYLlevGW8qew7QzapzzO/thMY2WA3Q3dd3ktM7YsQbDenepwQpoJJ0AL55/Iy3yZnFi
BnpU1OV9JzdV+zZtDXSiparpErPVYAzS1rqqpHEILLleF/mvX+vmHNqVBOrtKtNTVbJ/uK1UI+5R
H6yL40S8OpzHgaXOwQK7B9ghymvchpHFQda0p6ro2ho6CKFDePtoCDotC9GKofgq8Gwl7K6J+FT4
AlAWE+JHPGa6jDqWyiOSD5jNxmsGjPEQMBMDHiacItsJ0HvnGEc7dP4YGwh69sLfsmMMrbpaeJhF
yM5bDQjSAk1pBtENgAsn6haChO3O1PV15rvnB1HqSqDx+objyi+IW9wx842GyWbPv8eNU3loe/zd
98kwhyA9jwkPxklyVpdbIq3CODvMiewEo5qHDGZXBuRrjujRhLwfAmzxwe7Z1GlKlsQ2fHpGsXCU
hPv4xtQ076A0o2YF8MW9BafekHzbvSZ7ZzrOKcyiDE+T7BBJ9EwsdfLIg6B0187C2aMMUGNV7jJb
86aeRzJimmg+5/r4veT4GhWyf7lUoNGfNR22wuEC2EQajsbMgfU6Xrg/Ro4Wjs5V4Ji/v9A4Gqm6
PIrFbSNniuiqk4ikoqaowgoeKqovQ6mvoD3NueY0ZTfMmhF6Bf2DZkykhuLuWfjj5WPoPjkHrd/G
Cl8JGP0vllr1ZVAal/0AhP88sqlKGFagJVvaTxDLQZByNmB4LtKjhzRyBk3uRKAPz0G1ENXf733F
dvb9cqO7urG6InKFTUVCww3KK+BVbEFw1sFPnd5iauKG040viv1JaF89zuSuo68sBjiJH0TLZwXl
oTI6pQqjDQQF8/BXvAeeeIu4euO5sPzoEvJcxUHWVa4BO8rgG1hGCFN6De+/WZgH+zLZP9pI3ysn
8zAvbLWquER1UAyC2Me7l/hrvVn58boWT+DJaqIkH3Ale6IUNRLvoKzS1A8yo/N/MdFoWjYd+jaU
jbyj6RjPC6cuATIjvTsqFWfBvnTQ288+jKHVuMrZeuOFiBxzG/7NyD7tVPfZ4Qhkv1XNYcCHrbYM
DpzH944YbcP53YQTV3A1xyidrRyrF1R5TZyTjh591lmbqIu8aEhCb997PRVN1x/IIAviSSf97X0Y
75hXJpiQSo3c0Pj3icsGPYHRWaz65JN/QPRM0Gu2NIPQ372r710KJnaWVJ6wqo+PMH1lzH16a3Pl
5qd4PJSV5agYnpuwlaKSZtFLS77Lko6ICS4XITzVCSrQZ8NQnD9nGhSuIitfq1/C/d1vtQLJ7+/9
DWng0QRmHUpaS8SUd9IoXMNyk2ItXOkkpJkgKoDc7rBnxX4gDaiVHOCW3K2xtG4s5SdK47OpUQsw
rrehqfzrJgARxOXO/3AlbFmUzak/6RYsCKtGjE6CEFFeipBqvt7HxgSzN70qzpf+Gkc1n1ohHaA+
33jxBbUePWXmpXLcjHjSFO/g/JIOM4/ix/jxDjP5eOXpXBjEBzXM166XGBU6VHsziQVtd3AZsEvd
yRLvKaO7ChTipLM+E1UgiZiaqbjGXmK/+92SXcrsu1qHmpVplxJky7hfB9iLSlJ6ViS4o0RqyYxz
jgbwtXsXS0NeyZOc4eVlxFuh9tx4b5KG5o82u21lCzCBsU7al8lVqDEPAQfCli6WE/8FTi8XFgGG
W6VhwlvY068NAr0EZIGfygzs7RtiO2Yw89YMFqQsF2z1fdieSUoloJDouI11lbNvj9iZ8DsfLqrr
gqPkKsvMObQsqFWg9IiVh2wBA9kxY0BpCTJnvHC5zk0EIFQcidrpKrPNKVRQt79QrjqhoffJ9HdI
chsbk2WoYa0y7zcrYOQUobeh9EQT5F24VK5lEkR8tkqNwFF8qhTeTDLQbavT0AZqGjI7QvqAFbfl
mO5zib+CDsGFqmuBJ73ls1RNOiI7YnKe+ONDasyjIeHR3FfbdjXsZMymzskkRIdXuF89pfF/mIcN
wLH7HSi8UH0J8tVBegfetl/YqhIIHQHmCMLzEZentVTMfVbifKXFC/VezD3rkV8Q5OiV/ClYLeDg
2QJqj4q6QalQSuQpxfFv16YwjhKvc7wp/KfzT4TCXOe0RvlXHtX8q/oTxrl44fGwsQlkE8y2Y/H5
IS7ZoMxxdGSseVzk7s5SNMzQwoBK3/5Myyf6oIufc6Y68ivwObqDZO+PC0v63rHj2buhFyLaTuna
G1me8zMnrIbdB6PosYqqgs7BAA8RlWO83nhbwZ1TKucc4DscKcQhYY6d+jOhIyZcWmUeWEZx98bA
gDjbQU+GrDPsKHX2l30LezbsGzghdY2pg7El4jjtKLUGDdpVqTBxoGKU6S605942TW3WrwKk9HG5
3KGC+ud/zhYIIcrVwr82lvnQitaaqTtLCN6skQo4IjLKbDZ+YHxQIsa2gPIx5CmOkj4UUfmqP4mw
RiqNtmM8rjMBdp6ZOPZHU6W0IgXrH1i7JzHHZ7w6iWNynp3Ecsv0XWATAj7rFL0tlx/k5rsdLUMT
4W/ZtZjRzveW3l0g1S1Gpt3itWXvzuClN/ifStS/H01YMAICP+s2Qj9KsDESxKF2CH3xu8AhxOYk
0iyWZpiNAGmqttWRU/k9l/0h7ZRNnQNGxCc6bbjp1Ve2gy+7VvNrWWNiDhmNXEWITnWXZ2KkMA5g
pVu81pSrizuIIqrHwjSb1UYSpKEByVL/lHTPX8egzdAxVKw9y+8AZVd2WbP8wa+rWdywu2GA8cVM
1pZ+na3zNXcBYNUxnbdUU3gcjgQdJpY9FtmcPEoEZiJgbC5jfLzi6Xx/lMGvhE7SFZosvPAf9hha
wg1aZtTndU5cJlhngpwDgOCkY9Z9dcVySDOaiax5AglZCvybcXE5jXUA7Q0oL3FtHWXGmVJsLCob
LivIgrCn+jXOCYVUZq7MrJ5Uti6LxtGZbaGm3HGpDgM0RhI4hTYksZ3nBUJ8vTqG1A/0KG0j0K1r
AKMReoHXeFo/07/ZIcoJkAJmrYaEpmW744ECt8i1UmrDfVgUwJJE187tMcxj5JByCadXhfJlFt9b
G8129IVy/6BN6Uk52h3KNfZOqPURtONHxFBFFLZekWZJ22mRElnMw3Ov+yVk6AXwnamowZPsMwV6
VNRM3uhLcO3bY5LZ/OSbONutyYYGOJMAZDeDIxq7LvEEDqufawfTmlOrrdKB6URGoBGvskRFZxrb
OOTBdzVDaW65/c6FTE/haSkrb+iufsGynBTQQ7zWieQ9nnRlE/9a+MOUqF3GclF66EropNJkWLJX
KeZF2DojeexGPc9kwfegbMYmCOUBs7adE2mBMWHY9Hv9PDfqXaGz99TvMYZ2h9nqdzWISQ5JEwDH
AvGcgn5vHSOsbKcAgWGt5bif2XNut2n2ZvpSxgMdEHNrPVDLJG1+AxZ5n+Z6OWG1Z/0iqFbtL1ey
leqQpcVHdE8BQ48KRyzitkfdgyYwr3ukhG4mA3ikZcY9t40yjHcEFUJokPSTs9HBEKu8NW0LRAgF
ZBRxOhQzYK/8jgp91RqJXa9HtsFpdGLR+ZMgDJDv8S9WZYtOH1AHAxZIVKwHEn/kXSEhgUDtzbT/
vz/uC7CkyItqZuCSXzgp7PcC7deYDxH0plEeG8fbW3ahMqbEo64jBLP5rIsWb1FDl0LfR/wa1vzt
wIzQ87QiQwPhCRSFEu9aI+2wJgVfq9+6VHdWVM6U9Im90ytwUofxlWXS3zcx5HBmSA2inijw17J3
nPdt8SzLArV8Y7BE8peVhv3Ywf9ajRVV5EnSGI5UqLi2+lnUgKlGOJAnoGEdLKSMcERR/G6/laVb
i/VWkacLIdXxvHyHbN09SWtT6PZPEkvQEk4Z3AO9UL5OmujVyuCPxK6DStIRX2J3ZOWbVQ8b2BEC
12QF3lKd0rgWF2Ga6oEUf5DEWpNm670IqpEIdSZ6bavNTIJ6uetNSsBU8cvPN6incmeCBG7zdhMG
QwACtnc1GneLmSgaPxdu72FVW2PuxkZQsv4ErR6Q3LzWWQds7crk0UkoXTVlF3q++Jc1ULRBUB4O
jnW8wvI6y8QyTd5tPaoQ/Ct5s1p1N+mNAbzqMMP0TK/8ZN67QWIfjHHhmAy2ayDvIi8moCqx62m/
8fg6WIagFfW/PfRGpal1Tjd2+wYrDA0796Zxio9gV/fY8/xfgbEZ6XpiXiJ1vTXird0/Fl6Oaf6k
6ST9wynIrQIVQnApysvN+8tcB6uUd6aqnxOY/ORQUKcJN8/jU31jlvU2EGRh3lUphfLpoedX9/GS
JRSkb/uNBCmAlcg5Sltp8A253btbs0eAN/VvP/bQ1KzD1lCVihidR5YsJjtQJulJ559xnEZuzeiL
e+TlZvVymWUhSx10XZnM33+9nxtkQRPE1Yul+2TKSG371BxHuPktceTyyxtvUYDvoCPqo1K3yyfW
j+Zd+M0QqwMpcp1X0KXp0dNoanuLoxBJhlbv6PlhgoucV97jAft6LlKRhC4jodRk7c1aXCYfemsR
dqJGsvIwP/GxgV2a2BEYUZeslU8wcWfpdusacbD2t5qLVzBbd2P5EVaBAXKR283iwS8AssQhgjS9
Un3Tti3XgEKZtyca7h2gDELoONic43qTrRGt+kWRDuDiJbiEqH30PBkCBDySgS/IoN+jgZDrRn2D
ElXTmAPOoe/KWJsIFz9lXdjWRw5BhsMswNTE3jeJYgqMcC7ocC0SH8qI/of5s2kikdSHsDd+SI7k
nQOLngg8fjR9hHN0OUxDdCuUo25CDr7zbDmc+XBTmQcPxZrKVYo6hDl4myBZZ9u2o9ThlA/s/GSz
K4k1sGwZeSctAPAntrWNayFVWgmNrlnxJ4Ehj59S4ho5pcolDWgIjZb0vRnyMCYQVJ4RT9L+2Xmh
hJU0yR7RW/W7tizut8536zpxJR+Nf8FKCouYZFdUN2gBYV3jcGvzEvzls/Qv+P/dOTZ01bfgod+L
JYbNvl+H8N46ESzi1Sy+N8CyXpmVuNYr6T9RtNTvuI9rQc+S83l2OToJ95ayxGYplczVQbglRY+w
4nYDDTajzVgD2QN9ZTghfXmH0tqjV7hbaqLoYb2x1Gf5epm54CWDs8vPdSvUuLb9UPoChODRsY5f
1OPV/NRpV0prK+lzShClMlE8NNJOR0TIWBMYe31XXZ8KL7j+WxV8M4wUht3mruq9rx28Pwe3SIE3
CqKw+9x0HMHEVx9vK8x+L1bk7LeKvWi+YGD3aigZPZRqlkCNKbGkRW/KOUg5y6dvlqs8PVVRcQpA
Mi0nVzpcHZOB2s8wxXEW+IGSwTAL7rZRy6wZcYC5LPLaBNLgq+phY8l2NwmbVsRHoY8MYAfvEQNR
j+kCvgdpfPl1Y+XFidcbyxgZzqhLvVK/pd3wEk9Mm2tpMvWqs5ntRUSt/KBYEGpG/4RwAN+99h/D
Ezpq+UQFKyijzvgDg80IZFDGeaD2JTvNW67uYfn5j71lq/yksDoM1R2F2m4e8MU+9Zl1XFV3c1xb
vkq4cUKzojgp3LGCCcJRIqgCJ9qrbDOHVyAtKcru5lAcwRF/7xRecI+5gZb8nsb5cC0teePucGS3
ca7DQnMJeObvdVwMIEzzUovEc8TYRtRkYIvzlm+LmCv9aQzFlRWOeDtWgZbM+Hmz9/bLwhISv/fN
HvuTMMhtTiqgR6yFQXYSiDGuZCPP+YpoBkBZa/HvQzk+8ear27HrgNxTUHB8G2hMPdmetax/bcNL
Xp2dTwoitJk5PALjFAJN9IATMaCsPRVBBc+NAIxm+cZHk+z8gJCXfmBRgRAm8JLmG1ZRCfbzd21O
21ONZkTNSkcxEGLN+Rlebf4N473UsVAxALPVIf1pXEZ7LdN/lbXiQmyyGWtqT+U8Q6ERzOSP8KY5
y3jyy1xvZ8hgg4+1riK5BrU44nAOR5UtqCfXQ2wsMliH2bGxho7/sDlINmxSWyPIMPPldYbFIi4I
HNBh7n+9PkTTMKwP+5Dow+cmmLL2VlGZndjz5NqNAhYWEVthwsFX1QVCadiwd3/q+9tjM3nQcnee
GGLr6Adfa7jzuGS5M45iRB8+5HvhiZlfjRro+srGQ0hF7Zh4BD8D5nsvOrGizyM7A9xZpkRYPE0N
HrwxcEHjEwxLtnrkvlK10gj4TQRvst0TMgiVCcnRv4GLBrdeiv0dyW8fHUoJeJmX7YJtlPpRNbTF
e5RFeX90xwYW1FS5LlmmDMHZYzABM9wePAiPkTUhGWqsVy+pXiubdNKFlo62TQHFM/9npHswAuph
Gqozl0cyTKa7kFes/Gy139aSIvA3o85xraZc7TmwbaHgw9oJZZNxZFJhTVTLf9zquJRMWWM1MaF8
uIpjTejnM6K2r/zM+M2pE/U9HYC0eea9Url9uy31NJ6YDrbgwqxSgYXyM5AtCk6BwCVU+JIY3y1R
SfioaEhlaHpLJyTsnmrkF/pGVqexg9EO6nGBr5ekMoQ4nZmkJ0pPCMnCP/nCBUeTCK7PjGaWinsS
msrF82fcUwFCNOhARjsOBaW34a0sYt5f6ea+2en28IbyEn/n3SAjEpU4af1bmeUjWszkKKB8A3Rb
xig7VRFaPaq4cC7jhbwL1jTh9jJn98wABudcKU/FxQ1THNgNc6AChxhAwzlY6M10su4ez/31lrMb
3+es0nHmMb2aCDmVcNj0GbgYizbBKZdu3mjzmqL2cqHBmdDpxW68PVpuvSkennSbhuqtufTeB5Iv
3SDqtnpHP76UdPoPELZXnbLibSumHKmDdpesBIpNMc6K0MOQtSbtIX+Umxe1TtXk+1iWf2mwcUHG
1OrRwLhIZEn2NOY7mgvuUfpp/VNxWPe/G6jw4mKT4nMBBkzStd/LABJD9tXAvZPCjrBTR5VkBce2
vSDtvOL0NYnv0/0nB2yoLnWIc/G8mmDzYrzHu5janoThnZjRd/PxKpOzPOdZ6FE4wm4lcy0agJkz
9lkUZo7WX9RsVyFKjhSfAjGo76KQGpKvNYBIUAMZhQKWxghdx5vJHEjAwwf+9pBYK45tN5k8Ct4o
xY0Td9g/GNaF+MEqsiF1leOPkUZ7sD9AtUsu0GBC+YX/dL0EWiLEs6xH1QbIz9A5EluBxtRVDluq
aXkUTfHjIXc8IrZ0kVAcik0uP8Z/t3txSiQNVqXsEI0DyMfDaFKTIK4aSE2OEV3Cvq8LCKvmepom
9ZwRoZCmW/IwqzUkmDUhqexGMybfz+oTWEZtS6qyLbgLhgSO3ne4ztonHrY+Tab/oIhi9Pdi+UDH
otxvS5SqxHIZou5rKbKL4yRvdIKQCusOKtsbhA7X1djng4O4gIF32WFbJlNISRweG0q9uH9tpds7
SaaOyHgXZLXFVYpp3UUp5DFtDB2Q+CsUMz9ioPWaPk31TS6s/fQe0u4JRMPuvpwzVLkP3qR4CLf7
hXzHEVV8do80AAqF4MzzK5lswMV0sKdq38oSmPMI1XnezHmRVy6E3GhQrcSmN0qUlJxgm/gnn6Go
XsHNRIzGkbSZi/M/vwUXdrKalnMDiyWyBDg6FMk4tadz2Wafj1IN9HxOxOVTflYLgj9c46W8tXba
obgYzTb7krLyy2wH6dek+mOHSGP4AmCIaNW332oMISeKoS6Ivh7/UVdQSX03AKQ5vLr+P+mLDy9R
cR3qZprqaSOKYLBtXw/Cvm1mIVvQRZBSF/GVLRLi1alMbo21sxvzZpgfn+gFZ441wu5P3s4d1pHi
yXAwBXTx+54AHMVkbgGyJWcY6vkX7oAo/Vcu2NB3RTasO35VgLp076QJlMW4ktRk3rPetB+CrvHP
2howg54ikuo+olFvC0PzozHlA5u1cDki6EnObUQgR7Se+7U9EV1twS76KBK2h3ZXWdlQvm8mdJUJ
Tt1uWGmEYqEOjqmE0h374dFiTLtbQMOb26zOZO7S0AwdcNLNOV8zsZWbju4xKhhasLkqisR8IKfr
U7uaBAHDDbejr33YEl1poS0K2V5ZsYn5R+6r/GKvtJKhdydgRpgqE/deQH0iFMY+bVGm0XpluklX
k/lSYIvADlZbEJzjQTKtyDvHosnAiTIbELM18xVbAwqIpPUWpq8nc9eLyRR3wWAzw5A8YNQvJMnj
V80mq5oDe/igZ+EIpJkkvbae+GydL0Cqe8sSVLq1MfIfz+XcKhLE2z4ld5t2uVuW8XBqhV+2KeW3
Uh0CxgCCcH8Q9WoR8XAidahWWbXM8vXrKghzhflba+kVvQ6xc5Za0Sf9Sca+1+BRxZdIH7iGbJpX
TYLRADFhlfKh77zZT/v69P4tVkTbW3oQ9krtZb8leXqx8A8oGqVJBY3PXmz7POIOdwejGTZ+LB0E
ArELkTWEmCv6DvraVABaCHgc/4P4+lV1keiqyeHNqkFGub/nwKZG4sVlcWrf/HwCYizCbobuj+j+
PROrl79IaInNHPMJKA6nVI9qWRaDhbT89iG11An+9lIIWhNhzN8DmTs93WccQyw/apr15THDzlzZ
a47Zx9fGxq5rMobWdRhD9svnrvWe755Rbm00loWdk18WyDVL3i8+UJ6i0bXGwKwvmFXd8eG5AxYS
O+jvPi6A0pWC1phAY9EOKj9dRIwbRJ+LU/I4q0j9taS4Br1EmOQlqNl38cX/R4CkXpOwPlyMv/I6
iG3q9UW+iAI/I8j16+HJI4DVxdemDonyzSGaG74mVCPE8aeZJAbzG+/YLt3f3O6cKLdad/r6AiPA
OLqqkqRVdZB5XmFiSeMGOFpOUDW/1KsiBNgOSvil5gXBlIrzkSjxjmz0s0k85iAJ3hReRC0xcMrP
T/+yZO4GCsPZXyz/nLn3zmXJBgugzpPh7z+6dcbAg5vO9+S0c2UQ9Ak1+gjkr4/WoazERQDJfC5W
8heyrvC9WY4D0BFkGDWvAJ5rZE06zesx4Y3cKNbOXvFzfsKuvAmDrUPp8I/zyMZDELoUVigLQ5G/
WZ9SfZj/EZl7Ynd0EynWmj/WbXY325c1O1TxhfcQsiG6fE5A2Id6AfWwlzOQXGmTkRe95TvRv1zd
PWzWtgiGGjG5rBWQTKnOueb6MXm2ny9WqAMnZF9jRpFq3J2+YG/CeHGBpnwtTVDXphLnF5IoIABS
dKV/Ru6YGrWA8fmocdRpgsj8phbbabjo9obkk/AJIYnaQN76ZuWzUNe7r62n2qQq7iKBe3GhBlq8
5MjiWnGWkyResxNbhuj0CotAUu2igr+tp6ZQymFXtj3YMua9hdv7aRhPevFrpmgpKvsXYMN7/VMY
gvDn09s9r3vNNJD5tUpqFRqBGQmNa7J7ovfACtX9yQyC6TMMQafVxWWKmoJ44xPc1TxNl3YGeSr6
/oEixfWYhQe3I+UhlEpAHqOQJdQMTJH+j6cGgGb3koQsawq+57yVvixTLPW2Yu4nw5vB3Vu3pQ1g
EkDufPdm9Kc1wmfvqNryv5N7PTSNSMFwnNCdYhVWXgZlSn75+Qvp6LS0EFWRd9eu8aky7NwFOOWe
jL7acOm2+bz1lC4V9jL/mzEgACZ/tea8t+Piteo0gCgwrhyLo2dbItXAutho6tI4kHCfZ18dnUcj
IDZ4WfRdM7hAqoxArAdny9cZuyymeRaQM7G6da9Z/VAN1QXX6iuwPVWvIjrrdR4arg2Ue3tcgJUJ
x6p46CN+Z+0/S03cX6qVpiQUYLdvjyZxQD20Xqqu4UsW1hjSWiWbMI1YBe5rmKRkd9BY0rA3b/X2
su/KQmoBKkV/iCzIszlQAgJjnBK2QEGP9+53oKCriMHKLpySttFCmt8LqNFF2O65qc8gdX1UT1fN
4PtzN/nN1DmXpEwu73v0s3GJV24OeNtjVjUqdqUcly9340Jyw0WXoZIs3Me+3cUCN3kTNenCINek
/hAqi6XAoyGSUrEeBv5hmTjn5zQAK9S/+TSclG1xRV2rwFrmCJWYVv7tWc/KzxXh533Gj8i3TFEm
66pqvkbORLslCH7VFctB/nNXQFa8aG/lUxad7uJwCez8qm+R8ywU8AaBiLFMjXueVNSxU+bUR9H2
l3jpvXGXjo3DLr2MDQfU6+sJ+BPUgfxHHwWA4tLpOpMiANq5YXUfCFGasuGvx2Ubbre9WvQoyWZC
TMDhDxl1fqr04AlfHlDCH2VEFojMiuLml7jEAePgnE7KxEGktzTbPwHHBA2jX+cONzULmuQQTMAL
TK1I9M728SgGy29KMu/luUNjG/SswLimcBBI2x5LJVd3MtWQSXyYFg3goql/K6zzR76rcD0Fs4an
UehjKUs0s655oDwiDQM2FY3/sd6lJrTppmhAe8aekzRlIAytFqTRVCZa4ZGlQXoQ9Rq/W1lb0fHd
au1oVNPLnKQrZqgrHwhn9fbVJHYmF3qTppk/Ao0LofR1yb8H9YM5oTdP64kUBEtaypzH3rAIPoQw
LdY/EnIyZ+ER8nE9AprKVGohlFvBtnllGtj4tpTBsTbZ8UCNyO333XqjPvQhbxQX0Hnx4JFI8S81
5ckTAd8+PIwgg0cBlrOyihK8XqwyfZvPBEV2d8vE6/iXGxmg0NnK6UtfJQAm5zGN3d6G4UdRiaOK
UoCiOeFyP2V2dgA8NbUqrKNzWLSgHzwmLt+/+Ls0ZR7pgjPHZv75vF+Gf9sotaMONg+5Kiovv/g5
RcFv8gesMBO+KyRVxQs7rIQhBQsvGiUNoYFGMQn3tM8+yxrF620dpWudy3xsO0AAi0Cuy7jWPg4L
f1qySo0GsXJ1l6gGxBu+3TfQ5Hs8oyyGPgvAiM1k668RSkoHTO3y9ZOWNlsHl5W/ssO+v+WZN6a/
Z0py5L4YDdeFO81TKYCdI7OSqQv4m2+lzZeuUKoWE2Qr3AuXI7lnGO5PQljehT2yQ9dBE43Vg4OQ
bqMgTtOcTJADeDvxi1gq1GeBOXbLgKdzy+rK7KnFT+xLT4xJ/w5jaSSaKXskwJzfAqB76DGLeuai
y8+uFJKrPIIBcwFe+CLVoACrU4c1XvdM5DW/+dbyQOfJHSiEQy0nZU2XgQTIlvH+yLWGBXGxT/bg
v/h5nPvs6HNYvv9dkFED3iWUCATahTJsoScsknNbxkepeMRGjWDbqgrRExs7NZnXFBNCsFjsf1uo
EyPq+EGmLsnReOYoBJ8faZWaDFQnWK/7ms1ZMvfyFq+ry03jex9S1LcXOKNoql8XxJutLM3kpoS2
GOZ0yS/BMGgaYbP9W3ubOF4tQtjudVYZ8Gte0po9PCetuYlSkPWYjEgUIovGt2LNxHlxokFPlNzK
UfJC+d1FFCgrJku3PNzk+ISpCYgNqjdEsCAOj8+g/e02kNx9OpuV/qf8OnPw2W8s00Ok2+kVJJ1g
hppRnutJDPbmwWp6OOXB/2rNOq4Cs1ogIVLa19g4KOzC1AHDogptVHZFYQbQkI0SGI8Q+2iso9GI
jRXJeO302mE7e8VIqH1Ngon3exPwtB08f6LjdGvcFfqhp5IITbabDtbnHsUIPn1FRfNCN4a/IVeU
c1LgUa6E/MNNzozhBd3k/1XN9ZBM68cS4dxWdpZ0p/pElO7WtomBdalx8botNTl+Ie49Y/rNum+D
uWInKC4LdpRjd814dmmwb2vIrSGFoCFG0XtcMPkeIc3Aoj9x6nsNXB4vy55maozh31oubYnutTdD
HlUHmz+RcmPFxU34XVqcGsEZ+vi9Nog+0j4Er9UUMi51Zfh3Msc+6zPyBO4+os+BmxkUJoG4Vtn2
+OP/TKa/VZhKevfxdV6JZCd8vJeND2IsdRmxt3akTB+yx/33N9g/0/e2UNf7D1FCkwgPCtNANccl
/ilxEURp1QAxo6iIyuRUKGh1/FjSDb1KZqIiJBFq5avCRrRrv1ebvGQEia9uYu1SSiW7DdvxfTxB
h+nrBbEZrtJDFhOt7qwwyVsUNCWwSfZNxvA51hhsQ6YZtZn1UCLAGRfwki1r9WSbfOyZHoB9NxJJ
liB/M3nAx7el0taWSvbL5oFCGeXVfZBND6e2l+Bwq6F1sVE2eskQ/I3sWSNGZvuA73Fk8wOfFQh4
XmhNUebzxOXly/CnPe1zIbfHqSbPsairBGU32juTz9jYdzhu2tcMnGNZUlHHLBX4+W9a96Ru25An
AFv1MAM38p8kbLHUY3fBa0SXpa3V+SJzo6SbtLYKicZxak26Vx4aZHrRvxfvRDtGn71/Cv+gyAOY
aOQ8BhrIpkhssOx5E1lQgDCxIn0BTtjh+2lEdEpuDnBW2OWjQH94GuUNDlVii8PyTthjmPt3JYLo
KRUQfNjGOy5cbWkRfHADsv/KMwziZ29LEhd8iz/eEmdwGxS741YcuO6eRo+npnLmIAItwLGzwNcQ
7576yyfZMonwd9jejctGJgBngjNFtFEB7TXIwrlt6SpYmp3gH+/PH/F0hg/KseyF1Uyyda8wOQnw
drbj/xrNVyndd+ydslXiUkrIAdQFYae7JrByT7MS/zeGEwY0I/ISeF50Cz9fJnwSUyB8hZ3i1Fm+
GhuBr2bLl5HU8iWxfntfp8gG46p8RRo+sawnvjpGQ64++0STrF1x3PDaeo0YgBI64DdycHG/M0aa
0q2ixj2+RE9ozaS27zxToXIEZHo5VStQcsJVIlmNAYzcnLJdykqHAfdz2FFEMFz+/iEsa4DVUlHy
mE0ZJA5+/9dnFhjF4rq7eX6FwYrq2L37UQ8CJSWWfvI934QARSJP4OeyBB8KOnwrqcrPJKSX+9Vp
L4Kwx62nWwpnpa8D5H++L6pzlQJfLhZG4mZ/sAcin3i6MhkNt13+yxR+zTdjxce6y9ETr7y8KWy/
YrseHe7elg+PWgWxF9AJd2Wl7Bh9fPgOMrxFGrrov7KPnFDlPdmpv10a9Yv4nw/85xQXZNMdrpuS
18wARABz0zX5hrjB4meXFpJA/A/YEZnt+8vxAyJla5oGE/vIPIvIPpnPZzBTxKxV86YqocXzoYPC
QfZTg2dTqH+qXUPYgmMojfb+dfN8mvcM4cAoQGNUM8qW5A3g7AOWM2xjOvDYvaN2t1KxAd2uceVm
W7z+Ya4L78liQZChmQYA8GWcvhQqglEn/QtwV3rY87gRPQ/3g/y6I6ozS1gsyw801BSmo1IfNJfQ
M53luza717KE5uuGr6HJhYymFhEkX+jQ6ozWf8dsDOD0Ulf6fB7VVTAsKEpE4cpt0fPc4q9GZu7S
kgyQo3p9J8f4Te19hX+a7gVG7vsHSsTHD/2PcoLoLgt01ekqLdT0ykYPv6upakSqBOdCFn/Btx25
k0gjszfE+3IscVqXwP7oLJEwgHcars1R9cIFDpUf1Cc0RARuFu4hjKUEoJ6vStSuk7IOijOtd/EU
f3LY53paOfqeIyTS8CriR3/vsCXjOuOm7IEWa0waAAOf9xm1RfIrmyTEWMssvJCPbiWfmo6DQtE+
qPIMk2q+Hy+QrFapMYOUDWBQMQ8mcWaWTn+rWjYtiH+Eorqz5eQdPdyOzlzS8TBdsDoV+5yfPDr8
OR2YLYmAoVzjl2Z9mbVkMhZWE40sJuKbZ3XXnKT13f1jNJE7d5RMiuBvTExVVpek8PJ3/Bii9Dad
+cK8ZVk11YJu1q42+XI/HSfG6X2VfPO5plHk3r8CGE8BUn1kl8cf37jq2ySYD5GDm1uXBx/3x6zT
/7BOjbnGfcGNilzPLOuXe4l00DzeXnkGSaJzRPLhIPS4yFabIRDcsbsjj6QjozN+aAVQy7t4zSsh
8BVIoAStmWZvAnjTFbSkSGUV4kT8eCBaqcy7Xu3rZLauIJTO/bgfglJDvnym3IfJsTV+vohOAQjd
tSP+7A7srqPXT0mP87pnkUZOyL4ArdVIgq7T8/U3moXm9N/RkWUb3ZSzvfY1ksxfrjY9+7aMRhJb
7YcLHXS14pDUvTpMg8qwMe/emtaRajiAOQj2dwrAKBDPVfBHrtHSW76JFbnXRaEXNzXoH+XnpK5U
zMH/YqLxydLvHalE6AlXZpprjLZ8B9MawAHQMF3T5wCawvpMGywOrW7uk/8c2DzfFWSZl9K2EGFC
rB524Wl1HYvB8c9WQ0a5TEy4I88FeZWzdZAQxCs9mru7IdM1Z/vx0xdBM+TT+bZXyHtZHmvpGjqM
BdOYTNEmdwa7aw6Lth9JeEnS2e8kSICja0hOK7giwQ+XJWjPGBvv48sndszhPL7Jqfc7ovDsw+84
xi71SYp/ln/fE4eItLQo7/8CJx9fojArwjLBVayO8D4eCSQK1QFSdMglbm2BUdqd94c1IRvV+MbB
F74qFBH48JY56EgvN6jJIVZthnoExnMI9W45mONgbpwB2kOLAKBlT75dFUUQVCb1CxON56s80ImV
jsh8Fdhe4g+6bSSH48xP5mwHR7Tn2l+ZfPruDw9Qw3dyZZ9gn8Fgfa6tLB4XMwHeCpqmnDUag+o7
yuswIkxuEpfs0RSk4ev65HqNAPkGacbmN/1BzpnKSDTc6cFO3NJYYuadxGSJIAleXGDcNubv0Wjw
n3GFiRUzmfq8HK1bF6zqaDdlCP2mg1oNdCQDBPEcJSnSJvv34s55qlPiDR1McT92zMWgLERA5MRL
4fl8CFAdOF8i4OMRM+vXT52GDkPWErRPJ+Q6wWszhsVdbLCLephB5wUdDrUQKHCVDAIbgEd2bb33
nbi1zRXnGPXkjbY//VBTbtgi8pYVUcIcXW8AlnnxT/fb3WpZKfxQVQOBfXhCHsG4FuKLNL5+zNee
Rvdzkc5IjdH5MZAB3ZrGshlLGOtz+lZWa2PGxHvQFZ5hXx6fhsAAoIgGzmUaTN8ayO7yCwgwH9dD
mavqHj+19Y5KHAxeXDH8uQn2AXiRX8DIRYhGPszDpYMWQ6cMPwa0Sn7P9WAiRHE6au3uxYQi/E6E
bxzBB1gkRa+ip2+otGajH3oKTCHtX4KdYzczhjoZzt2s0AMcwgfWEbqOkYIWCiCr694N7HksISIH
1kY9Ct0RkP33bK8yCFRRKhhVupHGVWrqHmzak5lD1wrCpHbwCf/ZDvNMmWI4ffWnoIFFAIV7IAG1
3wAKNTFszq31lAfcpVson7txKyYunX8unMGSLie9SUDFrU7wyhhjqXiLZ95CnIUYR76pQOF070mA
+VBX5ck6JFAL086K1d8PqHVlFo75g6U9w65cUBcfBn1WGwS5TF6q4MWbDJascNi3hfa6gBaRnLj5
WUv0VpLGi11Pq6knLlT+Pmszqs/iTzA+3eGW2hgDpgpo5Ehm32ACS1SoTrQpVmL/h4anQNlSjglz
3hkD7P6uPMP9p2abWT8p/U6NKbm+L2ikmdcp+zHAOM/7fBi/W+Suj3+KuJ27fh9OWIX31cj7VsyY
yzHW+pZ+lru/gSc0BqYayAijQjAonu93DUZFt6dVbvfxSvhL4odT7tzvTIMt1jw3I8/DZC95dYM5
O/ax3FQGIZEsh0BU464n3u+HGa57uguniPzjPamp+++HsgkoQTesl6oVRIwwzSMi7py17E2xSfe2
zMPs/IXbjJ604laCOkfNoesMJ+8qMnHP3i+bp4LbBS0+WlPSqPFQJp7RsKII2JvzKSViOpJfAm5V
CVzWtnYUcDLdDe/yMi1KXkflOZ92bOMeQA79FYkOzunke0KADVDHTIisxMRsPGyq1IOiQ/+DKOtF
6PSmSB7cTaMCuMxBBS1AqJrJKi+79GyL1DzUs92VnvdR4nU+UqDhKegGNvLElsV89DXHzmFuAmfl
W4qJX5zXBZsnvEyqgqCiqGlUFQBYR8SClLmLOxtdHgtYG0CqWUBp126CdQ0LbRFOZn69PuFclLkD
LUkoQVpGa6hSS1l/zN71TOMj9fJzqJolUR12rEFPF2o1Bo6MP2HK9Wv5vIJs1GBB4IKzyhNxt3Aj
5s9YhGIiYcMc7HFKRM6yuhL1FoINweRQk5ZnSCKn7kA5MOn+Ki/dUuuPxS50XEpuQExx7M3GIGn8
ZP5nHCDag8Bznyr9rMn8T7ZKd2bIw0Fw1m9S6v6GccK/Rjojfyt9uqq3kJdxvitOeHtmRn0z5yEn
qsqb5KB9WHw4edcdXC72UpxdkIys7+/02yC5I2Txy3lzbfs8BofsaHAPmjTro/Ygcrm7gBUXImme
lZCYdtfAu1nnWbkl0QXcbqPxBYBNj5hbbu6lv92bduh5Anh84pcN4LVEE1PVwT4dNWImpNuYqiYs
nfwxmroMRM6F+xXHxQScrKYbAddBKlqv1zya4cbqHQ3YyWL7ElkBxf083ISGJaCQE7t0ixpLZjg6
Z2FGvFirctShrY+T4eFhHTko27KO9WpS80oGy4VvYxYRZlzwUaCdTafkBeVWU4lCvmROTRjoBpJ6
pZm6h5o7ADh+sY0nZqpI435WLHjpdUaG+Inu9rc566OLeowxu34QxfDCd9Ra4tTGy7NPFvx4dNGC
LpHbteHjEY0UOYtrr5aj65tJftrhgMPR0xORPi9RTdz7poYrd3LEWDcHaNA1Zd/Xxrh7pHeE2Zz3
qEOTacNJV4gjbSOUwshUgyaF7qjJcTC7EKOG64Hzetoqzghi40eywIAadTCkV4Ge+vYUuYjPh5Jc
1lnvrmqnF4h69XiEscf3tQ2vNTOTBPZD8Wb69Fk9G07iVXn6gCmUdwPmLRbvu/rRyYfJvzg+QDLb
SrEmbA6zF4+b3+kURj1gzQLHIgnVM8fCcnlf936NEopF5tns+pkXidAF8HjLmmz8AlNsTr2YIQEb
RjKea40H3JOTN+rttqt9qTF+uFRCgngthjQpZmp7P/1dij8iwiIMVC7aZObyrqASdIgklfPrzRBt
N7TecdB3ZoUVwcpDavpnT/iF1Prx8dEnjIwoiHYWn4NnvUeP+IA3g6c1gTIg8xOBaYgLinMvHWBr
BzUb2W6LWO8lOBdUtR8AQyDNnkOmUPuaOTbgUE6atXrRHEtvlv5h1jtmysiDyTJQ7BVj1sdFPHaL
I6wJ9vabzATtUh2Q5HtximAPuRX23LQQ9vlVuMI1NJ1BE3ejwx6gaT8e+o9jgZoR8yXz26KtGLt8
S+YtEDs5+bQe2ElXwmnra6BqW+cSJIfKZM6kBJ+lPfyqYnEX0VZSsZXdSeG7E5+/Sub5iwFjxTHw
fHqR03a7x4++meqCKUcJAO/TmDlmizHfkmsRONaGzJMdo7Tajkh+sqqFnmJPj1MuRsfcCw03oPCS
T4fIvWwiFB8DQZ/VAuX740k23GtZJyXs4MokcwnzyknYZpqskHtjka/fdUkKaABQeJm9DCB6KB42
qPhgmet9U7eXxBiR+1vqZjJUzEHaDRvIOY9vl0xLuMoejZGG9i9F0fCGQ0Xc5zwsZMtVTxJkpyLr
IWJ5HY/R7JI2Gh+lFYeeJCiaOku1yC5fkDfIpmSfMzC8II5cA8yj0Rm2NFx0fPmWlXkIn9/vHAkD
NK54p+FchHRPkdNZ3+akqYVQzwza3lQnPTxDkDG6X79Eg4/biKWkKVKDVvmofVqLqWtICgXf/jUH
PdCD1HF5TTkeo4Rg/56ziARD/m47GNbVnAaeRCl6RgmI+7zqiSDVAAvKt6oM49ffIwLacIswNwiN
laqj4PxpcD4+y+4w8a96gfcCDMOvyZK73TypdGtUfndyh10vOpbcfB4lBoM78Cqy6iEadnX/w1XA
Cst1Y6JDeuHDQNUCZkKeQ6RsrqE1ynqt1fqcT6rk0ykuP/IvJ973fu5LGzNjAMFt3WH6RvuS3VbJ
V4FgC2oopuNMSGKSusyaTstmwo2YLLBNYswwNFB7Rkmh00wcChRbYSFpMeM9L2RGRs7CwEkMxCZE
bbhHvY6gTO2/XHtCb/nye/dwi3qYgUEqFUgDeADbmTrpLO4D56PUM6K7T5cP5W09Lrh6h8UQCIWP
FCy2OqiC02VLV3LWi+b4QqNamzpLGVRQ67LfI8a0kN71PZOtsbFP6823GLZmdxMDCrPk7SBKSPVp
im5PQKy1ZjlofmVzixfabKkqkcQqEqd7rMgSsr9agqiCjahfSGFw2bLwWgaf3JpJVLsMmvQZO0lU
G8PsxRqCskbQjdnUBUItZPUvjK2g1Yt+Vgge0vKkRt9/L1BKCMlR2MbqEkLEc3I4L3J0Fha6csB0
VAjuPZK1v7ZQkJDSWABNkxQsR1/n03pNkpszbpwFBqcvkXQOOuU+nlr6D4u4OHxoRBnLsIjl3JYb
AM11UQGlj10UEJBb22Nk55gjzMs3fzkaKICnNOS020kJFUxDsPT0UKtCTaD+5c4yThzrlQJw5M5i
bP1K+tk6WEhQlZDLrmGCsPi9cPstPKAf56S9FwKQ/BjrzjisC6HOigkHpQDLWZtfU83F9WRCnAkT
+GapTM8I6/u9VfUYVIrwPA22/B2mqs+0MjPEXAGmI7ad36cvdyieyR5OtsfID5XxofcD+R/ELdV4
VJAZzHjntKCUA4XQ5rQJ9QnW7t/syppzfXtW3p50Pq+ZSZaynC0vRNFpxSVpdp0B+s+/vyrv9Zo6
4d2fYP/fohM1VEzmh28A7KIlLfNV9SmYm3khDvBRCo3nbgFgWRKJljTG7GutdV95mxCi0zh2OF7l
2rXkU1ZZlzgkdXQYnxqFSXxQxsWHy2YPh2r1GAB1qnMSf3mddX44m/BeDpa6cktzfmDl+QghMl4x
aKQVRi1oPYh+rUAdubyzmmoOLjQxTv7XbJW6VCtyg2X6uVMX4t75oOe2K5EqE0eA7NqHD+Li+uQp
M0MQ4e6vC11q3x1jsrprlxk4R7e5OJvmZRYK/pillFNE+p/uPS8yXZpfrIBns+U5BDcKGUJDW44u
+5p3fOpTVhJQeaI9IuH3elDwCq1f617IuQsRt5VXo9QSReQxkKodx8tUDhnURJy0s761liBR5rYO
XCCn/bvoeJSWnm9UgtoKDe5hrbGGHYsjLNHgmtURsk0GFn5rEMGNEOzAQyf6cASXvWSTAk10qEiQ
m2BR8Hor+MdBcWsbPxao3ps/jiEXJZ17yNxfucNVy4uMLnK24jGDjmK6t8wYDm2uGTieURQSOADE
r7H63FXkoGk8TFcbs8nuc7G8f0PNybWjAQWlI4CdTeDogfPcWH1k9eCJgBkTJoaoyhevv7eocP1a
xKehRDSRBYxl3Izq5g3hnibs54sFgJYOuVyUT8gdzggpAX3/fk6XpO5eoTKfe6hRcAjnAJOPUbjm
n+RtRZBvELZUK7tQJ8tN9ydmgqQANkBqYdp4rx83ndePZhoQsMwj5JG6gNXRsSSKfCt3Itbytykx
5oNlsfROwemedt+23t9/VJoSy/onx0vNVVRr6Bi1wfxZi/+nxaGSrFs5TFC0yip98Ub0W86q85sl
0Q4EKrBJnZyqrf55xglCr2OatIekEXORz+sI8GeCSFWrE9qJXgKyiRY+NefxB7o6Tr8M6nczc9lr
6iBP7cPm5GBRtHdclTfMt5EFxH0J+AXi5e3XODexaF+GgzShJosbom69puWUFghsbcGcB9woAlXP
Vsk/OS0o9MAmW3ErsI0NFLih/1DLmnoeBcM+f73gFfUve1UT5ezKb75B9lu3yK57fsdYuCkA3KjU
7ykvT13qDwBXUzB9g78+9ESjyhxOqgk6JyZojBAbRl/k54+XA7365Vy93G9EIG8Gm8m5ATucN3w/
ZXycX9zw2k4/Hy2dm2IVWcp0AadRJPuv0HNp/LRPHj82bbZbUo00DJFPeZVqcLI+mfIOonHec5S6
i2Zq9Ynh0HVmR5tMvkPoaWfrABVpiIn9tUZWBzfTdE+BRPcxc2LAE5LoiBVxuTSVjrCJPwuPu5Do
zfebklDCxsQsb0srYViI3iqzaiNpFxeHL5mzkUeUfcTUhEkzMb0g1xnl1i/9l7OcqVc0dOacMXA/
/nVn5XCr5DvI3FaC+IFDklwDXuOque5bLTboiPksWKmuabveH8pym7gdeGeyRXBHn6Vf14qi5+3Z
+p8ibANsOEYxNSreF6duoW/g9gXKJDJ+nx8QnSwXI4HXGDhYDaPNMfPq1OLWfj41UeieZ4SFcNKT
i1eRUToel8Jw7dti5qTAegqUYxqVmvpSCutBXPA8x9HXMnlp+m5LtS3paP71TjGhv/8OiLy00ROt
oiA84DXhXTl3E+2yNOTpyYK7C8BcBOIwipRiFct4brI6WGWnfKaB9j+EseUEC5nbr9bnSg28BEVC
hsK3dwCxRv6zHWTGqB3XHgxf0MP7rJ58h9ObG/Vub9KV2hxiPOcZlGyjzoMo3IMqNGHF72f7UbjJ
BKrEyUi/gbpmFAwGGLZ6Mqgox1nKy+56Wn2vTTCcybK9lmtCuYOKKeYJj/7lWRQikN3cbCee+va0
vMwpEIourXTslf12m/j2S8wbq+FmyhRUHAm43uZ1n2n1Re171+As2dGTYJfKzkLq3F0flnx0Ob7l
BQnpFHj5c1SHKVGCwiJRiOFkWp0/VIfvLmNuN3dbdmCcJ4HU7bdTwYUsmAs8YNHvpQQm8yqB6uE4
zk7HF/s7acbDAvDd+r24E2Bw+hO5gWdAAKv2wYPymKrz0DokySKDIW5Qu4QJBPpLwTKsyc2YcFLh
vV1D29KF6PchHUDVneWag6ttdffvJpyXrgBgFnohZYY2jPfyVxjUeEbo0j0MPUY82jN7UKjR5SAv
PUm2E2UzqCSQMO2dygblQYsQJ6oPupDjUuvSqcigY9FyeTmoFDq6kl/jDSte9/nlR5IDaH36DFU9
3LXVdKl5jxUSAQruWz4iyIU+FxHn+dPTvyk6bqfxgkP5REhncpXMeXvV0+Pc6hlEzxDlFGxMxoQF
xJIn1aRhT6ykC7wr9aSmDE46tUjCBOzA30SQulig7segSk34oypF61N5IwUXRhFdaf61eIHDcGTf
CZVz0/RPiy6YiUEvCl7pmIE+K9Xh8Mg0flPfvwJpoCd7wr06AMTZ64gV7yC+T1G//DHoHHOJGmsn
aAZZs9umEFpesfY4YqvHuyjiW+h6UgTFcL/n6YDycdefoOk+U+xxH9mIqJVr1AnO3CrXmOuGV4/B
lZGnWEtNbzZ5pKCqhTSnRbpwov1wCthjhFnClddAhyRJOVV230ELLUTysHgnqNNIzrB4GCzjljC0
RDEo+DXEtuXgPrgO4yhVmik+CLSiiavHYtdxjmSmiEBKrFegzM6RkdlQCEPk2A8TH7OBJg7oqeW8
IDa6hpOYxOYeaHRKcSxz/lJttNhIEuBgHMS7oQbf0KYBka7dh4Z35t3f9ByrS3FQVFXxCyI/fK7H
MeRutNWNA0SoDHxJ8wQoI0FZpkx+b2iVrFpYxtS3DFwGbauA8HUMtcdOHXGcMx3KqOHWdoH8xV0L
7RNXOfjgkyLSMv3GFuLXHg7NiAmbAlF4TsnhxZcX9txuhPOirgLhbBJNzBJ9hgqH/pGDksTE/A3f
BpJPWLH8LB5qLvil/J5rCqXSGFNGPNAeIssHUJgXKJ9vfEmgGebFuSQ9w1P/LRTPVXFzIFxreo44
apzixUH9Z/3d4rDVW9WMEWsvM2jIsucNyIstbSJ0Kqyl8H0SwNBXC78MRy7wv8JcuWOBKlzT9j9J
FGiTOAaml8IaRsL7Xf0jppuP5csdqSDuMBwy96LgeF66QKPJRYZDR0J/INFwKbx6TMgGFKVUIr8q
prQ1c9nwJYQ5LuC4Om4rW4+0TDY+eJZXwN00W5VaaBD3QBFVJA9ayJL68Cl6cqnTebMMrE/rMJNi
B/qCg/CEECWWUti19xAl7ZyivNDO46FCEKEPLqF23iF6lSwtyJpsfFEDIpWzi0i4zF5mAqLY0zF0
keN9lcLYbhpc/BpxAssBcZHTl6fAZrVWcZ/yCJlDugdBfiJeqXw0ckchI4ZO9XYKIMYLoOHKvEJ5
zAO+RkHWjQd2et0ZCE1cVFpdAKrl5dAugeAQOrmEGkgQq2BY0vXWTso0cpcxiZ+y9atur9vAlucv
zM+BVrQb7xKEAlCbNVKPRKzG76wuq+tujkXhFy2z8REJDjXNfqsX5WVyxBcyQNGz3AGOKIEYVARv
Q3eBOZ0acezr96LEZItHMFItSaJYo+Jgm8WxcO2Y7igJTsktO8KgAxOx/apXB7SYalXSFzoYQwCX
qQIY/YnrbnoFW8xuBlpJ5dOcb+q+HDsqUaF8A6jH/Ok9yA/+3p+km8W6HKjD/SVkSoN3zIzFLRln
TonfIciH/6Y0jqBzbFvNPAZSaar9FDJ7CI6XwhKE0FQd2LM1ncByHUPw0Od7mR/hTcqQ3F+WsGM9
yuIRbHm4RhaZtopmDJeXVHMj/F3fdppzovO0Q4QJwbJ1tT/2Gtw/divZdd8u0wXSVg9JIfOmLa2t
ml0RqphdSrUFjQYeLemZZuZv29SkQaN4WanDHjiVuzK9sLzqUMeZo4mLwqg+lUlCwCmSnaAmqhgt
Rx1pDmnQ+yxJe5pO+MjjbiaTwF+GcGel/dAQh5sFtQYa1mpc5TgUBeuy1Cy3JEsDwKwIxdL2u0tO
k5FS1b9J69Mw9/1E8IfdWWsW9GVVyEWu19st805MX05b1oNYVysBrddMdCG1J8QPoCt3cP2i8A8B
Zhn9fWWiLyL7sgpmV7MxLFEL3tSim2r1iYWspc+A6VyhnZLq7dl6d3hXm0r9ydXUhs5iH3uEM+/B
SVs/IF40hR60wSVgQvcFO66B2j2ArCJ737NwskwQrY6o+kaErs9pPZ26PCJraIufCfQyIpXw7yqU
AaRSG1+wVt8yRR86NYLRMxAGPk6QdMNSLZX6VahC5fDnqlLk45785FVGLSvQLh20UdFYwJ8jNfUI
wjw9PwRyHuW+r4s2RMrMMUbdKcgnoUUSUjmxnjkWhy1uyV2DyGjI+ta0/+qvS3no0JatJYrzWN93
emLE/z1vKNUuofy4oGt/nBNzqDveDdQrTyXT4HY2GMj/UwSenjGBAk1OQsBct7wuET0Pt61TxB7B
S7biZmlomVp/ZxJxn6xFvlUkBik8l22xWN8V9u61zBjxXznUsbjPdW2sXdNZVirfQa+BwlsJ4sbt
5XI2Es06Tu8xDCidMexKd1FMUQPa3D7oBOLNUC4/Ol2UM4f92xAOrTPY4WFVnHNHG2zwmGFX9Ig+
I2JZu2nKbZzn/gBX+KRKpJs02XLMFUPdkjwd1CviuOFT529VIzlgPI9RKuOe60cEBFAqN0q3YRob
ECRCqHmf0NYt1a5fenNcXH9KPXzvkZYzPbn7HfF7xOWBvDfxlFCrfQYO5KWrk4Qnwha1V8X2od9p
l51UeiaxMmzRapEAt1+MiOuyiROk7cWwlSrSxBaHsN/+zSl1+5MhbbkUhTxK2Aw6ubgK2zwlEbr9
LSR5HZ/FzHLpV55S6hriTQ6qWBPSKnIpG8rskBswQ1wYAbfOF8gCsuoEnjNMa/g7yYYnKzQHVMW6
8nApGzh3P0V//yVqk7a2mdok6fIy7R7rxJUkTBhakorbFMQlDnRSOoP728A0Y9eYtyOUNny3VoNl
Rp3m9pp8ImbSrnskS/d/7qGP6uCFhatuj/qh5HiHJQLMuFR8105XVFYwELBg06OwGd/S9NAGwz35
oE5VBLzRpaw2lWp2nbQPMn9KLO0aSuaJ/S25kBCgUWHgiW/zn6gpDP0DsztxN/9Bbre4w5RCIxPv
yfvSNrhCZJ7Rkw/aCjReSDQRBJ1J0QmqPwYy4asyvWLmfM1smN3HBbGkg5DIbcQydIlabEXVE08a
Sy61LxFI/byJ0EBokFYJ2LDUPrC1ot+6tL1gn+p4+iHwmpjex/yx62Q0zp0O4QH8lRsg581nNTKc
B1mhS9qGlhNAhzKGgZjSSqHK9Px8lk1tuhbKkoYEOJULGxuyohAQ22LyViW9e8+divONxnQS1/EW
YIkDIQuCWtnNLMBW13FrvgCmZxgWa2JudQJjMl1QoBJsYBpgS5StUbcujdJSNziwSwPlLgXODVl/
5ogoo/EeBsJE/gKZu+UIhwWg0tXPz2WUsON1r3ectDRjrbS1pNuXIV6lizNioMGRPyBleBjVOeo8
Wa+S2jqKo9oycxy7FovkKLSEoFF5MnAjTpsXv5fRo1ZO4J+dqAs2ZPw3wgrovq2oTsNiwKvVbXCw
xOIiAe3KVYxCHFG5pz0Iy7bWBDAmKctH3sQWBrliotytlxGHbsK29wcroPhYd0A2Y4mpfBYHtPYd
nrYsg6Emv3ZP7Ie+ypVkKbsYpGbZ5fqZWJ8lcR0Px2DRnkh/hft7ITcMZK8URg34+ZJcxoKjn2Rd
qR6i1d192m17el9UxuYcGh/Mz38z9j4uiTZgpa/ytNc9loY74G3HToBOgDkz5Sx+WYoFzFzPOAes
aOdxttul6cpjTBwpIrhKFgwbY0UJ+UQM3EVI+3WqrguRnJdGX275yXcuej8t+kAi30edAT14JV/T
7BkdasumewGseKDxJ48S3aTX77zURlLPdNCjR/x16EDPrd8xALm3svKpKpzkElPVmbaKC4rP5SDw
1n8oX4W6rwNxiyeqmqT4a+EZokkDRqg58L0uJSnkCdzSeHlvCr76lzUsW41OmpLBDUC4hr7TO4JA
s0iNWGVCXWdqKMABk/fDyX6na3kTXl7NokrQKa1ZXbNeRwFJHcReGvuH2PoilvUysE/+d59eXD30
aWkUR0hNW976WN81zXYF1mCENINOU+jLEbu/7ToAmxqq1BpLgYvhD5eOCuPym9ljpF4ueKa7FlFL
RlrJNUq9QSwYEsCsKZf5DsivZBbSKYfVMCmAXxFlwoqy+W0JcwIW6M0+vq2JoZz5FBq7KpVZxPXo
CTVJYNxjBONgtuoOJmz8yr+GJMLnbe/5SpknIbHOaBWcmUg46SFXOTmdN/c+X7TD9X0P25F893lu
2ChMkxMuYxxyMrEQWp4iIlvWMXywCWPCyOGBCWWvzd+Z9vJ01TjSua05AAUqcHKa2xnk3tCqtG6r
RCdll/6BqTKoBl2YLGez3mZUvaDx0mhoeFxaHcd17gcss3+m+fty0n5C6+FFB6fHZAGYLKxIV7DN
YGY5zcs5Ix7b/xBT81fFnun3lt+GkK2qiE/34bzGONUHThWoenEIEFm4SP1Y2bYBeiKwK1ULjnVb
5mjq8euxHsklpwfCVbj4MiEtBcGUdigleyss5rQwG4wuzq5Ni/tB+fq92biZZESj+I9uUwBus7n9
TQ7cUln7lm5CKJ2PY6yxRVoxvt9NsSeyhsQnz5fnIW4G8syqU7o5TpQ8xvUg2BfO+Evpk33L8r8R
XnOdkek7EaeQbMDSu3JXNh9L5AHaOhOdfYeOWVX+lNo4ZA1hV6TMiR337IQxcrhtHWimg8WBrfwN
D7k+MlpPb7txcgJriMbP663kmAOf7VO3MO/xBmPe5aich4LxfAsKAPBabPf7edoBqUvtTlAsPcuj
nu9+Ri5+K3HI9vFKJOjY/GJ+U1yarbEXvr8uw9sQVc1B5iCQLeb1888cvXHxEOGoJmr8CiIIlz9b
O+KnOSYDnu2PR5Ry9wC++yRzRqOvsPihxfgLcfirKMeX2y7Tv23mUX2GqA+dlpyYFgaw0ICYuCiF
NFALsQbKQFfI33zNjbxYXnW+FYG1d+BSpnFT1K+vCoNlTZ4t4j0r6gadi5nHzvj6gYSCKGOBZqBt
v1Gw/Oqu6FZQxEl3fksDEN4jLlm32guZws+49cueX05iVxUhsxfGvNEzhrWU53gLUvYH0GMUyj7F
xrKv8c2NM8nB7BblAaXG7f8uUy9sqHgb9G0lHbgiWaN3xUYRn5ZzIhkmdLV3ANp5Lr1vk+CaFbyZ
6KwkbXdgg5mlaZXm1iJEGyzE8whawf32y/yt66rr9dZbLpVCxbjJlEfIcAN0kjXPE9751CvJVoD3
BgucLsEOrBD1pKyJq0CNtn5A36jKc322a7WgglxICplJF8gv55DdLA5smyInOdBgfJDZFnuNrNSJ
xGNg1mNUrrRV9hz3oa2hRL/AhFlrZsMnrWKM6JrGV0ZlkiJxwauK4+z+akdvzMadfAlmBiO3b/sT
8DMXgBKw5kueeTDXRbAt12JjhM6Dz44TsAqeet+4n7l2siil5r8MtpUwKO+h4OwDfcjb0wIQutrU
It/qX0F3Iyl7WNhMGRvYNPBgJR3aKShzuN+dLp1Uu5EEb5IaBDn+6QRluGwEDXiU5q6TYK6oDFAI
QU8dkcb9eoeiN5ARRxaZ2ECi26+whBwYACebhdAXPQFvjZg6fq/MTc7ia0GnGMxTdsPwGeDdHOf5
dX4wyNEP4wXDlciDkYKP1eltir778lnHf2PJfaT2V3wBqU6PdZqXtJxBXrFN3Jsj84SW1zO57TF/
aZggLtGRUX7Y7tkL9sM/aE4srBLsxbwjvXto1nnYPH2w1G7qz7Ly/daUhUoerYjt2PS2SAFkrQJM
kKP3dXA07E7h5NJgDaGfRWioe7SLnPFipOeteTPkEEPgDMEtkxW+69XsQ28tTPSYM3yqznuzJOMy
gXLGKdBO+XXIY1qTeo/NIxQv3A1nlSKuOGTqQRubYgHZnBJG54n5ERJCGIk/tj9ShFt/aALPDJmR
A1adZegT0qAIWzZ1siPeEjv2DL/1+gfhgxGc2vN1IYERoZiXcvVSuOzOyViz2WzcMGEGLLAWCA6K
izKgGboq0iREX5Mcv8bb1nAjpX3vS7xaB9BIToG3Ogn7yUNXy7zLL8gRepcK6UdlQig7dHMahpcI
/EN0tI+T7EWL12TVsmyxMSVA38ek/mtpeJTI0GLsV89ZjMMn0XXSGGvy7Jq6o51oqknBfBN5V5Ab
R1M+bP4flxrmk2Y3lKxTg+BoMaeSOIlOCSvIqhH+qUttx+GFMjE2FIrCz6/vuFtfW71SelYnu8iW
VHryL63KE6S0M2yEEkE+ARDoKW0GH875g0r9EZagXSE4BXmrcsdCOu2YZjL2fVz1mzWZEqypqEk3
nfmkaYgGwCBSJUbG3tt9W/0ts17H6IWI9ter7v4dFlDjhsU3zWm0XIZJ6EuB/e6wa//OqGnzeFVe
qZ6vZGWjETYkzcB6h2kcuBxMn18tYY+PJOQ5RVtJbvRvPl3IoEWl5e3+BcpX8GzDoR5dNmd6DeQc
99MMxcHvunXNZbt1qJamKUf0q1OkMthSIsRcXpoJGUOHy7lz+AOYrnybE2hKeB4GhBJX7hXya6zZ
VraUXdbfg0u3IXN/Moy4sh4FNgDRoajnDHnon/qDQ3m5VBClfpKqzOPq/tzJeET2V/xo01ST9H55
DSDJjVaARQ/QXtZXl/qJZMEKr4FS00V0KTAJ0VNgcy2jPENXvKwNTJ1k+VdVd/3XWBdIn9mTPYDw
lAq7PBJGDfWTQhtxDIrkA+/+H89Dr/aquDxIcW1ZVaVys0OA9TnLcyL0oMfblf6Zkh7W6S11jwiR
Jdc8mS1gFYdHqlp/So+U7b4jxDjZxj5VllJ049kfrLsLwT9qA/KnXAYR55qm+faP+RX2HaBQgHDE
SdQhypdI/KwmK9D0VkhxOs3d6N8bRlTWov6f37p8DbIhtEHbwAqng3qjd8sN2Z/SHT4CVSxmqoyG
vUJtzmzUSh0AlJTp+4pKVQfcm8IXongBqPO3zExRADrz++DF1Z8g5CHY1TBd+UpcfD3LqLhJrFIs
ZFBiyiDWS7xdO8ctFRZ75dVcu/l5Vx+zl5ZfUc7yaFbq+5gQPNmMOCiE0yIyvOkDciUHmmfuIg65
z+Bh8wDyYKxjw3h31IHcwghqIRVK4//Ax6KQbDwAQiwg+geWfog0g9hhCnaP8fQQrhaKE0Ex4RfZ
HqWRipsDf2pmmgIPZNQLFTTcMmzYqVSjwP7xjsF2yWy5PA0eUGXXe1O8oHylKn9si3w2y1ANsd6r
hqKn6u8P/YYlt2FDrVSrddIGj547L03QwIG14E79UcqW+FuyFYo5swdRzLmwllAsJogzngL8+uJ8
3az0j47gqmM+hdTYw3C6nmLSR1UpyzVHlDxdSjHB7unXm9j+HvRLzG/UjdlzubVV9tc7B2AITRmH
aMRtDt9yr/WqmuXiiDPpGXOCCkKu4zIGYmX+DLx4jI/lJ1Y2zXOL5TU4RoH0tWj4HIp+ibkb9D7/
bwOwzBcZaHSPUn5y3ZFyzA+JMi7Y2OpV27PClgvrslsDRZXOjzHz6g9vW2RaRpWLcfNVhy0sN0xw
zobLfQkskXREMJVE2U9+EJrQqBG83GRn0ZCM3vVIEMGwzmEZNg492Drp4ZQkM3Kj2UO2+lfo9b4v
M4z0c7Mc09OUENHi/OjQOYWKEie440lsjNqRHsMwsiWhrhMan1ixdtKJ0AsOB1yYdWdgQaiOOLXF
lVL5QfT9WKeT1hwt/bzl4KYXNw3TP+zDMtk6Lz0VYK5oCO3nabWPFwbQcpMXD3RVV/mgPNZ8CHSV
6C0ti6w4KT3JGMigk4DMQ/TUXFupr2MJKSOloHcNDoSbhWsLSgrU688egen8UpLUCjyynyLkiJ9h
tjGwVnjk+e9XyhEa5qPaxzXEYRBpnuvHXdxFBDtJg2LMkmQBNpEoOhH2GeK1oB8NOnso+IwXOXOl
IA47TvluVR/c1t9A1YQS6wMYtw5S45E6JX7oC4GJq/SFNgkuCkg3+OgQB5K/SHV4hVejG8h4kMfQ
h5gIjRW/t7bC5ou5I9rtj8yd6pvECK3kbUYq8XowiWgvk4toQJ2LcBUpHrlrqNzcFCgijbu8Qt4o
lg0LiBK8gM9iepwS0L9zg12gFXYTZL1Vgxth8kRemgxOWdBcplqcjFHId4DEPh1xP/B9nyBxJqR2
pHkTqmqYUbcMY8OvwFJ1+sB5JXj47Us18wRIZcl/xKkJpFgbRHFWa1xW0JcDAhsd6TdTwARkaeU2
cIWACWDHaigF/7rOWtYgcJ+OKjC3qM9qFNjqCuOiLKA2ylm6P730hlSGJBZBBBtMn08t0xjhkYke
8o7y9p/wf6NHZjdZrFaHbiXW72bB2m1ej+VW0yRsWAf2EIVQLYaZpac2V4RvNraZ8pJckZbWG8ji
faoAU9bd72j8g2YD31QDlyrl3EMkM/T1QiJB3UmKwPqU9LMzAqsPzk2UwTctFUfwmdMztJY872OI
vkFNSqmF+Zthv3Oljd9e9WhuikYSyn/Uy9BfAa58iOLHLiDv9wy6d+dboZFho0RXzhvU21sXot23
xuIhsm6WZoEoRz4QzxiuPdIk0tGG1TJNPh/1WtrJdB9hbuL38U0nSeKjZZqQYnd3NPthZPjhHbv1
V67iZUEexj0RiQBqunkNNlwmeWzO5peCScplyd/5tnpPPdNLi2isMdTV5kyjWf4+EvDm1MVI+hEJ
c+odvOxMyUl62vy7/jpWQyd0IpCz6W51RWXk3/jQjWxKhGW9DARxmuk/D9dKTnnEj7spVpMPkDcg
FEE9TG0xVnoHrachh9mJnGljjLGZO8zQ02fMNZYqUf6ys+G9CS267wRZsnzxgP9pPyvcZJlJiId5
gs+agi/FXKhcLDKYj1agYy/MYgddzP3eyrFEI9N1Rwbj6JOcyT6E4PUlu3R6wkuT1xesrBkRlwTW
KASnnZrcKhRT1lUvumEYHjpYbI6hGoytM1nxYqk2grfsP1TTYhdWnnHywQn2G3+os3EZcSodBGAd
SzTcmOVX7MsTTIm1cqWN+ul4lN02c2o+efxosU4IXeaT7WVszQq9CVHeZ73iTD4g8VJQ0wj8bf13
OgQR5ouTFZIhu8TURnhyVJp/Kdk4gcdKOpghdeqev8cXPlRwmyKQO6wno6/D3qXU89HkKq3Dhduh
L3i4lxqTDQ1nH2xUa/qChOtp2byCieyPXDkecw4QGT0F8YzanZ3sbX3X4g79EQE4oE5pAiieBcRb
tACSwPbG3aywGcC8CO7Ga43v67ZiObcrYAMlJKalnYMjxABNbItIaGqZ5StbhoyT/87qIvvciYp2
jhLrQMc+EL5cJ/rFoxh2FtKGqiFV6XjyCpUkJo4KFUIye8vqGjfgVKn6pgzmy4Gym4IzqAFmyPLw
90G2eFL8Yi1xyZFSsKnePniUMbcvoAI45/SGp6pcXq2ucBSSO4ywMylea5JN0jcECXpJdDvp8n/L
YlVniVoeWcsZeINDBH7kgToRa2bMO835psEzmD+Cfi9/g7MOoMa5C9hJuiEhD81H1//qqUBqru6T
t9qDpet5WRfjNRF1TSzd6/qLq1hWSDpxqC1adeyWL6PDwr7dikfZUzCaju4zl3GfYyFXm9TTPqRg
gGsIIwy0zEoctjYT9uPAacRJ1W6FOw2IkUmLguMkZe2RBmbYikEIRDx/zSIMWFiLH6wEcI3uVvpd
AG8y0UcAANGJWf9OUctarZH2Jx8u2VAHKkPXxNHxMgXwENDzNOJG9ifMa4irYD05ibBBM8abJwMj
mTnvSvRgENaxS23rNQnrIzM2Z9Im/E6pSR5yQ4SV6xHDSjlLHeuTUwLqQj3sred6//BBbluNajJl
uWrPLIRhYM5lIOO/9PI5wFJVYUb1R3awzGoKo5uwvQAVcqd86WBWC0rJnGMsQ08BvjEmFwOXfQ1o
sMv6Nj2tzzxtc+qtrN08aGFleQsFkPXenn9nGe2Br+DTSFZS6UPr422TC0iylMFiZgMuLyoMa3Ri
pKfyUV2O7g+ugFQ8q3DbXBhzkSaHCZBe0pLA4ZInbNIyWJru4ydufqEBzV/XeuMGf8vYuA6mxBbu
zOEMOYQEAaB9MJgVZklbsKq9ixIA+RX7BhMRI3Efp/jnkXs0fQ+/ClIRZjj/KcSFxo/05Aclj2d9
P2/+S9BfcaVxUr5VfRyXDYYGItmoICsTyZyGFrlALirLyc6FFZuWCEgH5Ax0T2USizlLBCR4vOyx
oqcIFsJFrxWFq8YvJSzteDxTIdyVXK6v4VFpqsThDdaYZaMG5Ki4AE/D9Vv5rMWz7pcqrkkRj+SM
XL/gQ5g4NWWk93lrNRjmG5h3uDeBm/wXGAo0Y0L9BbTXBpp8HDyDYYPRvd0YzWPKvnB+ZZmwKQT0
4XDc+flLtueS2+/tFbOCCNhMtd8RsxekziV+TvWnEVnrIkoIB/vGaUnURvBEamehdRY3xDHP0v3g
EB/fo2Jj+u81wcLVfeZEPVKmMPMsfWw3xWK46ZTLXRPrKjdrachx11eYl4WaFg+LtnR7wpJvM+Mb
LQBFcrsfOLmFvzU6+jMoscObnyHx9LXt1I41wnn+7zjhoo78lxNw6Tfdbmd8gFf6SVyUpUvlEDmH
x0rjVogyqoht2/cW1m7OK4e2DRx43ocZDXes7QUgE08w4YNjX9zr/delbX1qHldlGSJO0NQdF8Xn
GdAdnDfCXWRvu4Ctgc2TXOt2M1Jv4Eo+BfPR2eiRch4rV/wGEUyNXepYfv8HgcnTwUJnoG5pdywT
gUbJhaCb8GdciGtif7Y2g/GMQ5c0Y2IDcl2gDvp57Ya5fzXKc3Nb6Z4s2BVGH6j31B1qAs8cFuvt
JbxaAB1W8HlDES0WfRPqXgjb3zRP+EbEDpE+NJZRacv+7FHRoSYE/8hFSFdcItDBMCoxvWFd+ZUf
mNEDAQt9hDlCtPysRrO9HW4nVn/B8awVsBm91Fm0KjeJTgRBViiDofT36JrnLd8BNILUNK6CDJM0
O6cxfbQq4ImxLvOGEivkToJ1Ewloybw/SUvKCFCR+oJ2DaTJCkQk7LfpQ45+ZewzxUh96FTNsanu
Xc085Qded+zZGCCtwMKg3mcYWFYwH+lzDF4ahPDm2VwKPO+IkrwNouCc2gTgugFac03itdJlpRhj
+kFAzYmQnU1j2nppONylFNBEF2czIGdr/KTywiLHhpRSJII2VhEIZCdrigCpsQQAVSR05O5eV4Bl
pFyuY6f/UHC2ce89faedkIoIxXlEI567KUARYMU1sUo4Io96Uxh5F0J793gkx6TyxOqPaeO6bo8/
zvyuoBlmVqdcPVTI48uBsW41Q6BpQV84Ef6ZE8Lfu2zUXYzvrVJRrqt6ybEWx26nTmiJ6moPo5z1
lHf9T0/V7Jbz+VBAw+qQRTByJ13IIRHVuCEFS/gCDnyO3QGUf+1eTi1CxbXQfkhuKA+FBqJOq3jy
HHJ7OmKGkZnLNwiO3VR9vejJhSESyjvE2GB6gYXlBuiKEnKH+zr7LryOg7H0YqDGWLQ9pPmYK0l3
fExw9aGPpsNPLnCE3dJnM6WIQUi14y4L45Ao1OjkfhdSegSu9A3m1KnNQEQ9ESj6e6j0s/7EtYUi
2HU5K/Fdxa9H1BhCw+52diU8zuI2wbbrm6YuFJPIGY5XAJwbScfobJ9svfwsJCYJlGGV2ckvsZX2
Q01woD0IGz5q8dV4cIAO6RkXhb5dPkCvayDZ2fJyYWk/KFtbYkuWLUlQAYj3BqFoOB3t7wkNE6KX
kwUGGQxmkWzsv+oYNevGC+Hm/evtqwd2s4EOobncfPhFj9BlxNDCi1nUfA2BeqmTJROoJ3h2mHLS
0TkPLSNq3XbWuCEBjdB7iHYhp3pi38j4dCZnZhmt8QOPTnXJSswqyQCPCAj7CbutaPuUiG2fxygH
WPcPtowPl25x94nkOnqQnFZsRQPvUCVm5pH2kcwGme0VcH8K49TFc6zYhvvk8JozlLIxG6VvVnPO
/u4ea1BB1LqB35sCGel0SqRGq6t4DpV+aYAwPebi4sToXa/AUfcwBOWtZ6BUQ0+TCsdjr2/3E2f+
96Yx4pysoBmQ1TDgOsd3Eplyxq5X1E+6F1HwZY9+15U0Vlumi1CXyA1VWnYELAzOI4Q7b49kyGEz
XrgeaZdtWUJtFX4ZEdkzAHT5NcHZQsD/5W80vLVc4LLBATnuPzDYIm/FGCG3bbwEUY2ip/xMgtjR
mvhDkBcSgBX2syEoj3imKsiilPHquK3U09+Rh3Cv/hiJ4O7pI7bFD16EdakF7xn344f9iq5Cj3+U
80y6S7y5NHH8t1q2Qj/fNNc+tm0ZammSHGjhAoMGTk3hFgvuve2JkikxH1xxSfDr9UmPbM5nLICj
JddznA/VWcy8SmOCOOwSpp2BgdJ0RYOSdcXNYEjwo1JHW77ZaOg9xVcXEGiVgRwYB7xcgIBwdNFa
mCALo36g3Edt70J+qVsNWcETzhPBtgGVRhWWeW8V6rxYtmsIxCipiWquEayxKhXmasq1UhcS8pdm
hLUmg/PQRZT6BIlhJqjGvyJmKecB2LCVZXat9FQd9fdyI4NN9b2hGEu6QTcDFesB6wUHbzWORAJd
4bzSf2ei8cg6Gq2r0f9VY79nX5wPU5UyRSb1HyTNciVkL7iH+ra54Wi5R+16m0D9mgQNWeZufU8X
zUiMkzvYodWu5g2CtaXU+kRQ/nxi2YM53Bjq/Hmccr+n2hsiZmu+Hap753AgKhgElU/Ta6sr63cy
MhOWmsWcicP9lSjt4wvmOTH62GPKGthJPG+H713GCzjrfWaNzcbue7csfcr9+Ae3FlyQ0rlTTXfQ
WMv57H6O4LVRSIh67CrY/Mfue5kvii/rv2UtBK3lxxtqlau527mwRP3vJUEjgHqbG1ISgNCcnLDp
jqWYhUP163xDb69Q4NDyg83MeidJ5zYAsRwkC2cl3M8ulXViFTMYsRXvaFx0CyEvFVQ8bJofBNtT
03dvgLh/ISGR8IXVg3gsD2LALmBFikRHshUBpP8yuDllqSxJeXg82MqVQHlYcZdkqyoa/3JFTgcU
91Sb+9DUerMK5x+fkcrSUJpUX1S9RLDdgzAAW/eKH/2RTs/7z0FnUUDqQ2Be4ti+HBcmivned3FP
37F6FGDmiz7x3fEUB2FRjGaStu80r18fQt7zrxMpsp59RcimP6SKYJl7QsUIKy5vWmCiOInf9U7G
VY5HLOS026ITVf7k7Y9o+nYb1fSndt3Uw6SREPIlrk0LuZIPOUd8mtsg76gxh7xI6HmfXIHojtQG
LLtsx8C8oyGg5K6nxkf0sAnzhsCAo9/TLHhrLuk9DR5w2xfdNS2x/quaZG1MKg7Xq6BFM2l40xh/
v5H6ZJcooKHbGCeC5uCeF+zlhssNWluBaHvr6ycirX9dqfhV16UfFVxifPRYbcMbyRGn9QWGr9Or
7w1Bc/kU/2cM7m1FE7h2wD8oUdg2Jup2QGnIYQxin6WaAGb4kUHtwVx3GSGx3WXbCYNuACk6ic1L
XcAAUIIKq89i99yhn8+6OMHL1HHkOpppXrVmYqt+LQQONQFzsvwm+xGCHUBktnTzGj7D9qpUFKIs
zJfYa9O4R0YqpeGmfXNZB3xnoY5UTFb+GCTRe9Y6REaFCNqwP7b3+QmVYeZlf4ghYdSQI4LT/kqf
VhmzXugjtEfBVFT0T3UGtsjM3XSO5KRUuwicKdAmX+sITIF2YEgJ7K4qCn6PGJt/6fuy1FEsiDPV
8Wfop24gN/BsL2YApNpjW9+9shQIIWHHcjIujB2ATvkMafmWOA6wN1OqU19UUgu/96HuHcTyUAPN
3XyZL94dBNsKbszOobzZXYUa1YuEhrtyMLOJKDveZuKzRi0AI/QPJQYcVAksMp+xxFXUf7wUW6HN
QFurjnxuNWMb3RyxO5tXpr5KKMNwUk1TqqXWeXWH04m6JVMRdR7ouqwnocMIf8TOwtiEKtHJIlSP
v0XFUZuhhT4/z0/gsK/5C5cgMgjKLZv6pTw7vLdod0LUHfyYPFxJiV3x8eanhD4esS1i8B2D9euA
7zflDmmPThlqIqKvcNi550aceJshXKh4VdcvcSnQI2KGsr4N868g58RYa64afxxFyvbZOxMsJpkN
yC9H+W39xr7Y84WxwCvs6hho0a8DTXkU1AHRfLq/RgiSZL63vmQtUAIZmyiyDFqNnbM0DxqXONBG
6j7i9D/HeeQDA39UmgLpsymn5qoYWlc0M5bkt0yu79QGifIDK7FcONDpTuTNW3ZG2bartQBn7pEY
Z6/fDfFtEmGJnIJrCrVg95dQ8IlfwnSAJDJvP8ii7t7P7vAuCm8n6+71qcuXXYnOD8ayPDYLBGfO
Kt0KD3vqvz9TU3N+aHvFDV/kpdEy8JtaDKO16hAB9VB1R1Yji3v4zRUTK2TYvhf9zYAONRMYbtPx
9GRPv9b60f1FKCAikGFmiIq6pL6yOaH0pf9fyZi8LrGEIipyfFwow1oIFnxdRhUh8nTvz3+PfDcr
gQSwrho5Rcevu41NFPKO+ZCEbaQ5oWIQP6Ndi7vCgpEtI71Uy7S9Ze9FRPrp8UsrlOIgh8nml7Hg
nzSozeQ9PzxeOWExvZ77VdUt1e4QQ4+8s5ScSSFwLad43kfvsgWavnZGQV7AuHQKM/pyUkulx8pn
Ed2miZAZa3IgyrFX+8HrpNtabU1p3qQfzPZwB1aiimIUfZhJo+0ZHd5lMOQ3j3uqfx1u1hwD2MCk
fMQ2CwGXL8Ch2BrBvCZNKhkSz38QN4JMH29uvVTVkGVcx3PFGTAECGOfJyK9709StRQCbJZnnr9/
Iqzvo2BE3YjkZIApCqtcNu2kcI/LnyR+jTT2NzFL2BagQeA5Xc9iomUsQjRSwbQ1Hk+fcjRKLgAT
vqXld8Y5T8CL36/iulUw79cIN+rH2KvoFvNzW4X4UKhPa5n3ddFuxMxewg0n4ykkwps5JH2QrdMZ
8MrhIPYGeEWLZaC+S9HYK36ttp8gqp2mDI4QhP93DPUeEYgQ4lQO8/ileZ/v8Vdm68J/tlAynxDT
E3nFMtJ2ljYFGMgbKbc8iQnp3hxDduS8vd1IDsEJqg2osotzo5tF8/tAGqP0lA3wkfzFGqYSykjF
ks4m6KcTlKxIG3ISsBhqKiJ4FvkFENGyph/eZgYM2tM1OKb9zzH/eTp+j1bNpUZRUiB5as8c8lpK
PqWXg6l9mJGvObOuOcr/QTYou5Y+m1bgDqZcCtAHECwigebHKxdDjehb91BN6/D9vKJrHanL/4Tp
k2x6xyMLAv0v7fiwrNLbhT4E/Xi4PCxKYh5qlEfSFXetcoO2qnvSvQg4VMTbs/GpKK6nIZ1jFVPf
CXTmk9cqtpTm+EbLOyhJLeBGcQwmSZ+JS9JR6HtZ/G4rUKHuZlAq8NFwaA3mI3w1A4Y+dI3PxHk+
knH5SkaQjlb/FiWPVZWfl7mXkSsO4wF7yOd8OLsVTxcIhRbTMXWuBqZLlsWRBkCRklY4PfcxHGYy
IUHvsRETGGHGBNiO/r1pf8PdgWeeA8NNYupKMqaob++WC3ca3Sg04gP99LItuByUx8R2gUvBARvQ
dR2ypGI8b/+UMUbt36I1LHnJabtwvpvndGwzDU8UuCIe8QX0c1xj47lB/Zs9rDgutAgIxfes5+t4
qriXseCGHJSw95gG+Ju4bGZuB/nd9svW7AaAs1ZCUr35kvcyCD8EX/xGGXomwZEVqV5WKjxvptg4
bUYBi2pGFwzze/21nH1A2K0Z4kgsw7nsngyVNDjDLWuaJVNp0b7CY15JoYfrpOEwxomlEOzaIX8j
xoVfFaSG2W2oYRYt4VASV+Um1CHpc9QbNL9YKf2S0Gy4/fdRUrFNoTPZsONuiy4o5jEzJWMwcmGs
lrGWMaIMC0P9F8xtaUeSUnKpGHdnaHD/DdijzV2KC8yhk8bCE4y88exdYZU7UmGm9l3xp3vlAR1G
jERukZYEjhe2P04dzqO8Bpzqu8ItNMBAeqI0M4XdKZFIqF0k+W4ImIxag061tLunMxNqmse4ebrN
aYvY7uW8iu/ytxdsbWEFl7cySpJpCsnXARaRP4mN4gU3dpuORHe4yOq0I0V9QGaYhJwKXSFpPXff
EUJe5JBmVQVx33yyGbt1WRjdipEbWDPqKoHVemCv9Orph/rEUvEi+I1+PqhhS0+4o2PBFlwbIvL9
WyKYYzHhMJj767CxcECeZDRGFce1Q8rusWxNmCuh/QgLJc/LrdcwJeznrdi7Ny4g3za1vnbhd2R5
lo9kbhrOFt42W5nRtBlx4iAMkTdq5T42V6krpDmXD94P12XQnPrTUYAiXKIYCShYtC8YtBAcO9Yl
v3/9eLxpIOFkUmm2ofm1kSlrGcWkuxlv7J6DlA48LTfDi6iik5sMDlWgE+KZ2yBElv843RU8aVuC
wFJu5Vl/EKR3ykEXB8Ta9/fb8QwtDsx64t7WSJAHshOoEovKdM2Bic+kjiNhlWO+2lYO2Av0m7I3
2UfHS4u1Pse1964chY5nJ32QHvkN8cMSN2bkufSD5wG0yyuewdJBySEzXE4baJJ8IZVdBKpaqIYc
lednl8XzvtGjENqCwz+6BmuaRPSHobDl3sUqX1VrWctWToxryRDDt4RK5QL8KCvzyn8TMiVw6G8A
xEPgI97AyI5YM8p12IWujxiAxRX7yxosr6mg+edxaa8h7ZkC3G6UZcjwhKyF4VSFqnTUIqMQ8cVx
Ty5a1p0KKCHHZsrhzTK1JF2csn9yxvTzC9QKYzc95s+051y+qsUG2+1eaCKgk2EbigZ5Sa+CCHjh
K7VFOHJ2rVRVynxYStJO6FZJqN1L65vYQJlcHCc6oVjhVl/hUVGywROMS+ZlCDEIv5rVjyRUehMp
omasTaV9hzC9g5HLwFR0xaAzCr8q7gOUpofdVZ+7+gNdVAhmHH/it6RNOfDW0X0Vxby5sIZb42yl
g2b2A9yIx9VFBlCqiTrgqVllnF4mvsj62TEEo7fUPpWeouOn/sftGQo+eeJ/AOnVkL9RwLpy6RPM
9SW9DGbefff6FcK9ix+y9mHhmXKrmYDieBxAuTC6GJ4iskoRlutiWn5nyiX82B+VMHvsUUS536MO
48z5lL5NOyKIBpnFQU0FN+Zo3FUOi7iblswLekUEQAd6qujgIg+Q4W1yiJt3kXLGZIIS+qXcXegp
I4GP/R62G3M/vdDx98vac9/pMTybtzxMHYgB7bpyRwek/gsOUjmwuw1jejnx/P+Bscpl6rCBUHJo
RmmdBg6L2BjzcEWEHnH9jaMf9N4bIWgR42tkNSKEahBc53bMlRpGhkZtUEwyqiq05USnw1qp6B/C
gDBvO4XmOJ/Siy+eNOaFr+IkGpN2qb/vhqLex7AqjvwDv9FTmDlsmZByHGYtzITM+ZDx5QHCuvH5
FYHZCjZ/z1Bku/FgKalo+nzIS7ZXjRk6Ijzy1PsUwXcBBih1nM61mZi94kshAQngamq6yzRYu3A0
8Ldn0eEoL8HvfgjL9hOsRwKddewdUBT0iR+sPE4VO5YwSXBsxAQwfuQ0EnhAahT/K9giGkMdamt1
w4Ihxf9rktjl6HR5+nKiXYNo7qy+lU52rXoKGap5LLiTlcdBX3gH+DcSJHwOtV/UVhwXLJUYd3Ar
R/AdGVMKFF/fQh0ytjJ5iciYI31YRgvKPelRGeylb9JW1F4lsaaGmP8SBOkGHb6VGJXeJ8aJxVYv
Hq7OApH70hO6+oDZrH7eQSS36TVPXe3kpUnowTPjPMpNYP/qJ9ZPrDA+QF+nip3qh9i3+rBQ8nGQ
JfDMRdz9hHlS0YT7yxzMnABcjpQRR9QhoVBS/nq+KuyLsyf4yehH9xJ0bn+0CZukHe6mOPi9+A98
Z3Pj3HOAARS72AxWlYGxWpVzkVWusYrRHzm8br0SJMmA6bt67+gBrTcX4XmuGr0YDGf40XO6+erZ
bJgH2wUyxvbLhHU2Kw8OM+AeNmIninNQGqrXi6Hxk3pzbjGBiDylgESduQlJ5i4dSLDO2ovfiUsV
VJsu/M8yhYYjAK/EA+kHMFgoYhBfQDTGNSji9Sb+IUf7zwYu9EQr23s3cA4n7JfQxbD55/KFURry
+IHa2KwbXkzA9jtVWIsGXwWqxH/6qr3pw9vdbE3l854GGHQoB84ohrEs38Cr9VaaUEJSV6+5VaM4
th4Jj/ztO0ZacFMIuWJ/sQ04vVifLfQhe3mSdG3gzMIBEaV+q6wBmxw3NynWlgylknaVWGqeLZ0X
w+b+nVExGlTx0/LrXFxU4nBuTovSysFakmIGoa42saRsyfNLzY0pGADF1FtX6oFI/sqwJwHmGQnY
wTWkikJuw0Xf73SBJEiLigifMzA4xoGIAi4vKH+re4rg7HJ8BUG6NU3cxTq+HGrxCXX7fsbiH+Rf
GMqajfsY/Ql3bj4fnba5dAw9JwKFBy08M5G47oB1Qw87VxbP4E96HFtAAOIvzVs8/+zcwD4UwTVv
+JZsJRmzUE8OYkfeCZR9TDH+10g6m+dYjb21dgjz1HqrXaPpk1gTB31Y/gfKyBY+hVG+Mi1d+aW/
3E287CMW5II+MVT9F133T3dAkU9RhmonpZYgAKuHOVOP6uUO9S7JEUgF/OtsgAM1q89jcgkBYkQq
apHXT8yr9PcgxJBFRfRPxVz3xHT+xpX+uyR8WvZfXjI4HBPNeliWqjNjbfCqJ9YTTNSCCZX0ORwy
+aiWE7hbPCXv7uWqizmy8MPEd4qRkJRZ2AcZadJ/SVue38/H4ceVPOCDZcCN7T7v9SnXTKCKJ5AU
l9xwcf8FbAXag2EMqwGJkatqACGLxxq554Xl8ZW4giA8JrcLRnJ/V0jLPvoJ1YSix3OjzkPTxft+
cYcTidqvSulJe0oubHYNjUHkyb/0xB7meeff58YGewfTCMxOXycxygPekeW0b9W9eWAN/zrt3DNx
8y7HIWh3jO0Bz58ypJ8hQEotSWdfXhP3IGIB/t52HOVFZ+VK1rOQTy+O8m3j2qnbZ3X/ZBwQUky6
83FJJ2aqz3mEnLV5zPRL6++ChFlsfAFkY6Q6YWL4zOM/0567TGDP8iPa5qMxn+Wn4PfYwJUnHDw0
hMgnBPZ/PPVqcRWc4T+8U3UEepzeiUon103Mg3D4hQzOWYXMSSWBmdU8UMnLnSEruEZ0R7eeFp5t
wiPaxl4X+sHKjNjaQ/oTI8CfNdXUuBIwBAI9jjsCaA8B0vvYJY+Ph3qNmAs5xLReBCURMpJd1sAU
ZdouRhqsK9xVVZiw80dWdlORDq7F7Qc4egIA9n4Gq072vAKLwwliXDo0tOGKKYuaCvWbo55mr5GV
JyX2JUdMJToLdcQUdX7wYWz+EeBRuk0jgGIf/H1GhU33LbqD6pMUGu/958xWSlOmaFUAunAYCku9
/Lx0qv5HyXKM8CAxYXs0tBYT5ktSOsQu/Szl+ULVqOB9a6FqqE/aTghZFIr+7ZFDemcZWCGEPJjA
WJvApqioES8jZ7tmEmZ8r4DBtQEfxLyrz6X92k/jocl+WOP5TYxzsDKcmRwpWUO9ShjZTRmKDIz3
YDkjh2i2r6YD8czw9o9K3UN6+Vmh7EjLU7r6hJ6PVFPZK7dSmXp02U0d1ow34cwdlaAg79o1KYJm
59tOIVu5gIF+scTJy6ze8rcKJknIgfxstEmdzGJQHBrTN9AT1sErvnEYy02aGTr6/9hUtk8aIBmT
GJB60Y/FAOTZhCynOOsTFR+lz1fCAGMvhN5Bnk1ZXMsRlfkTHVuoYi6GRyVjmVF6Qcw8p2l2Fj1c
UHIAAli3QegvS44U02p0FweEIwwvqx9shdyXWS0fM0FB9yvaH8xwmoOHtgHW5g8LnNjp0E+oSJb7
8jfAdJowDcLEnmLCzaVTGjxZVZsvyOARWxsuUsFiLAMXFvjWsLfTC8i89kzSLfyAfOCVckhiF5i5
YeOk9zAbRkeX2dcL8NpiWbWMIwU4rKto+lELrcG4GgeDLyj5rdwBP6TVKCAg/4pRMszeOJrUMQ8F
uCrcV4j6TURCiwZEV5nN3Jjf06QIGjTz3kSE+kh9M86vXPT0YOnBbMHD3yGF7uPmy1Re1r6K872P
daAxO/a/Z7phWLObqImPdtktkHd1ccagcIDNa7MPb0oTLsVPky4wJU+KfQ289f4I8fYaJypD9qU2
0MwAg08vQ8zo0tTHXOX+WyppKsRm24Y3LkQInR8fkXq5l90IIt4wSSywES6MXS37sw5TJCEplxWI
CBs8vJOxcXPvgZRF3XJ2V7sMqUYBAjAycvupnsYKSive/jOiJoHCy1NbI0X0AhVepxNVPZlKOL7p
keO2Yvlsyl+7dJv/USnXSjXOupWz1nxexVX6hKAcX6Twxl7vnm+swkkCriSRGgKScuNBw/4okHB9
M06+uwRESL9YZT6RlR1IS+j17UC1wZvh+v8Hi1Vt4cLR93NnoQaabRc7OqDCUcd9iH69S6ZihaBx
05xSLIBUNDC8/WM/76s+5IAaA+1PJjnw8bb6AlWMzQAhjdGrg/y68b6LA4VLi7c5/9yWvhJgYyFR
M/js/SfrHNjDZgL0Qm9YEAQ2rzPQGlpoVwAK9UsNQMUCK85+vFJT7H+yknh8bIfuP/pxZuHtdpqN
6+bl4XQz+kPxs1JcqY57xdE/gDt1lraiMQYAIUiNA3de8gdcIZoVpT9/f1vhF3C2NmuPs1QiMFp5
33IzVvDwo17dIPb+jNgjUrWiK9LWAskzYf0SzFfTNWC7SdgfqH7p5bJ7VUTavPCS9efYLJOy5Be/
EQ3rBlCA5N4D2GokLKrBMGj2WI90K5nrKIgztDy6JQK9CKGRbak4Q8l055cSF8m0cqd/zxSFRqCJ
Eiprt+6Wgqi8Sep2kaT40N5vzGjM/3dG9JhHOEd54nrYRJqLLwtb5S6nWEEQAgKEmxGLC4Zf6Mk1
HsTiqe5oI/wrT87J83ibxIMVQ+iYE9Milnjn7vSgDAxsZ/+q/mYfdyQlH+KXrDZ3pv/cgcey755t
Savf4lauGOFXja9XXBZH6hm4VeyO5Gt/XAlwlN0BfrTA3N9l5JtZVFN4O0JdtiVKtcgdvdQaNzNx
EQgZbmpIXlRQSnffWSdovjRCRGyeEsVXGUIDe4nlRDzHSfHhRfxd2Bjw5/sXMvSs472hv5ITRamT
vu1H3cmJQDyk/9/9xJSBt2RVwEKCbcQkT1aJAJ4FykcvgxGroKRp0g4U7c3itz81/OQS/KUjCr4/
0rLirtxLsAl9m/LIxOnB6ovENFtiYBcj/I/8BKT9xyoUKshv+w07rwV+CdSdKa5kw6EvRJHb2RjJ
eMhBF3A0JaxpbcbqdilaIkRX58ycQ8vcEhTQZC1OmyRrAiQXCzfa+RwovNfRrAnrBXz9pXcQ4C4J
ARl9XlojonG91eMqShLy+ISPtdpd0sLcUNgMuu0ARmHTYAojWODQGyxF5wABOMNuu57h4KVFcHiS
5VRGnUQvJB7bWVgTJwrbq4gY19rbvcYudFb4kiL0ywhlKA9MeiFwshp/AL92pgt6lWrXPSgyiwja
tGLt7Ej44HgX9cE+DLlje/hHwzZlKlLP33atPj0HeJQ5wqXFFLfum8sYB1fqEVp3N5jUItyN6Wys
XJcogfJKv3GrB9R+odveiPF3TrTuaZKHRRGEi2ZHWLTE/+h7W50WEDTezt0Kc6wwxpdbJSdo5UVf
hLmR0lQy4yy/d4xxjwJBKQ+i1LSNKyQM5Wi44dnajUqisG32h7/wHwAwkuqvu9ekVeasw7PdVscZ
VAH+DiR84qBAfqjSMfdPsuG2J2IcN2hbVuOzrkG15BDi5RxK2WswV6h9KclEPBqdgWNKFH1seEwY
5XhNPYZAQJuWAuZCGTDtgLN9Shg6neEOjaX60aKVkGYih5fV4uV9ufU7PiILwpNeIAgBQLnX+ueu
LZInlTR0e3IHaU8BgZoLJ90jjrl2EQhxNBQAGIMf2TKjrQp2eZq8YiKYldAqeoksI/9kA/rsKemz
TuX9KT6Qd6qmJ0BG9+ZxujN52yBcx6Y7oApYn/x0KMVkuwRZJsqP8EmPrX6ZkR8BFc74N6dLP+Ui
mu3xhaUWljh81jOyURM3BvQ3iOetqtP28KBMjMNRhYI3dT68znBLqYaVJTzUZE9KdERkUDUZq5Wl
bcBA6xaUNbGQ1r2bQpCRY4GAZY4tUu3clzYjpzAwVFTCXAFKXYojipJWbQlAyvhX9Jh9A2JcuK1x
PFoIKzxxEMd0GXzGqTOmCDBUQnDKuTqHIommHp//KuX52w77C2/27OLnTuDA5k5YZsbkWimJ187a
kdOquX5b13wSUxq/YZ3yhx2rk0HlrdDsOqV6eZKFjENdeGsvCLD4Pq90DM0NzApERmQ87i2gIVSN
uLz53d9KJKAjOuKsApK+9g0zVRuRXboD7iI5BwvDo36J1fPSspnYpwOtcD9ACpDHLJgnwXH8b9bJ
V86mg9UABDMzj+CKcG4PJnbHZLBIESIgHugCyVM8CfKLkm0wjYkBNu5UmYoqTzGQOlDAyT7VnYdz
0lO6u4gxE7GG4be29+1qUXqo9b4uLhDSWjjawZqWbIey5QqCmi9O26VROhN3FjpxBkqL9DVi8a8W
VLS0R4+hkrwIAkeG9YwK0QA/g1tmsKEWJDIX10lDOxZx3fAHHz4WNHUiU3+2PNGPx6OkzEQjA/aD
U+JfvXG4Kqk6RT6PKBjPU6dNuRisf1393QLXovgo7+GT7lTG9dYg7FYPQQU7O2ajC4nRaGIKkNZn
UX9/x/Ls3Zu/YWh+TKuVnmBLV2budZA7ljW3Vus7EfMKv8GvP6A2VfvxjVvSAB0yFdQATeTslqkL
toWdtHE7BsfTK9daGeDiuaI5MtBvHAcMlZSPJL6l/o5ZgJs9+Lqp78GhhtbeAAUzA667jUA4ZfD4
dkOEntFFx/6pIb/8ssEek0rfO6M/lhID1EQgIzZitc3bpk3Aoq+sqJ7lcweaG4GrsTQoGWWNlOex
lRhlFVv5fXEmDS/jjZcDmDOE/jVWrKHqhVWHDHcEp/DpcMZx0ZqIN1X43/vVtB/cBXEKgo93PJFN
2/uFAQuxKnGrOii5TtiRcFP71M+jtioTKMgpCP7WrhYZfB7YEfPOVSfxwjZ2buiKYMFtTd91pdZf
85WDcuKrc0ZFyUV/ap6duBewh4VpBrVGyhwmU0TN+B+m5SQrPtR0nQMHukeeMUgkzNjYX7MbbVe6
TlILINKGPTJ70MEl6RJ1HAosX/s2KUXpqi2mQv7gjVwtI69Eq9BL/hHHGXpFTDCxnJdvW23veQj7
z3PNQ7NwH3OXVP7bI+UD52TCkIknUCEDL1p1lb+fhqx/mOoyO0KsQblJEmB3hGjFHdgKzBtU1ZMY
vrZc7Fx6YH9PpucB6JnUm3zJSA/OS8mK2vaG5DKSyZRf3rmWhWL3O2H2/jLqplMvEbjdhI58ugI7
Xcbu2De3LkVx0mtyMyTnVhcC5KI/1ealsi/xoQyCI6pBgsNE9XVCiu1/rXM5S0MqojGURMBvkV4I
QDxM3caAHgSH5oR7ayPUI6Z2Xp29X3KcPJKcQ219+EYLzXwDZ/JnC9ZOVtLf1t/k7zHxqEe5OSJJ
sPNfTmQLi9es+06hJVNhR5BaN3+3S/5GmimjExYJmw03NGwEooSR30Hrffdu+2LtWAWicvbQO3xk
rgDeYE9bq168Y/+TG13+J24f3DX/MMlR8hTSrzbLTEeguuUhBbXebdXFvuCI+ByPATzLXGkUxgUt
t9JMTxMB8H95Fl3Tinmn1unSsJkfEWk7DUohxH7AW2yP/55Ia20sBPoJuBRD9wHb/sJYoKxCjLyl
JC5bQUpucmPrfH65bxzEECjCfmdNdo66ROUWH4wlmxX6nS9rVOdkc7itKsSYdGg43sT3rlqm0xPr
Pn8soPh64JEfZyRdPPa37XbU8QN43bmI0+QUIFdAaqS4zuqivj0lsG1pjNAWqaXbLpMORvQ9T0H2
G4euyiksIEBaEBrgllU1LPEZN9zYV2EUYW4BSFMM5GKKhES2zCJSmKLFSsmzJZmrUPXLhmAv7H0d
6y3rqVrp8JQesXaQmUDWKQeFGBc/vW762ilBJ/Sz5gxowrDoQSi+WSSTi0XMbNiJLF+fJvLCA+1L
VryoBrjS0XYsLywqrrDsAB04TOrSXWjDtNVgI5weAAE8MTQ8N2VMcGNNDD+wg7R0/RKeywAAb06Y
vDstwWTxG+QpWK8NfDM532Fh2HcTBtJEOKqYd4pddIUcsPIOzKnjRiYn3huaK6zTZ/9SA6c1ZU44
RCBOKoqagykJhebkSPtuPMC+mXFTR4ZlzczhAH+hckMrF7dWlkLby5ru4SBhM36MDvGokoIwMn7r
41UXeieeWemD+qty76L7wP8sc5kuYprjViWIxZPMEB+OfF0/ih+eLRCxxPJfEFVeuaUkIl5z/QVq
Xte4YzwgNt0RPo5gSRiwo1+Ru9KRkLDfxNH/J4+4sX4yvzYB6zh6/ZUfqMjVbWC6nC+DBCWnfyos
Wq3oE7FyabIEoKT73YLZsbIRiE2o2OoaZgVucaIGQ90qjenRwYvDI+HdCDIH+rrTwP9dbVyyQwWC
7iHyJLn9Xf35u4v/ZmTDnJS9w+vkUuJXw7kBL/P8+7qGmkn36GGE5auZd4JI0XMSiOCsJEeqfu9p
41aZObttvP6qYmgYc1Gm4W2cN9tBn+QU9jYWpGd1UXTVMpIsTVE6Mb4BB130rpEmXlOrjOF4FPcC
lgA+wjjrG2Mmxkq3HBQw6sTFenIgkrHgZrGGuA/uWnLZ3VrdJuBeStg+vcBjWlQTYAupE2Ehvi/3
HB6wmlxX7NZ1x/i5+Vo+mf7SuiHB/QXBo9OlSehDTCFe5K6LHe0AsQA5lALR2orGbnJIjEISThc7
Sj5fwEWq4eWvVW/1CULUPVDei7Q6Jn5rLjYeJ53Vjo/R+iaC5+u4gICrZw85hzy1Gd8EinfaSPPS
KWphc1Tmu7h7D9GGvm5fQu6sTsTWl8x1OCJIS/uKhf7g2/g6pEQhl8a8TfR3W3Dn6lxMvDDnHCtg
rcjFR/MUj5r48cbTGcxlzBQFmxjjRRYtFmnYspNg+MWnbSTNPR4Yry3yCcdaVs2b16UNP+xu6w1P
6LRc4Uc+p3IRopgs8UHX2ZdU8ZC2mIASM+cSyA/XakYylC23eUvNuibrx0ocVl+PImTQDH0q6pZG
1AgVtRHX6WHiNvkKKRizReFb/PI2ilT/2xGjOGs08C4l4s7yJmchWNs5xmqKOwj/M1YICvROcdPZ
LlqytrAjOgqOLwrougGkVgqckr54OduYTOeWGKiJHEAbttJ4F4oOrudQoID06mpOR8JZITF9lz5Y
5Vbsp3/X7UvPVygNkrI0kV+PHXtJPTl3Nn91egOhRtKhBI/LVc5Y74L6qhcJBD3LUAH49Jlat2lN
RQy5ibyrqw0dnfxVIW0Gbe/rjOXn/WazPxG9Rw4ST3KRrH+DOU8jLfoGe0oXt+GEj4iDNKO5YOjP
213AY3ZNq5ipt+b4otfw3aj/Ke+8GTgCypX6SLTFvtAnca3Fajp9AV7JoKy9lEKJ1vpAiMdSTWId
/wd4TtDZkngxKPbSQOOvCgsh3t4sTtNLrleTdRNzTPsG8GiLWgVC3fHpNo2px2cE95O/ibAcY1X6
QaZXc1CCMtT6beLTTYmw3GAES5ReBu32+JEjY7dB/kFCkeWOh6gyzwnAekVMW6t+6ZL3sIBQfNGc
GxH2ognQbNpnOiIOyidNz+DXf5jmGI8S05CTXLr1uAf0lg7bYjcqtRXn2ksLfU0oEcwPkBEF6lrw
VvAI5dTlBE174edlGmR2IeMiTVEYUqUQW/A7dnkRnK9Pk+6dpsv40vo4cUPSDoSGBVEpw6wxoq5g
D4TB05nxjs1KRTi895P+JL2iykOXZcWhxaEMM9YHSj0tRfQ1a36L2sUJX4m4wtfyrNbLvCDbdlZq
ynDwiOJ7qB/yYo8r6vd9qp/nAdp7yB8PiIt4Pptzofy4sHvRhjfi1f3s7+wm/Kx9W9r8A5omedsI
0Wc+nnLdKBpXdvTbiwiMHd4QD/JYWpEWyNqi8P2lmP8Y0w3E610d0H2HpSQuJqexmxM5k8xviN8/
vNH1fHiIilbqONpm56hsV1eP2WnjmZElQLLOxx37mFny1s30CwoGIItAT8nFOkK6ELjAcAS31l8J
pcuu6LpuKRggU6/eF0qVqOArt/xpeQ3woalIh6eKqBci9Jo9OTZR7rnU/mD8sETP2NAoAgPsSHG4
hai0thPIxROI6PYY0BtP/kOrJjjtmds4QaRgGjX3gw4Va2yjfhSLXGekEq9WCK5XDOxlUtfL+4J7
w5+KPMfwVVEm9bO2kjmBAgk/Ds2ZYX8uYkrGAwjerpnGPk4kX/mXJQqTTyjdMLB10YDP/rejnNxB
2CZ9yr7xjzdJhT6eoku0eILeXitv3Kwo7+ssXRsRV/QheqM89aK5XSKe8TXCBq2LxIeyt2txBUtu
VhW6ttRxe1k5DB6IYV0ClHIWhJc5PXjpczhwW/HVwKl/UJrgVTx0yVZmZ8o0PksKLik2a7wKbu7i
u/oPIvbjSJRwCLnyd5X9u3XWfWdtbXXyPpUAwuwlXjKCOQqh1BiWcKrWQU2olXSXVgG6AfJchO/P
M6O0yR71UxG4jW6PI/SVI68w7srjaB5FBm9pfK6wo+F+3UCikdQA3pSRqw8+xbvKDTDqXXqXRr5s
mvOnrTJa6fCf6bMxTvm2K2bGbNQrgYwkOJjRcC3CpFaKX4HbTbvGpkCh1sJ0BlUxfIs2oLIzONsX
6kpT27aBN459U3aTHLV4qqOOivmJ+xY6VaHuAM++dxR40airxoC5T2Bm7U0BJrICuCXY5hHcOYOy
I2fHKFS2yDil8OzTC+bHk+eMjbU3IaK0wm7F1ZHwjDITtBNXlow3x4OtcQ2VvfQVQrL6hQwh7Kn8
Lz6qdBBCN6d5lIGYyybnQ5I/C19lN1HLM0rECifxdBuim4UVUffrTkB6An2IA0+e7Gqdg2+tf1hn
iEzUslxV6wGU7vSg2REIZyv5fklrd5jwjONlrxYCPOfOGyeATUzjOAOrS27nZLQMpD/FTsYAuHSO
vNtGPas0G6INBBuWdDxiZR3AD3NaqzPUU2OKn/EluDtJ+OMRa3EGIelHgbUbQby5GRlySlTAIxtY
tv8t4DnVTdbPJCk/Tmxc0GpnfM/7LeBNncfrZsuqWm+gJws4HflFQfWh8Amq0hKrolUkGwhBvC5k
UpdSzjLNqKiUIZOvcToG0eugMM0mxJkTzpeam//0C0C+Th578meQCSklMEACGGrKSswpzx9nICSR
Ox1msPegGwrTCcwAuXxcBOpPLgawv8JifvY1ZwSH9t5DP01GQQjHS1DvtnewwCjDGtPjijs3Hu21
/9HGD820xdjpfsb06I2xR7DKSjREN2xMeDJInr0rcTWFqj6w8exnwshH0ncfckzKQ1DteCQg7v/R
2lHr4DimLXGHaMv5hPo5z5463CsPcExFeSzyvIVJhxJDWrBO1I51rZRjk1aVkRQ6eqZQ0zkHwXh9
b0v//os4OZcTntu+NjKwEKWcJUND00tb4fCykVmzdnsOgw2OzAzZq3tMmcrqY6nBuBpTD9t6D7BE
ENNYtJUv5evEvpMS83hU7x9Ub2Tss/lO/LZkd48ONVRIFzd2TefuhaKPUgkE67VkGO6IILZmCjXt
G3Hieto93KSx07wdV/36yTX+W3U2lwZQXWRgwOkdP5ll2Gr2sjw8vZ7QE6xr7sMjWSnsZ9OT+E/x
YClGmrZH/4yggdr+Td7TkIlYkVKOthTfcNKlBa04UnPEbdNWFSeEZSNnWMSmeelHj3HKLQfoOklB
ss265YlNriN3iBWvXBK/u90c5h0jWKNGxSVcK0Z3d/A3n3QWjfC4ZawHMlwDGMr2q4UFJUMkH87n
kMkmA8MjnEgZow6sSMJLqoSnc6ZxpNE4Lsgp1SZFiq2iQJMpvytzao8tKNdfIhiNIZYuHdcNxTNn
OxrnX8DQ8GFPxSU+dfbIAGAYzcSU64s4RK6ZFwnUZJlxmmbOwNA5dh+hXq7lS86hllWEbp4zrsFv
GCDZ7n+/6Q3jVx3kIJqilR32VayGJXFuc/kvXqTk2MjGfo0dsRjlOUyauzsOtc3yIL2lJK9NCGOG
m5FKlBKSuO+3Sg/yaKr0JhUWtH2WYj70mGf1u0v1jxVqYp79PqSZWvGUICDvZhpmXFWocRy7V4Ix
wv8rIoKoJDcmC8G+CfvE7DAUgc3NRR8yG9izIkElfr0rJNDMKGBYaKUGDDGLWfa4hD/qoTa4UeN9
ZK5QgiajY57B9bEPM3TbgbV+OQRMAFQpmZPjRDdFrV1GjDrXPgp7ZezjJc8Fj4CZAnN/JiLyRHi4
BTUBfQvgCqg4jSjf+MOlzbZWZ0H/9Xv2fR4774WNUKjOXf5xkVqDCDjqjMWnEm16asriBEuAO3Pm
h309zbxwZFecWqshS3xzIybyEcHBEXgtOSbaM1yLhkIiRSo1Rl1Jz5VdwyCETXzgjN4649aEtbmY
zEoBhKPkVWCFTtVgjhC4/ptJAKeQrkweCfZdtemVZ1+2/j1TBwHBx3kH1ObWKsD4kTyGCM+bKwMN
XhgVPbyeMOWyLG50mfDDQSd4fgHK3SEocsNNkPCbMVlLir953VX18/k8FzuysTad1G0MYIVi6rQb
nZrqNnavvBRthKnTxrexbnbzLpiaRFBheFRJloQ28KNYLU1IYmTTPygWb/qq1bi1qgo/KCX04cRa
Mmg73wqU+iAu7OZa96fvxZMzCQ93ogJZ0o9g365EW4ehWPL/wF7X4dV7y3r9oUe5noBCcehMbI74
LWxTC4CG7iIeJMAQH1VWctKj6z0oW4XBCjktev7Ua8hfMcFl8mmmZlLX3jVhY40SaLv1zWZhEQRw
rLE3gXCqYh/0A5m1H70/mLROcgZc/eXrSVm/H1Cs7Ka0xFGfyuy3Gtra9xFLLAEvA84bpgGPQ4ty
vojN9QH2g8wD0egEe0aQBD3Xl1rlE9642eDNfC+V7FGXiEQYn+oW2toZYsVop53ZaweY7Qf9ivP1
sUxeKaLuW5/Fz8JvL3XZ3Qpzda+1+6ZOZrzPQl3OhimqyJh0opaPlmnNxxECGIKzwZlmagsk2H3V
EJKjHhPIHLupPc8j9yKyQE2UHqkCtIqkutYY+RJis6OTpHtI9dub3+fFhbDCWn/a6WZq3JFATxOd
jLrMQzVxP7tuZRKPQnOsk4JSzHZJARhdOGTmLh501OBsadrZKtKTXq4b2kF6EmkB0qHM/ysaPVs7
o2KHHAQfSwjBHNatRrq/Fz0P4OXXg+KaeFUMcAjwphAOEONF4BMtr15KLkvfi0J7ehJd7CwSkNT/
lZyr2mllgeIWLxocLwQ6Eyq6Elod4NB9D6Vm3RYYmekxywukp0UoGKQKrZ2LYCXvMVHwjsDJWZ7V
rG8y4zV0kjvx58J4ARhOXrKOn+8CPUxgsn8+HxQgxXXt6DIL1IyO3rSD1oHZWrGrobRFZdUG8+/p
z3DpaXRoPx14adjkAM/Fxz3y8NprRgUSXPdGrbFYPEoQJ80nE3pvKLQdkYJtEoPkmV3Qae1LSBUH
4iQ1As4qxrY1t9N3eOCHc0qRmZGJBjkp1qZRHbNFM8ubaDIZv2ah/8VTja6qYhdOVSNShYD9ZLgC
S6tu01JBpt6Z9OVCVt+x7iR/1N3jfOu0+LsP6NTR5eKH7aIcoKwGu0gGchuim5LfIdlq/vjuCajL
4HEMajVzbYwJbDYLeMnofm6RFXdg4z6d3bC4Z7oDEce52qBrKd/Sj71MX6EpmxO/KSnQLz/RLCXt
tmr4l4ZOsQcoXdBDtaqaD3yUvURWqK9K3VkRgUBr9HGVvdxFtYple2qQTBor+D2v1sai4E97Qk2y
7MtBYboaYGWkzuPRa5cdqr9ekZaQTzxupGO6wCZgLhH59J88sYr5cuIUwNZq1N/zKpGmdTTAUFpx
wQI44DftWZE7qSqWWqlA5IvQ2yUWuSnyMhnZeecuztZh1Bax0QkdDaskIAiDja/RAqkACg6TtcXt
iEG7g+WQEuVfDOuymN9utkurvIvQC/MTZnwB9akpaNUqN9kTPtl6syCAPJNMfhQXNSGHc47DHLSx
wtHwzWCWCxUzsyf4B8JvATnrGdQEO7/qq6in0O9EUD+4iLOMstZRQvzMnr9wDtM5LOJwSsLvfkUh
y5MSxDqSXasdvcaygiSf03XIbFLT674NR32STyG0WJXXRpgAMM1pFXekA145RsSOHreiusi7dYlW
WWSeX6NZKArXYeW4kEXPQdNoVxnzEjxEte4PDi8bJms9Qcv8oV+chJcxsdt6ZTKFvnwtsYHjv2ja
4Cz0meJFCReCZz3rd4kPM95+v5989FzRIEN3Iz/31iKQBKMiMAUQesanzFYWiYo5vZnpUTABKbY6
qn9L8MhCbTgTLMQtCArCKl2hLv2Re9udrnmrkk7bWK9sCUJG9xzI27QxWDslMH8vGZ7m1ltBri7w
qfcLSWmIO+rGcsc+W4SBgmwyXWGhvVHONBo8vzZgqQR0kDr1F4WJzMUVIyn2T6fi0k7N6OlOqx6D
0euWpPhLm3GDtdX0muSpGDZ0tC4r6bSyA3LraevVN6sTUb0u5lV2Il44I1RHOhXnH2UzDf9/3ZWx
HED4sf/yUaE6hqAbJPQFGOA6xQg0PBqJHLn1Y+gNyZ3X5OK/ibDsy/hcR3wiHz1EfonnmbwU8Iwf
Sp+BSqem3bbYFTjY5uQFjeo96sqXrk0eoHvSf0ur54YRlm1UqqEQJF2v1LA5ukkWkSrAWE8+YGVj
Rppawjv9hzbFNUXX9f4hmf+FrLuP60mdlNxXgCYDy5GoXcYVBmb3KBYLTbP7VwXstv+oX++vNGGC
O/obaBkk1mO7KCspz/5HJrpobAcPDHDv/uO5DA55kN0UROKvgMPZ2Fo3NHcfoP/BhMuJbISBxHJh
eCFyYgf8/8vsgUFgYSdw14d5sE5624wKBNKM28s/wbslscHuTL3z+bKEK5pY3uhPNscciC6d93xw
CL88BeBl2pQ+rCMzFw7E6RDJfs7mJshDsFT3TIF1v9Cg7IrsSUwnDEDZerD/As7jiFLEqtCkIRit
X0rpDWHCgzlGaXvNLKjjDRVAHwPLPcFI23O0yzIloZG4vrvT9M+6FeXAo7C4kLB1qmLWXN2ONZEC
wZwlyX2R4mY63dg9pCE8A4Odcq+Ebgjq9NPCfH6AZcvrXNcL1oPJIrhA3pTt+6Ke82YoFvjkQiMS
bv+WqsTDXUlPtdAnw8dvJGRS2W7X+AHheV5J38iSq04/Ozlqv5mo56Dyzb1ytaQpgiDNG1TIBv5s
hvU6bwAt7bZgdQF5Y2knDDos8nWMXA2Iqxz/3vNYrgu3SlRspix2GVGvmF7y3D4eD8w4JkC1N2cW
gnT+FCjA3uOb6D+UGdx4oqupzBAU0vMR1VGLzCI9csd1KPXX8vynxHdkLdkdQfN68CmdM4rqukjw
+GHwpACo7HKMySZcizGQmcSwj0mL5q8tfCFuLsh1aBLHvKVdEAnig9ZFLVImyVtpOSiEAAZNMom+
7+7Znd/QskS4aL0IgZj7FCscKc274nDtNF/O2yxcgtTjwDVObx3z9Hm/8hQJHdf4rMe68PI6G5pK
NMkgoQ0Uy+BgsYBwBK6rNxI5ShMxVMsZakTnu8IFteCUIFv7qc0n9OxZKxlXTex2XeXeVenUPfCz
SgmVYq0dqDJ4uc/cHGxAV1bETc1iEbRrUzmFI9eQtQL6g75iJz5yjlnZ1f2mGsldvw05VkQFKfhZ
hxrAkywJ8lfyBwztGtXN7Krs4vkLqU2OZHD6dhRghd8BbOduN5dH5LYFlQa+jaV/jdXh1zeoiRTm
oUs8cu4duV0PdrsmsukoNaBN6St2SmohkAc9PTMpJWuJoLVyAYplUffzGSXVldyxJkh/gMEj7Cp4
b2tCL7TPDa6ivxiCifOafqIYAHaW7DD3AW4FkLdMRqY2YvhCSRpfYzQLIFHXd1T+n9fsUiKMuXyD
z37tlZUcuJ/1nDJj4rz507eHA1yuo5AK91U7VHVesCpi5XvxOfLf/DHbl8kP9UKaDWvCUSJDoc/l
9hwRTKxSFWHXBspykjHjWmQkMrPf2N9PLTt/X9rATZ+eEehzy/TP7Rnb1UxL9uu5rBfWqWmKQO/D
7iMqkuTC6Gv+naXN1BiJivgRBH1j9qJTANiHYWwAfmBEWXujmzTxOpyFWx5LzIa82FlxBmBRmyab
PgeL6rKQE4a0P0+EKKzOwYPsJespEujLrtKCvz6UXc1IgxiIV8nJsEI06Sb8QEHH7ULcyuJbz7Gw
XqV/SqWqhTEXdZgFFHrZnvkMtnjBEcyegrzFJhnBwwbmSfdeXqCqi5nX6tXNLJ4lT3enqXShya6C
Ju0tgKC4GFKcV63SIuIHvqj1oba9Rx4qIBdAZcE86K/6+hGQX1XgnZ5cRP2qhj1I39xI3DvbBXuu
mpaWBasc612wcmmiHeWve9Gq/4lYy+fXLTbbbKX0d2ee+ECNZCdvdXOyo3rH9XtmB/PGszKtqHpV
N6bcKa6kRrdUFvn50YfG6o7fpPX0rk5F734JmEfNz6FEFKYAljV53L1bZdzu540RfS+KhhqUsbM+
DT+ZaELyFk4RL0rT5qFZ5bvNK+IzPCKRmD64RxM9Sl7lrk3kg7WbcPAH4Atl/eCjwBJl3Bxj8fY/
HZUC+q0GPWcvfba6wZGv4+LW+SVT62GpHL7LaqdhjwFfqxRoT0cdhySV7hua2dR9uKP0y9dh1LBn
G1vCwuFG0/VbUwk7z/PaQJr9mp9UuPWuwv2yo99nGnqfBNIuhEKEglZxfh0w+oWnuFjdL/UCqI2e
D7ArJFkpgK4iIRzUbcYky6xsTx55FlJFu/hV44t12R6opjw0MmQMeSPrUfOWyqQDbcmwbKFCGSTJ
Zg0ORwR3y9cdyz/1U0T4CRVJcrLc6koMx9LlxcwrCeLSIDxGiY3IZdW6jO+ZZkKVSvh5TTk6//5D
RG+YUCPVQMgJyU4NsqsL66CslkPEZs5s1lzZNKO+I0t0jKQdWtJA+T0HwLKn6V5keffT3vsWKZLj
SW94sEzdLevimi/A/LqStxxpWvg7lBTuTPnloqYqYM9oo0ggoeDSlpXnAOZfdD7KScX3lIdxNvnU
WPFWkIpD42xQeXY5AQz07kcz54/gXgFvBCAz0AYs5JzRoxQpvJbrmaMyuteSr2SwMWHGR0LwHo7h
4ycMZI+IsYaAqGcM/2mh39ypQornik8GvbN1G7HtG52y/Sw3NQTsPEkgswoB92o66yBGQamBrXlK
SXYTGajKXnxFd5ICX6KO3Ki7fpA4ebcuER+QL2tNfqWwh4xas3ODLNHhta33ygJyo9igQq4kVOHX
BDfQfPQVhdN8g4UJMUdDNuThl4VmQr5fbF0Uc+HyWEWV4b7JSqje0dYpc+Ij+NaZ2fIRrZ9tYeqM
hKgX5oU7h8YuEPZJoI2VISMWaAezgjeJvysreqh0LangFcd+lvrBK17hPXa+rT+zoEqOP4jHagUu
9fNthFKR6cBXq+h33bHDyHGYIsakmee8PJQL+2TZbzoS7lwD0YLJ4PkJ1SuULxx2a9fuPc3hE0HM
xeBadZ8WD80mC0wVHTS25LbNXMprKToCLTMMiEBWpxv3n+l8B5AVhDhGMA7mWCPMLa9l/hIg+vsj
rGR8Qw825/3PisThJJTlewfCMwu6nJTVkHYKcJbb9qRqNHxxmuNgz4795x6Lt1MsN9C2C+Pb0Dlj
2aTBN4sAtkPVJG5SCuG4hp7/TjZuopM5UG9/WrodB06I4YHxDT+S98SyHl/saf1qbmjx0ZZvusXV
1jvbnFl8Falq3gyBvOCLZiLFf4DHfBc3JKxx/mJ+JVOomSi9DyGDVINPYsW7q933gSONSEAC8o2D
ZF3yHjPZVH8StLfNvfXDIGyv8fY1dxJTvHcZ+tyWrTHpAuyyBSN+DqBmMXt2CRofUzEELiTp2cGm
RuNsINOF36h6kFAe6aVTciZA3RUiZPt4R8mLpLKplg6M8WDAepAsmSWRaUHNbqVCWERt7b/2TPi+
wBHT/EgMtPwktQlTrRNVU/n0Cv8OaqUnZDIpGUdVB02m9CK8Hj5YUpKevwXZO/kitW5ZtLmI4G8Y
gPkHYoeAS+r8z9/guu4F/E/lIf/hhszqEBoFg7ZzwhvHgpwigjf2RxovNIq4eydIVZ8G5nfKSjeI
n6pko+PRdY7T8TB6T214kbvkEIeJosweRm98Yr/RrJhd3cZfUbkjZseb1tTzEuiJfxnA8Gqf8Wxl
363qM2BJl2U7FZ34qCxefJilC7aqHc0ayInVW1905XkDYe5cli7DByNqTWtcF4WSLSPcwn4ae/jy
GRFL0ahu5thSwI74aoa9Bgf/6FhHsrIPysFpaZXsIqK0JoKnhaN+kuzLDFP9LbEQdIIvoHhuv1qp
QYAhVJMZxELITwxvPNJqmL7rgSUFHntJehlAIRlD31Yb1i73aXRuySnhFCNYYwTk1SH0ykFwBokU
QvlmTsA28YPJbp68nsQV1h5IF+X3uLku39IhIFiRFBKD4D2GDij0wf9q2dJqoVHG+YNICSt7bXt0
ukhjr3wVu26dqzIzWHpTBs+JR2YVN3CjjeMLXA0wAJKFpHQshykpp5/om0xtqeE8adDRInG2g0VM
4whRxbnp19edtNRJppZ6C5/i+cOsWPBGihvVt5trYEECG7t9VWWPpW8vB+jiGJ1ff/hf/XPhfzBV
S2MMHHGKPiFDiyAaipXaVH181i18HasQauhh5tzuqv4+EQIakOWDtZsVgM7ej3yIvjNAv56l7Mt+
/KVo0z4wdKJXYHRp8/lT3HcoMDSiOcrjGOzjK6sIp4jHUzbxULlTU6qZhaaCYPkh8OZLOqdQqBMe
z1s5bgJsKaWSddHUCamBoST+pLxQJVu88/VLv5HDry1bslAUCzXKNtcIEkypNQJzirQYzk3OH9fs
NkxaLGULbp3BXvJJhj7rjuyYD/6x6AtgZu9KyRruq3eIDkB+H6/BP8wK9xWYXRVwA1ur/1Z455Uy
FsCZbudSKw9Ia9gpIJ62I4EUWI2jgGldjJNoU5CpJA+E8SI9ab07cXpE+R4FxjeirkKz7TltvuDs
AhKzAS4eUn7NSrYGM/rE0Nt504wdwhY3he6yAj2zxXL/Nh6LqYCdzPP7otqh9OJqxjv4GdiRhHgb
L6MQ6g7/xmti1LDCT3Nu4E2mIkXjwDK9Jh4Jhd/BfjQFxcdHZ8ZNUfCaBk0z4fbddHYhNGtt5iXo
sZSDhakVKwalN3cCIAB8oFIvSqcVCIX2dh+LoM7zqZfmmKktCBUwbXAvAlwHjEgWWoWa4yrGLvv7
h+S3e1bYg3d0A/+TQ7tvSSdGHBOnLMEvQRNIJDAIpGhdaruxeEC/kwJeGD/mAj5dQu3+JdMoA7gC
/JaOtb51uQChscl4nMKADXQg5tf4s2h5a0GN+nrUVsR53nKJEsggAB8UQhzXs1dQdrd7ZqngIYQ1
tXv1cSxOPkQJ5+tH7IQmLgasp8IOFTPHBbgacHke4iJPKsuNLBP1UzkrkfeP0upCm2EW2q5Valow
v6DaLqcVvC+q3yMv3MiMEhiiIgqTbnt9hC+1LfJ6R11PYb8qGqc7wAuXCTmqT0W81sl5baIZRYPx
4UWSL5uo1Tzcwgv6t8XH8sJXLCXDQI0p5hYIGaZMaApY5EVlqMYM8ZC/WUnK3Oov3AKCySh2KOHD
+AorPkQYT8PgkYKCWlWSNZt4TaMUQYZZ1M0f2Yj5RWPIELgjQ3dIFK92tFuFsLMvwfc3X2GC2StV
4E54IW90HuxabJPJxD9/z4Rouesv0smtt9VR9Ha50c1dB1D7djtKO3Ad/jhWQK68IgGwF1C9eYmH
m6A1DQjFYb16KhZ+TGm76FCe2z0QFjIUpcVwFfWtDlcJ/v9pkASlzaK7JUjgbnxvNjsGH5Zy3g8f
4MO5bQw7vbSgEQgBF/7c6uaXZVzklwu+SX9DlQ+rM9Q89GYZCq1bzAQzBsUe03S9NTaA2P7R0uDE
+ZHgq5vuOBZAWeRT5DbLs90dSkpzvnr2+GVAmTkJeu/ZY0j1jYVkkc4wq/jpAB1ERLw2knFTLAsq
Jy6wzBbMOlvr76rjcdoOdn/5O+oUezkU5dBiKqBVOwh61KDXmlErFaoKA24jdN1856BFRzR6Wdh1
pSMR/MYQAIksc9hHqLyei5C2Gl0m0Giy0+ZRCrW+rcdc5pi54/RJ1Tlt2OJfW/t8IurmZ0th8gDz
hC8ZHWwhvXeBtgMSTnjxIuajwrCEZLHEGKmeCGK8SN+RdhKrWO0xg4R4ZRQDKhC6TTMf4d6oUPJ0
W0ZtmJjnB4OZ519y/icy1GAN5Nn/ve3M+XpQ2kNA8nn1hitEhOp5HdwxbO+/jINxN/NorvnAuyOi
GZuw1siZQXrEkHjRcWQS246C6ufJJ5tIY9gm3vz73spHtlyieXSE2ePpHfiRjAHlmJLgsgHo7XkN
EZtHWCtFSGxIqrOLACJi9yitajqxNAAaDRwvufyY9HhPm3nCbiU7kv/dZV5xoL0jFXDxpw2xm2Eo
dSPRJt9aQFb04LvgtMnzdvmv161nFQP79z4aDtPTWZobvbdlWZgD+XdPlfrt6LPYr5qqvaIfPfsP
TjOtevc02vAl/VrKO798MJozHSs6PO9hnzfmNPydD6bTvRgqElYeFmm0AL/COf8TsGH19Qr56dyP
22BdTKVDoUExe135HFCvlz0jL/pJyZ0j0z29A52qaG57yg8t7YTamrfJSyY/cdSPujbte8D0c2W5
m7RumwaEZdIZI+PVscnhZRzwzVDq9vT+g+9ytBNnVOYlrlBF/LEi/GO2j8e400RzPU8Eaw5XHf3M
oy945L3ewt/ZrrEQZ8XUyDBALMQw7kEOCpo+wfJB+61L6KIEn8jFJXPJLzfDqDUFSR5yRM2i3dfr
QvijBxZI8dIK0kUbZmUDWmAG8aiv7k16B5ftV6pyAFFwC9kat/i6tq7b1M/XilXjevDHoRFa6bWY
SYcFI9MhtXoKW/4B+0Q2icOMPrKuhLcCVagO26eeAXpEzg8zLTl0gRYbPhvSqetnSNyrCfoQmWMz
wWeG40gJ0ONkPrfGJCzLVzbVppZP9X792yXn8IcX2FSLpvkF093paT+zLdBva3hrrnyv9r6OsCoW
XX/6a1Ib53ewjzqKtS4XVfcgC5HQdxxJZlzr6mvBAD9B9ROUPcMZqHPcUOae4cDWj8dvRWnr0WZQ
fbQq1FTSqoKtuIqObflu/HdgnMXdx+2GOEDONsxAbThfUzwVGn3QQXjhJhxmrBSf5L2gz/kaNdqw
SfyGlekxgD45rIrHVfEQ10u8wlHB9pTk6+TKNkepwncQ2li95joxJZ+k3jFQXnq88hIvEYwBTtjM
/C7DSdxPALE9zv/aLA9se+9hbzDklXx+nL4cUgcAaDHG+dDfYcFU0oMadoMrHKmHnvAai6blOXyi
deIGgtQHEiNPgfZBQ6wuzJ+722HJ1Thymo3pIHLGVKgrHSDVU3WjM0n9DaXKj1kmlDgSlgF5R6cN
0gggMwhzc/Sywt+vG/OtGRyGPStwPYvK4p9lz/sngmAGb/17BPW/bG8jRQDbunmYFa6y2aka70v9
1sFkM7A8jcvwZdoV1nOtVnzTz9Kb26gdckedmw9TxQlf1N/d1kQwSBJ+20dJUo0cWfFiA6mIzHzl
NmlbCbpVX2IjNfCjQO0PcR4JgAZkzmsHP755Ncjobexyve26GGZRfPtTpp6gdxRO+eqw2n5j8fn6
4MLJU8aRK+1CiPt4KTWvyOYLDWi0NfimDtnl2C+YNtE/OKBnWCEMjTGHAw7G0aHTpPhXH8jeZ5jN
GRIL84o0LB5jiP0Pvhe3MZ6bz4VDVMeNjCSUi/g2SrbqF9ya5fbLOA6UlO7tUt3JlVDxQXWnqWz0
U2bEzwzicvTY46MeTI70F8tnIN4una1+EQkJuRuNN9npZ7ZAUyCzNFd7MAeixnazsNcQoyP2bgxD
pIavT49b1R23wQeQWEIu/lU4jx5a5/uByXbvemqYO8Lk88wLx4iZODxPVe+/K5GhohOpr81xwx0e
XrLwPPFGo1uu0MmJ6hFuhVKgSyQBd5ygzayc43ikqqDBYZLfOfFCnkcZ85HvgtAK9ke+/0/GirVC
0GpNS6F3csEKJ/5vSxHjq/rzxPB82upOKtYsWmZmzZ6kizjdROK8wU8aYIcDoqeftpFpNgoAmo4i
85b66bZesvqWR7PZ7+75Oq1JQjNn0OrNAVtCUr9zGjGvZtOaixWpiihdinW5PawQ+E+pO1mEXF36
eiElYgrZNkKskNoWTcKwB5oXQLau1SlulSJA4nsCz22IR1yoLqpzLVzxl+CvbwsYPi9fXcX+dRQV
+Fi8sEogir09rOpIfOY5yk1HgfeljwKsqE86YZpJ2FEqfwGW49nRYJasNS3/4EfpxyfYq2jKxYNQ
cOgEizifGqXq50lBeL1/bPF8S/+eSvuSeSibFDUzamfIALyWIdv12OHL7sYYFfCVe3nzqEGcnnGq
ANA1viOZk/riRpWBEJg+jcfB7aPvOWPaQU+Eeah5cqg32sw2ZUP1/Ccupy76n1URvcKW0iZx5X6S
LouQ6yQv0xSbkYbJEE8UJ4r8h58ujtd0ce8eSzsJQRrpPFHQd+QtrFyaM2UsPOEVfsIxe1eRf372
2wIdV0DecSuOxBRQJ8fiw1tCqtxExZFDTVsd3lSSYCjxNE3AHxNRDT5xQJ4FFZwF7nltyVQk1xcd
Lf+sLPfu41smArEJPzg0Pm8PvPGQ6SfELA4EwwysdNNu7aPn0877qKIP5iYF3RxpK4upMf6UN06Z
AG2qgumFaMxwCOREb6dWVH8Q0zO+WNCkRPTgb8eQI7y4SFCChaWBDeo4zPrZFe2qoUBRC+jIWb1X
FqiD/dPvoLbJZUo9R/fmO2dJHeUq3ZIeAKGLf7jtUL4E4mZMkljHOanmH1Bz4TN7fCyYhWFCZnc8
z3ieIcgoJ+dJT5xee0BSXWGhxmuO8M2ninRxZKFSGpH1/Wbe5RxuWhlPALBB8//EeT4JLQ5CHMiq
oTrCsrHGSY22qiK4YUaQw+PcORn2pMzZOr7NV+AbEODRpb8y5Ctx64ZhB2Ni8IoWK6alqB/w38rk
dL82b1cHw7olSOyakrCRtaHowb699DFGIDW4T+NJhOL47wlGvPfxCPlq3/r2lQo5iuxV55C0IM6m
ruzXfVP24ISayMjNtQivyJiV3B/OiTN/QqdqJfESCvuFySukYdRguVSyyhjbZM/iAfrbrCmYAXb+
LxJCT9F3sLLE7Wi7/sA5mh33ownEzMgzBkNH82S7aRzuJ3zwXO8IBkQIYE5D8nihFFAdPmOvCv/n
XwHX/KDPsPtfhY45FMqLQK4DPODvY1ru6FQviISSfqWP7vCNEDMEuzzLingstqMhapuXHCCbPxnq
fIM5dznNtco7P3uOoeUshvO4/Gn6hHkPv3pm/ekzHcuP29RAInJdkJqyQScYmtQOniAfVg7qQ1lg
cMYu6x+MJlxrDVIjNm6ZukL74Zv4m924nteY2E63pIQLLJWRl7LI5ucrxgWUeatqYOQRAgyRB9JP
j8afJdXcLXcqsblmjlzF87lmGnThvvBIlPqxqJlmcUQRhOV4ckOhZAgfMV8/UffAP2PZEmtJhOol
FBNezcQ8zWoFh8tN/ZL42e67YG/zWTeiBA1jlyWJT5hAp2r4/fmHU19Ntazwv34virdQ8VccsaAi
SnxzPNPpfwGsplFtcpi/S2LoENsN4GzlJqr85KdTKf+Fg1UeW7QsYhRKtqCq4amOEmH+vV6E1rM0
YehD/EBRTH3tpYio4jP2L+L20i9PLGy7PnyXOMecCV9CaK+4hEyq8136gAgqAgoIPxYeJBYiDwBz
kbIUbOUjJ9Cz27kOe8/hsSsIeoMOoQP9m7vnFj2ytDcHLPBZmBCz+MORkE4tuZ6t6rSUHwzY/DT+
y6vCtSz0ItgUCLv6jevq/OQAPDdmwyX3ynMFhSyySvVZT2Tr3WX7YQm65MhZJzXeMSSLlfBkb9h8
Lldl2bSCl9z6mC+ScUpVkkJQRbb5IOJ86D0YGXIeoabgSpoOQxhrYv25yZMSRs6BaKfNzIo2Ma1w
Ovp/+Yi7d5JO7GITUa0HkfUdcuWy9gnlOPLbkfeT2ItVK7Q36BHSiRPAZWwMkzDtJaQlG4Ym8KGG
aIRSnprQ+ZEVoPUovQ4hvi7ZWR1dsPEX8QLH+aZxl3ZODsy/o/EZtgJy88lyaMGsLxkegN/0JpR1
LuIGTiFDjbNyVpv3ZkWvUMj6YKkP6k/r0RF8SgbsJccil6NO0Brxc6Y9xWySp2FaLzalBMP/E7YI
AmQqyCxU4AjSiB6w8irv/AT9MsVJ4hIddFzaRgswCCyvk0kHaKTUd+ebDXdeV434lcDU/w6G19Yf
nXWe84I0+qG96GoQrjsaAkd7GnNnR63tzfMN4iZ5TW7Yo4yr7X0R2x/yksGGSFZnKtxE19R0EWD6
A1qLVwlDqrkywopECkjBW0RK83yvhdH8UPvfsJKEiUqRJVGjLvPyeScjPb562AM5JOMqHZI68sMe
NS7mxuDhDQpmL0QVMoYSZFjJlGytPLJ3zR1EkrI71jPine7ThV6u833aElPJLez82BN3WRkOq4wc
+0K3V2ahofEfnOCv0NFullgUIekcZVuL5mafoZRGMJpbMh3fEcfM6eCM+jkQFFN0YwbJARlNiuKO
YZiMPgOL1XlXb23UWDQJ6ckCY4m+Jh2xMPKBvGB0pk5sKLPuHQ2mimZUvTVldHQQMDHN3cvmRDAi
XFVlxdpFhPVlY4RWuaKUhLgzWbZ9wDXLfVgqhpu+lJcKMo/s6+PPcK02bO88sVq21Io/M93IblTm
0PTdY31e5/2r87eyqTo7/GPPBsXoO7nGBPw/xLfzF59DiPYP31MXdQ8WwSzz1PEhoVqTHX4TV/z7
eIown1vSPfnel97Yme+LxyQjrHzkEPgygUdKy1dq6xU4MORdpG2oUHjQlOE+wpTa9QQFi3o391Iq
whyg1v/zT7qaGBCE1HzeIdcgSWD38auW6lUGziS3NDgBWCUNYraF2CyYrloHHunnl0vUKHMHzI5q
QJaxNSyUtKmxigZi8m6tyB8uzbETjXa4q3/FKXINl86RjCJPmycm1UmApgxUappp3G4+tZxYg7wK
GAhSz3W49haTZChwgAp5fjx0gjoBOjZsmSBSOyt1r7+4EnmQ9KcOIevgaE6jFnAmLrqDbXm8qRUt
/t62Tu7sM1miSi511tIxT7XmfX0tTmAEzwcB27juNFH8M6ws3YqXpwTuFOXo6ltwfot5HOgmzg4F
b/0SWImHywo09ia76dzCQMHLeYx5H8riFO2XorEMBgtI1V+9y6hjwYHhOz400Z1Fa6IIFd7mkXny
TcSHW+oh5x9t0iPtYk9lNdlNRTwi0OjjxY35yAewbJEOYWpybYICSbYj7cYh10qXTahPYsBkmk1k
wfXxy2X74rlLmu4Clptkm6C+07KVrTc54k46cl1fk3061LlWbq3Ai1PbW/2jzdPN1YK/OQrGMjP+
rHegVj2FYMeM2AxzMka7w5ePx7qZMMGegFu8ZvqALEhZLryZh9Cyi+RWLMrsW1BOMbXDJfVqN07D
8XQCiDkXmNhoedCe1tBL80XR110XLwc+PJeQqX70i/8v68Weo5r/kkDKfI6DeU2n9Mp7jQwuF1hO
c/qmEc58yI0K1BJuaIB1DcubYxloXb2aYFQtbLH30n60UYhSYSAWKQYZq5gLzVFbFq3Vavg2Ubgw
s+7n+lx+o4OI6uZSEpKAvqmqYq53NOufqK/lriDjyMjmO+N8SFzzfdRvF0gfvC4DuJh9HUDhBuY6
9GjZkQ+8YTV32d0DVbggd45xmUDWFPR4GSjyutM5+TxOkJxPK8elWj/lF5l8WPZ24BRu1NU0hN16
ktSIZx5N2NB4t3GShPUV7eSM/3SHkkoI/iU7zAXwCxCK7o+48S4JLnDnad5E8DEjuYuQY/1oCxis
mqKBGA32noXLrotu8F1YVgQvwkhtXVhPfZxCXYUPu3exwbBmzc5X7/rOKsVM7HK2YFpwqT0Z/CFR
wDS0y7v+0aDxs1DiptmDBOd+j94vQ9l1v0ePSnaUVi+0Hd5NZ3FtNUWEHIQ85ISz+vx7AZ8exobW
H+L7sEdxlwkCc2TPp11MxCfxoUgdXx4KJGUQv5n4ZGLzlfoZQVRf38+QCtnf7PsXvNig60nRpdYh
xkMQ3oqvSbHpyw4OTBv4H8I3Q2W9ZFXz5Bl4j06Rx9xgUXFtzNtqJiy6ImJbY4eYUoU5pNUonwnt
ENS/o7+1ZpbU7t9cLn2t5ID4Y8wK1JtUM8WeGvcfGZVkEq3nyGtGiqkyhZBmJ6plLb0VRWj187h4
JRf+QKWb9kWV9AWcNIUq6D5pyRMyHysr62tUsvp5TECQGiJzFeWhCdYQ4025i/lsWAu6ude9Akgh
CqdDNwaLlAE/+qTi69biTNA40qHR4MFsg3MsWQHssTK/OrlEoXEPn0PxvoXugJSDHu2rcfYKu9BB
nJv4cW4smwmMBWHs/0ESEmOFI6xYTPE0fuwGRa7PrmgU2LS2Uc+jGSMkctensRxHXjxyheuqn3rF
c2hQSZLmcFotXGq6MKvzzr/F7M58aXjT4MpezZQnFvQHKxlYs9UAWBWHQvlNZq8cLZgNbwFBtQiy
HrQlsJYk2mTd76v4mfn2ELL4x61lF8YcM3tPEMCveQFmb27GAwhHYZzf55n0sRhXOmD2B7Vb1Ov7
qnEsHSo2NL3YRUKFtpuyYXMQnyQ70Eqw028TCkeWjJ/Gjb839QXQW0CiIs2LS999e4A7IXi1xV2v
6jmLk6nqZeAt2g0+sOa1Ldf0/FAUIa90/R2KhIzZIkN1hE0DCmdyUK7fre6hP8DSxijVp2TGyzVh
kv1qVlLkbiph7sIwdnlZPhbqnEp1evH4bdMt0smXy2BXetBvPIzo1I1hLnRagNP8W3T8FHkCSV09
TBNM7FzzwBtMZKI7rmhimC/zczKWSZxhtLkVDjWQKZaq9teO2dGDClD8YkyGDf40J2mLSwUQR4bk
URTf6NIQulHjADkcGGVZi+wLrz92KVfYNE8LTL44H0InMyJjQseOsgWPfkWswsu9soTLTUGZSU+f
kwq4DThlCa0c2aVR/OP3KplFdDjMrjE7U7WOD/hPJd39L8hi4ngXNOYJNaeQwFK7h2wMh5ehkpWd
Z0GBP60OpnVUxR/vSMd/58RrDw4lZQ+edn4OqX74YaGGwqEK3PhWQthqnDiwhprrFAyWl2D0tnWR
SYpa71Ts8jU5pk1ZSs7PAGcQVZJl1vWqBGE50xGxkOPGEqCaVumMWQrsO0GD08334uQBYkJtQJ5z
bDROtN6m1OConB4TgO6ALYrGQGAQZU0Cw7Z/hH1Tb5aFq5rG0uD5eshUQF6eixA/lA+GEEfkoe0o
D35qlSaIWzTiK1+qYaNe4G4VF4hARLU47jTu5nw7+od60CuGHBBVrgUhpUe+/Oyg/9iAwrbkmzka
QeMy9DgEdtOjYKVoV8n+8lcSTxPIaiXmB6EmC5zrALbrOoUzRb0DcYXHpZdvpmSOoJxUDg5KXW6D
kTg7w81npf0YAnDIxLelNKkbApmIBnSMdF8Qv/LHFw4znBpdVpr4D9I46XSpF359DpebDQKSfT0O
aFEGRHHfi6NxbwYFO1PYop7jYyBg2jiPRb4A+0gFJY3D1mabPxnEmOso5lumHFuFRSoirjWwRija
ql5YcmNe4vDNYDorVNvi+Wwey9cXSpCHAmytPYO6n+IhTanPlC/IGo57Sr4grGmT5lGsIZDXjkom
D/QZLO01Z1zEMbgrViB5EQiV6jUFSSUOxkBue0WTu0XJf/3w302rQ8eYe6/1qVSwcQ/TsRXxPhcZ
25Ub7QJA6KthJwu+ur0441rSdXkPA5Qp/S34PpJCSpHy3A7+gDoRFKpoT1THfcDciye14KyenWiF
qwbYUCbkLDlPVM8l/AgNbYEWgCLjQBEad22wsaSL+EpRDihf/rgpamaqEFJmlPK65Hj/gEwfAfsv
XbYtoCr4ar+nDcls5GPfnp8eGG69l2VEUqTmK/kcSj3q4ThY0bdtiJG1xg/gCcQkB39CBHoGfEnv
W9NM/LnVy5kNFo+mRky0RsSlDYnE0W6YVqmC3cltG6JMgBrlP9zNjJE8Kn9QMY49UpbCuJvm5hv5
wpPNWG3EysCICsqLum2DCNzqgqNmQ9Qr++UnTHpNyP0/t+ibgYNMAJ4C4LdZzgvS+RkkwhOrWalH
hSJK8nmj2kJF7+IupXDJEbpfIQMWdNItC+iWsrELP9VBuOfy8sasmToPOsbOe+4FLtOiOwBGFFOz
7LTViFSZNXsSQFKYdR1xo7en/IPT6wZL6KkPEGhs9DPmVBAEI/tvSY9l7qYHkgsJhVVnpQvJHrjs
3nm9goGWl5usb1bsM/Kfoa92LRctnGV+sN7z/qp4ZCDW7luj+8ndhW0K8CekW9Yl4STOuXC8MyLo
P1ycHcX6/IOSE9CuqyMKsdkXd6dXHuiZE+4jGjtZXPUXuFRKs7MXOgyD4q/Aj1c4roadigwWp5t0
hhbEmWgFEUdaJnWP7kxgsy88iN8sgRDty6KmMsdGdSSS5PRw7YizpIydVw1t9jwWgZAOeGTnuKXv
EfCdKFke4D9is+PlzAj85wwUIdfJsGG+4SFdwnEwzGOA+H9lRRLemlMWAAqZ1vLWjiTfWfBRN3T6
dng5Q67aLfF6VNJssCYNe7t2SL2OFMlbm1DKnSG9BGFKOIHEQ6LFLt7IY9OluJDfqJaE7y1rZSP6
puUDolvR1yDFnsJR8VcwALFLHUMf7cKFQVy5w3F8IuGVKin3iNxk7mgdFysOiZYuBEv9GcCtCtdd
anFfzS/VHM9qHbtAzWPmAvsDYugB4kU0hqOAMtiup9Q8xpY89qD1gQN1MiBNq/YtspGT80nVeA5n
04xbA5VtgPcXjBzau7zFkriX22uIZmgXuVMCAxcAnFwGU1hvbiELnnG3b78/pJJq/+s9+FnBHv1u
lSeBjBJYt6eCgYaSOV5V+bqzb7E0txc2Z0o0B55U7BMhMwPNEK0T/bk2xbL8WH4jr/2/i9DBVaUW
qTjXwLWyqOcnljbHdtx/0Ozsziv5OCpq95d9BMZF8cisMCf/vSaO+XVPcxxxxoKjndqFZEeEnAk5
hC5qMijNvEG/PLnwKYNIGRlxijUHA/6UdYx14ClY/GF/SqWaATfPkDrt4UnrCC+1fLTIUlzY5s3/
qcRLdkhoJTj04JgtZIW8YZysx2JAzFjv4zqkiTQt3X2YPNnuK0DQ0LGGyC4jl4VPKM9mnYLIKKZb
CxhmJqEFc98kyQ4VjrZ7b9jf11ERXLTaVvacAut2TPu4I0a34AhaMuwZigb2WDbr9ieNVuH0vDR7
ktkCGTw1kzlYgkNrxpb5niJ8BlmiIQeT++wFLIKiesluY/8QotwqcSlM5Yoa9fvKUDxC6dxelmkp
b/9zBp4L73Gj0npzlsJc5b7WpAGzSoXBHkNpnkiYJbykdFAyYhIEBTSaMrt2uJWyCSaKhMHLDd79
uPHxb1LjBdfJv12iXcKrSUT+r0c7eO0VTkJ5nd/V9mSxgQeMf10vzJrTgd1MdvMqbn6zS3wzXwsr
jrkPumZnn8MvovbKnG7mI2NMeYxUNX9zlRNzhgdxhmqTMGBdW1Lpspp20/KSjKjXnNJbej0rolki
oSWgfrYxMWaNWb8Q1qC2OOEOThvcba4lokwx87C6LfPeG+nA+HoMdj62Q/FVOZF83XAPOSNMY9D+
f2wEUo7TgWIJf4K4tJJxAn6jt+p7j11xFrpfdGuxc96ldpbrZBCmxAzNOPv6EjuMW+I4IEJKKETc
pf+OLGRJEoHj9yKJetv7pna/LURX3EMdAqcpgrPomjuEAJtgvTs3qXuIyV8NS04IyoaRkNfm8QQT
UKGIMq0rjrhRLV3X2/1j79Ue0K8P/pz2nzHsjYlJeKSXfYI+G2uxJSFC52PA870+iNAoqX6wJyJ5
DKcoJQmEdh0oDr+qC9JQw9HYLvO0WNcOz81lolSx8OakNUHg8+YOvbTmK5jIcX9LEf/OPYUxDKio
uhcGQWB1Ci+XdwQcUof51jAcK/xjVC2wZgx0oUwHPw2PDuBrNtN8ZLVe/6uIIX3XApt4CfYBHFdr
2eBZJsVEySUGrLYz8hoE4OzKR+tCQhHrartH4KwDt+ZS9o655eAybaV620IUfr4yp7fjgGp8Zqom
HS37fs9IChB8bAza5PmFOCYAfnZPS18Ga0zZvg2C8aNIPuv5+akYdX4xdnWaQxmUSb/mZufVoHxb
PuT0zQdQswX/vJv9CP2K+GFrjF5I93H0KEkLoQM2+neWQIbXc4VOd4LuhKiT0WJnWjvNuTkVfbuT
buEV2HvVfoQUWCvbZY/EIFKf2rU78RC+1d6z9BZE1P7WGyfhob9XObbUGbpjxdSZhuuy3G7HkdjO
uuW6ABViLtmJCHJieBTI4kxW0m4z0vg4+bBQ3/Ht6ul9coGLGVjWH9iSDxt0tLpnylYEOtKCjrAv
l8My/A+nu5i9CXanTZyKppZswWqyBxvUyfEgm2r+2bWYwFINYWXMhhYpyf/LmywAk4Q8NFHvdGYo
B0PYsW6RpAaon5j7BNfGVlLqqQo5ik6/ucUpaWAb9UlG+ii01alki4jl20/xnicq3Goe0YAsBbFc
wAweZwd6gQlpahjKGiLBa5SNxLeM6eHy25mY7BlHElVndDgWwV33Sk4i680Gsz/tTwx6H29cfg8A
msW/n2CvliIAVCfZr0q8dK3ldhPG8BPuHD3VaKI/ets/AWxbF7F2QZWbPV9taiWsO0DFchv/5WwY
1T65gRF5HyG1VEBUGoH4MMvguxQRkPHI6Ef/1f3gdYsiHJjuJyljYF4sRCwet2wkMD05Z8Ehhq6Y
TVbiQL9CfMlBzS78La4VagvvqONdanclFirzcztWhpaL550L8K+SFqvO/I3KT/nSGHB4PowJbtiY
HahYzXQa+YRNHQHhvJczVMytYKu6I8oJteIRr3tCTon2dX9Xns3aQHx8/+6Mp5G0uqPdaEG+MOlk
OKhFQ9lw15O3UBdrWlc2pn2ocrso3umB2HfgwHxhkOVoKDczH7s2iw3SB+lspanFh98wA0UMV3Jt
/LS8IyaV+9jN0KXiCaY8OZCMejCzKLDIAnZiTLh6LK2fiUA2VpbKvBCrUuP7CdUFeZ4jKQQPk6I+
PIi6LQNjOe+yDn04OpWXDW94Nq2/VmB0xhBg3bB1JmgOO/kyhGisVzbaT48QMgm49A9uGaNMTRYc
0fCTpIV8L/696ulBDU6WHE+WQqy3VO8XhEgGl5wKIdLr5EJt8hzZhnUkc3lyKSFJM+LqjBoMc6UY
ut8JLoM8qyMf5tdI6u7IHyaSkYgCBg4m8CmP7R/WrHjt6GWr8AoaCJgBtFzM6l3FZnop3qIZ7JEx
yPweOdv0YeyrH0dfqBA03n43HtuOWdpn4eGrCOfYJgdkLqFjWqaslov6E+8+xZG0C4NMMDLOFL2e
JisG19bD/ZijyecL6KMoedtYXCMQR7ppnHd7CPu4/53Ov2z9OYqB6ajeNRxMnRWMxYCaIIulxNYV
jcmKSoG7ZdiIc3qgmYXNaZAAHDyn5dZAAaDrUjK2UPwSCys7aU3R2r7CujGYdSeiYDhaYA8sKgbC
WDrnPOr93wfP00ExIq8hFJZULD8nlNqCCVIAHEP6BkvwBWQdXf61qz+5LZBjaW28bbtA0bpzD8Hm
xqUTeemM14ONYscEE/eqlo2ZZfUf/8dqfxsIzGIELYNXLHgxhEFAQ1a3xxbdZGQ6rCDK06ab1IiP
kNrMSsR0fQ0C+92d+kR/bjZSKc+Uh1tLWZcnBntvF2NOLgl+CfvLEV2IE7T5ttzZeuWCOuFLpLzy
U/QGERc79MC5SLgzjOXqakH2yhzeF30o8asKvJD5vKSmLqgcT8pTu3qIq6f4U1JTAv7mhlPzbODc
yL7JqBFVd0mP8/QYIYUZESAU9kPzysJY+5l0Fomtlpuw0yeHsZjU0cmxlqWItFWtkuSd/Kep7Am3
iVwo78GBq8DbKp/U6GL6LbzQl4zeMkGxaKn8wGrSL3fLkn1xS6ZyYoou6dn/9ZHIxMckbS5A5Kim
TYYnYeaclmLz8VSzmJgY+QRFE1rR93uNbI/4g82XCCDjApLn0LXMFwUpXryZo4lF0ZbIUBxBNyYP
0MhaZKYnUWzf58/N3aKoGdolNlOLAXSdRlEhuJa4CG9hVR+urBQ0jml6l+Gwz4c5Jl2A96niJT1G
TwUu11Lv0bEVosRurOALmDmk0H/aNBFxS2PxKS93a9GyoFYbpv5FZojOIOSoPdqj7Bm9yS2FgPqK
8MhRJpg+Jhz/ddJOaHfB/Z9In8Ic0QkApSx/vV+NiryqEEYQKSpfqJih1dxJW6sHypVkZnh/xYcU
CT/rZUIRWhl+In3Gms5CFdqTxl8Pl0pZefQrqHi6QcO3CzYfQPtfkoL5zhZa/luZ5GMOp1wHTU50
jWcXSrrbs/fm30MMF53eoX5Ko/kMWGUxgSvqMG7bxRQSMHA6duy6XjjfNefLQBeI/LgGedseJFfK
d4gZ4GQmBGYZrdqPetMlRfC0ZoUFxHPh+2xdbqaJtiqYohJT5GLND9l2li3XVZfJvjn81u95yjWk
gppS74CLxUYk79eXFJjsrLmkWqMiZK4ASmk1k6GplFyySIJYxp1B/jtPi96w1RHqBejHRuS+pK4i
R/aF2h5DjjIMkmy3ie2fVNrJYH9+CXtP3Io1tOJQfq1us4tWoW51SodZgBqixgG8dc855/SCob9D
P92ElLmGAVe9vD78tfOIr19NQGsunPxmzcbIBDE7K0ff15pUWmd4c9WNEBQRwkgvrfYAGv+UfixB
huqN4frE3aK9UsCz4BXf3ri+7cAoE3CC4KMoaviPeJ6N1Kmz3VxoBug/8ylAgN+eQnXwg4nqjWmN
J/PG8UFQ9e9eMU2dN6mMzgnMu2zL1MbV/JqBLo4LX70Mb4R70FQkLzsLvgzhcKk18sBKTq0ZpzJW
f02il3Jq9eCZaisCJg6bnD+/GHFOqCT0xnou46zcJiYVNLWAh4Y2dOKfcFaeVt9hEkJMDq8XRmOh
1LAFUxdg7TkOkMEc8DRbdyXQH7dunpa2v3jylACCN3OTcol+Ngia1JmP5ulSdV5KA86/mjXeUtLJ
0JScU+JlfE1WVaBB5fxpFbSuvL6qR4dIEeNEEhnIQI55YCJSmujmAu98Q07ILA5QRfQGypzXwmO7
Fn1St1jI0AFm5B/qM7D22HYS4BxYyNIFawZAKyQpMjJui8FgcvhYMpH3zeebflx8mqDwcyFgIbd0
uI+2zpINve4T3MX9XoDAMMH1YcHKKODy0SJJ6FPY8PekkmgBzURRGQAg1+5wmQhwnSHfX9Or7HyU
yg2uE1refDSsr19HO7+veR4XWC06uqEr/HG7fdu+ZCnFjIC+hOzLbVo87ZlcUqqgtaC77Ju3x1dH
3byXmyqfYuquM1pYfClr9LEBuYvPg4mieWS+9T84kxLSIEXEozh+ZsLZqLFIeU+5yGhrDNwz5ttC
Y4YKA8ga8iEH0kTSsAe338X6PAOwpRyv5VVljfqP536+nJScXTUrtx8neaIllSCRi32CChIObLe4
ho5CIbQct49ITSPuAGElDPsRbNHLzGHK8Nckt4RPQuiECHLZ2RL/ZDd34ItZ4Qa+5hjYA5FeH4QB
5kkkZCn0ZQ5JLsNzUtCLgE/ccyjfdJ7bUOrPFz5Wx2pR3OLAaXOmKYdrIBV2Ujqg/594wek2MSZQ
gSvuPL/LosHqaPI8JHVTBE/+Vlij9Rt91NaiVW8hRFD4A29Q7l/oHDk8OSZVR6fhzAqaUHIhi/8n
O+PpUdtF+xKh2otoejJ4clnLmDyKUGKZjhJC4/1Urmp6ld1tvxcfn9RI/g4Jsv6IT2kAokMuld4C
F78qiBS87waKRo+FLGhrqynjqO6segDjwGf1KAbIaZP1t+ck7Z23JlfHjLgFXCwacKEUNmA3bwcO
zEYjmXmQszeoJbF1hFZA9zwNJv284QGZdOpUi7tnh4ae5QUv8SgeSALRYE3IwV5Ti515YiSsLjbH
t8d3G+wtd1x1k58lz7b7/XmIP34kdGBZn56fMkX7lo35Lm0ShJhr5ScxDcpYckDAj1X6fYh04jmO
l8YcuWwKrBKkPRbMAseZrvF2puT7RA1DwdwIF4PlWqWGZZeVRV9zulkccCMj+aNTKG1U36JfWCKC
/796sM07aSGteLj1pUH3jOsLaWOUp1VzVHqRomL+e6QbUEycjAGvDTxOVVMTlDyEnP2W+prZHaKT
fgCBZgegOBSCOOYQq/soOeDXj0gpcjs+hRiHfxbDwgyTiqZ+Eo+zcMqzyzie0Qo8H/TGdma/6YvX
CnpLpSnkjdAAgtEdMn+/e5+OSNCyfP4gza1/S23vANUMgSBlhaHKQE5G8p8vduBBQ5YK5AUvYfqh
9TjenlVCE4c8ysiHFZDAyvHzjObxOK7vemGq1Rgio/dxD0kCpKBfsiAI7ted8CRStMe7N90Lte/6
iyLp6Ew9O+lgfBU16iJPmqVBS4Iy6XyVn3B/T0MuGkN1EK+KH4AS7ZVBj9Mlh0b7KdMNp2SWA0No
bRvBkjUlErq9KlOTjnJgbqR6IujTDwoXz/k7X/67OcJisVZLH+xj33OuBbRp87qTTbxtBD/BXpAX
oPR7MyMvOvdImA582R279IEbLDHw6otMbBQUzKRgj5y5JTebfi8RCfLsISwQjyi2MXzyGpxz/tRG
ZUriiYJPKJLM+t0nNl/eMfc76CR1sV6jT3WzJymW8QZL84GLcwF2uhKulNKf9Lb+I6zCYj915HAO
bG++N4fsRJDLHl1yq+vLGbwi9UmvINnsLhovEXCVVl0RJfn6Iu51p0TnA5mVdoAVw9kNDQlouFIQ
cT155LEiBhePIYhQObGonJw2tF774o3GZOO1Lxe01M5exi6Rasxacjljd2fUy3B8swMYrLq49isr
JsLPlm45XeudEr8a6P5SBf0a1Eh/gLK275Q5Ik97CZcP6sq7gRXgxZHLfHx48r9trCJfcT+WX/s5
OhlcNcrWlTJokxPK4WyANM9D+YtevKpkjEvrcR0+9DzintnTsRa3pmIP+9jC3GVDd5l8EmG21IAX
QzXpRQJhzHpUF2J6UFer24Jw+XcKeZpiwURROID9frhtRIayxog6Nfgvew5nu33pXV2+vmvk+3yQ
Y5QEwM2aLLhwBMwEYadpGVf70S2484QLC2HfZs0uOEI7+Z4bLv/yrSzg8wScHr4yGgEf0lOnQoo4
vGbjHGBG70b97Nayz6YTC+tISdCc4hl+Prf+RCranQ5Sa2UrmrmCZQdQS0U8IXBoHxjFSbtXv7EU
UeVgx5JxwObz8HtDrxJwaJVRX8vfisAJ9Ou6YKx0W/AU+0bhZnX3hoPFlFOocWO+oifyt2xaDrwb
WLLPu546wXtgCubdZQf4jcigJBnneP3an0eLYXAnuEdDRJdMIM2Arq+pQtkNmrozZK/e11v5w0V8
nRCJ0gF1/iUYPofWNv1SDHJbGM8jsEEJ/5jnk04Z9PDD/srOUiBS3jsCA4Qe5baLRnbFJHXgTdRv
Wf0s6+3iKe15P46moMdlypwShxTt0D7dKXtkfvBbLL19lJ1Wf1Oi1yOn4psj1OU86rLfKnVnHHcU
4DwxsRXf8FpSL7Wou73hts+6h13Fn5tJCzJMSBoVz7NT/qK5PU+haQPXSyRWKGRc26dGkwRbzl8u
vc9rgdSD49HCnWAWRaQyVd1Fbb0wNbb5sVTvd+SN4cqr4u0Yq23QKwZTIsEM788qWp5q/e/dVrEn
NyGdW0fbBDTlJZGCTMNZ5QXQjjvNofTAzgrgxWen1Vbj56+vHE96rOg8qH0TRYYserQDeC3F6rTe
Lm0F2OeGCH9yVCfavEb1AnvqKMCA3N59H5pTubnIleex22NB12XRajGDDvU4+cmWcLnijkokz0Fj
lRuH6rLutI7jePmh2sYIpD6EVQXzq5xlydd/mqh0wb4zSCNJ4cEqafIJLpkv6WG5FX8/lSaNXFxm
wvdYLDs+H8sVjb0QjqIs4hj/0LEErP4yU3bC3ly7tttbGH7LiCtxQixQC9xtBNaGs4c7lDRx/gJL
od9jjbXkJwfDTs/592yeZ1sqXFNG8J1OXPeuMyxN758QCPuBOqFmQxz8e4IkLCNFRvYux5P0efyB
4/nQXFB7xKOOTcVBrRy1XADcuTaqTWOOlNNEJxDpf2E0uNz9Z3bjrZumeobLNMbyzlB9i/23JN52
1+4ONq8zkIHyPtafRKPJY9iq6q5opvEhm+WL7avkMACSaMfA2N/NjOmSpsF6Ap+ZYLGAbZKgr0Dg
5qcj9mgmXI+AKy3FmTHOSW7a1iXZBJKTMZq7cE5PkEA6X2YJ+ktdRWNCXobgj7xhafbxnb/d/FkB
ZR49+lgSZ+/QNXqmtn58lKLba3ufPgKZk8G4UsJ61HVO4d32Ycv2sqIrK8X71HccCZ7l3XJ4QwFR
cB2HFRxDOXLP9odOSipvAgOwAyk9NwVxW3tqNtXW+hvgZhpEWeJe0L1H1kCxvTuDhzIrtquKLWTA
ateygehKJE82ZWqV7/T/2b0NzVNkyYKS1wDQF/g67SHmJ6NKIWua/RejtaVhNu6wC+4vgS7dEuJx
dbz4csDq9fAi2TPB8fTcWlruNo6N6dfp7DltXqf/YY0gT8nWHVMwRnMNsSR61f7UyHTtLhSkxo6T
gFJ2OXjG68IO0XJmuj9PjUSLfs+OkLUn1lQg2ER6uQj5OwVpmWoLRtNtY+0cS165oPy0/VlcptA6
o0VWVw7RlMN1DxWwGuqdzTzhiECNjb7idlDLuoZ03BRKaSMzOvzd6SLB2Ys6343ZwxcIqiPK3Ftq
z/Ltd1px4kj9v1F51oltvARByxX8UItejuBnqYgviIy5f4Dp5UoGh7X5cAaxPYitHfPNN5wiyCwq
M7a8m5KcjpEbsHw544rjidGXFFStYEIxf/e9t5F79w0mMKDv6nSAiCcRJAti7RZL4hzL4IaXaNia
6XBnKjfYcNddMwEsyKkMdDMoCi9CbetUO6nzNvA7Ty6sdN6UxBhH54geXIW36P8DHQBeYcEU+E5i
8k4Yzr4rPkKHlUdRbS8NAS/DMFVk8mbHnuenPbqXV4x8nnIEMiT1Re9CN7gOz6B+ZLPba84Xcmlh
WN8eHDx8pAZfP+b8gMIpUqaWBjoIF4GvGgcIQM8XFPEul8ZAFAnI+oxP3KGKsQcGWcctFoDGcRfS
095B2n6JftN6l2OzKiYWzUTWOpQ0iNT54yONkyBgywxYEmrTWoayhS5ursbcWMemkgbeBMXjsaji
Djia2Xj4+NMk/zgvNMTyl0RVc3AlWRmcL4KTL+5hsmqvyr+yQ9v4RdiMMG7cvue1ApfP5eAKhV4g
gUJ+WW+CrFTgXi3MyGL5ADGrdCpcPGYFsQxOUcnVvNSKOpF3/tSYC7J84xwevhaESi2lBA3Ed6eu
JiIYs9SQBzJhBRu6Vbpu/a3ZIGFOiRhdfc5Qpi1kTXpLnfBIXIrSU5UJU9oyTO658VywATbdzPqd
iVkT2tUvy0IpmRT63H7sNxNcs2QZJ1kV088HUf30xNAzZJfE9y9eQI/1tq4VmO3LslSz+9A6aZd+
Dr8xF/Peo8zaOoisY1njFTiNsN4If5bwZrg5d+NwXqjobpbzFuq4R5xwTwhy19F1YaUuYmW6w4Eg
lsIUhuafpU0Xe195ycg5Ne8oyZn99JeHvvbQAxIoOBkcKY+wtMjXOOd8dtc6pfmJJKguIahJ7b4H
G16yH55qr5p+SjZWcH/4tE2OAOmsjIZ4i8OJdZpl8oTo9RvnxakJdyIuoCex7LMXd/BQVr/wnrGz
1ypEB2mIK+T3p3chA1PzI3BMbbE3qbG97ocRC1HWMbHKu2Okf90sIol3ysDeUe2gd2r21XtAHNdk
0Ue2nc28UtLMOYgg8j8GPLzGk+yZg4+caiAoeh81T0LPa45Im6FrxCvHNSBeJrg+EP6jET5rFoU9
MxtR2HkloszxG3XdpEyLlHsseU/PfjusVAnd81GzYiF20B+U85SIem346/36nVJ596GWmRbC0KYk
ATF6U/YW1vg07aMTQtgJwY574oSBPNDb4NHcwzuno+GjGO4T3NllJKdSQMz9VXZ91xafh+Qcscio
ss+vUv2PTh4cTb/tx6yX8KFn7uU+WvNpKqEgLJm/qONsPt1fw2GCIbZasrV1Gw89ITARWmNjEiw6
C5nEvIKIsFgckpo46ur1uiMfpDXDqI79T30wc3jLhBarQ/DpWSWYnu60NSBfkvl8GFn1jx+vTD5B
AFW8g676A3B0q+o5wrx/MteWD29bSTxfSswEMGOwMrZbQ2WDrYdwejhtCFnmCioe4kvnRnnNxGd4
s4TkJ12Y7ncs8+xSeJG0pAMKLib0za/2B7TQojxV4FunpCWOHqp0ff2fRXX6ErjJwGchs1KRRU6W
ukL46y04EKaAlQ20+CGqBdXd5+7I0XqLZL/7+OVDdvj/5b2FXrUt/LvFDeexFIbr3OQlf/+GvhqA
2+TjSiBQlio4fBUItx1aQMI0DlpQu2YgVwpHS3DAO8bSzQJsv1sM9NFEU3W229MOJtqZCgDwyJNQ
JdhNoMaNmeVZhMmyhBNVWE7jok5eAczk5R/k1SLZDmiqomVy1wk3Gw/+z1WV6fRTnlepWQobiX2z
lO7wCf3bDPtpi5oFjCM6jWuJjIfDLElA54NoK1IfiDo4z/OmM7FgQzkU5U3MGhiqAXNDcQfnnJSZ
IkxAtpOA7N0N2AaY1GlFvSW7LOIkj3ooEr9CrP0eFLnK2oFJd/EXPf/31CdK9Yp2TmZGUyub61+3
fr8129nasiRPsB4yFmGvYuJelbUqLbiymnjaE/HwSUSyHr6cPthp9MhLwS94026EXX9u/UWE1T/o
wnsz6gHzsMzrVIPy5j+dm3c7dTSeJHE0Ofa746Qx6qO95DFi5CCvYXrdptu+AzhK1/iDurHUKLv+
OpylU9XHLP1Jk90feY0wmDPxNtAw/Rm+AjRV6yqR3wRfiWro/lM+539iFjyv5p/eMgbEOv22C/qg
Mkqf3tFHi1Kt61rG8fcXq8uQCRdR3UL/P/cywxKVA7jByGh+Yj9czvRCIKByGMyZ+nYS9xS5vXQd
hp7ImXQAhRNGwdtr3iMCV2QlPKLEq2OVvW/48oHFg6dwTadmylyqtJOnJDTOxZFQMLHIIF/BzIru
YTTuYSFdy9mzhoOH3lnrW2l5PS4yKGf/EQEHPVHxkcs10BJp3pVWumgqCVMFnsBOPTe7Q77xcD3/
ko544VMHTuRzODEhAvjegHaJjIooN3xtC7uAOMfPJ5i5jGr9FKqP5WziL0Q0egMR+CzeqmEojIPc
s69pt15OmHc4elmatjk/jM3lxNxphZAAIf8PzuR759D06jtlGrHngkD6BRusbqSE/jzpFWSkYim+
FRXV4CsRfFjM9iwU8sZasvI23xa/UF+P32eDVeZTDAMvIhUmbtG6rEVZvYcC0fjSBjqqab0O2K0E
ojAA+R8iGg3ntNu46NEq91P8/pKBW4AG0TLmfuz+PnhzcAzIkDUeyEiQX3OCkTokmQtEiwPpPS8l
qGSt1X/98ybX5v+5G7ge7L3Njo/TGFaC1oRTFwXgjFd2RDlprDfeCRO/+Gnv0gGe8l16KUh9yX4K
yUzbBGd17V2LfTtoSHGrYK8vhqgavVCVkRvEsADoO5lb0jn7YBmmSeJbNx2K5eH+CpsYEJBWyB8P
4ADmcHCPNkXuCiLUaweIHGNCggZMfRUbd7faxdzjb2329MqSVkckixKgJ32cnsjab4eCVAZnUuGb
nU0EzTbLOntEy1RIZYzzZ8MVBWvs2o0b5dF1OPTKoTpqm69bWmHoKIN76Gr9IX4BDsuBoLSNWqq1
BftiNBq9ch8s0Zvp5ygCqvVrvtls8AzT61tUacish2j0tB9SQwxSq6jW1QyjM9VZ64bQOO+bDpkj
trbbsX5EShqYVF1CZviJmBE00TwmldMp0a/ONEr7jD9ZvB1aFAnbjnQGRflmadGrV9+g1bL2xtWk
2IaD5KtaEIpEP/Z4bKhgm2MUB2jhPJtn2RPo32Ko+fGsvJoeWH4bBP0EdYf2oBS/nTv+NzCZ4iIj
o1V6Bo9C3Qkm0cYnpACWUMnbhuNut6B6hFzF4SQdjzOds6szFdmrfpt6GqUBmsPuTsQNua89Z6YN
+KabUBQzS2DzULhp3Qf4ojJl0t89EylWxdjfgLGe/x1AK0LxWTx+ww5aIxvB6REXHHtD1MaJGVVq
zQeHQAuyzUFBx4bcX2D16XocyYSeeYd1LNCr9bYb1i+WA3G30NZWxaLFbNWSdXezQxD5RyLecfNd
JpVhCZUOY1VqtZqNPoaK32UnCMpt2qE/J6CzkiLhRhyy+/ptaAyQQ+Y7xzQ4OFOIRjaSro7ZN9Tq
tLJMVmwUv0nGOQIgT5a+L7Bg5s+GvdVpkJvtIw31rGzVgNZg5oR6edHYWSFTUsdDKqY58r5XBDMn
LRVHv23g946BhCjxKIhQ/OrDVqkBPzi0BDPQZeQsIpgCwehteE7yy4UUahRuj9F0nuYq7UZyM5dS
6iamHpSae76nY9r47CnmxO/pL0VJ4Kh+L/A5hTsI3zt4cEQVjD+xNMDYLUA9gZaYrunPvtsMdIQG
hR3F/hLMuadFECShxCnO0UCdwqMlfxcWQV3itmjKCy0OKwM3N5ZTH8ey0GG5cvLKQjwUTjjQ5Yuz
SObItJd0YYQ12Y5ktjgV7lxVNXsuj7lTZRC4Pg6qw9l8w9tIM3Fu05ypP8alkyiB8H69vSosGDGq
56LpOmkTS2vpgFues+s9Qzl+t7LLbnHisTBVcz2vwuzWj0JmBexMjCmPSn/QuAe1bNrqSG6zMoeo
sYofVS0qKXcfO1Ii+WVcq88B/NSK7/F0TmejXNj7k6Q+parvYwVFrmXA183PjTln8GVWW1SQHbIJ
tYRHhT20Ky99cPLl3bCL+HYoLy6B2+jDN9DbO5l0yFBQz3ogyTFq8ZMV57hpThEz8oODqkxeG1J2
mYV3u4tgRsls0aE2p00dxumz+jM3+btl+Fgk7aMfEtv6coMDMwTRMEsTRF3SnmBZ+FvB7/vUw3Bl
jdpJ6vNwi3uDErApdf/zVFaVfMGtsL9oCJKbpmw5fHToH+2ZaXO08HN5WuDbsCJCEFZJe6UPb3dN
aqicgWSb7xiaV12K7X0GdeZwamxgKk9cp8LiqPESn3ZTrcXXiSF5M/B4TWnhbCetHssxH8uyQb1N
/+K+1xeHcEShteTquugYpD/sJicnNPSe/aY4qI1gAd3NGe762j2+T6jcrewF5xEEJhj7wY0WW8o0
PtjqU3cg1HUeJE2b10riLCJ7o55wNQ1SJnFLagNCtLg/CZ//ElsuvduKkjmfOfDKO8KvxHi2hHdl
cG5My2+3puKP959dPXCz/euHGhUBAyFnRsoq+UkY2o6WC2houcVCp+59hq4YxGcXlvbbrXn5wA35
d3GyEhUiBwQKp9jsH8LHoK1PNEmj1nEdBy6FLp4KYV8yYh7VjIZLyqdhLx6kzcs2zW6prB8boW2q
VkxvsvXBpUhes2rPesAIPaasL57u4B9yqLoMBqSdPsEJdklcX37Zt/PWPoaI3Cbyti/hWmJrNz9C
sL2YZ2xpIGO5+ST0U3c18eY3H1hrg3IMF7NuaTjxmQzVsep15dZGLR5LVsxDW+Wd5aT9deXCRlXD
f4YVh1oMW82Yyh8eqBug4B13KUwBa3SdYhExEQRUYQi6QfFc9svhAA+8aUv06J/UzWG1OjO+TZ4K
RdospNG0rwDlVm/j6PuCcvHJT/jO17FVdmrB7G5+H9QM3sqodYoo9clVR0k5axslNkCBE+PUFgMo
UHlkATrf4khkAjdePE5s8MybUP+yNP7siXua47t3KCm/Wj8wbbMpfwIjq+7sOswL/fJKMkD60sLl
0A1GatoZSI/5A1rwmyYHkC+KGwE/M+dlNH7OBebk4z11R2UM5KgxndMPD5/cZU2+kfkt3Z5rtK1r
XaqfZM0I1UdcY6wz+trJIOGN6ZMor4Z0kjNIIncJaPVA0ejDXRThk1JxPc3HGK8PA1s+7LE2MLdn
2tczevT1xMPumY28LtLsgV/vb7cr2n+9kvXWUOAo+Q/IS7LK/uKD8Kg1KbjH7YyF1J34dte4Hpao
rGTxBDngHUbZxbF3HW4u0rGYQVv7uWALx0Bvc7D39aaMx85fbPOk5pI+Lg+B5uvSPMD145QGfHMQ
YR5PtUE93tt8akNS6I6PUnw4ps40scljHHTwRbNFATldgHhK0gQsIx8r10oM8g5HD8MXxTOh7qey
JoELc3dwABkjlkjXoHddgvVJfkXbGS0rWENL4VKIZeTUCMYjTDTDHwJ84K1hFNGVKHlId4aOuKrB
shTRXIYx4nQb6SdVIOiPXoQDBjcFzSqAehOV7uagIkkAjew3nUmz2Z5CbRSe/n1rIP3dZrUjxmGA
tndbM6YqZFTCuJvoHLqLcZQFYNic/mGzl8/+riTXApX/5EQl5LtjdyVSJRSVa/v86+CAMn11678I
qXyM3FbdOw9rGElDKJRh8XR/6aFhp8rHgGCyOAYbHRqan6PkJJFeLhZydbjqICJ5Ge+xoLnLMW7g
DCiSdv54ZiBy6P9Nq214fRNJF4YH4fr7/5iMR2M0ljrng8RJcfCNyFHcjaodXLiO7eeNrHlsxadz
h7MzeaXMgLgMG4m+4CRhMW2nn0kpu8b5tL3B5brUaN4f+cfNopOosWbXDX7EvR3xjZEbUFp6CL3f
5VH+PEtWklzi0cdGEzDzGUh9wv92cIc1lf8fA9GLkTjsfN+DHFE1jyal+V925ZIAACO1zf1Iqneo
VsOWukuH+494yooVnn5K1JApXIpHtr1MHDDIGsDhJyvhdrxjHZnGdIcjj/GoR2DGlwIJu5TglPv3
PBh7mhdaYEDWJirYSLGKI030L3W1q25siI2OA7LwqJ59ZbyVxfQF7n77JZkw73+jTYooqlGnIuXG
81efDhLyW8Jf2rJiv7ZNqrx4U7U66QVgUUI7+r9+U55etFyn4PD807+s10WCfefvJyqBCn+5sYYz
HNO6yF61v7BhJMI5PX+eNGBvZWT60LNxqCgmEZT4JsD5skisRy672rMcvFILHgVlMQg7lIgWe0lj
1cxbCu6nYr5MXCQdGq+Rs0I6+d8i0fJdqsGJOBzyey4AdBdpY7h0BdoNd4FAVSLmO/vlLBWPVxCe
EMqEchoqmafboMht1Y8RaHZt2codsKxf7AsWJmHGzec3bwbwf5WqS4hW5M9L3lFn+07oakTqzySY
zbfhVL876y6P1mRMACHpIg+Gzq5u70W8/ST16Ixcevclxsl+DBl5aluLXHHu1KFVjiF1yofNZYTW
GlO+fRtD2KiVlq3zE6QFqIPwg1TbmjsoOc7iUrK0p5d3Tb1TvgsF/tAyy0pwc3xqDDvH9BzIyJLG
drFJnrXIeqoaDB4r42/QUJjX83OJuVm8kkSmZ/mSMPpjMdog7+fIkoz08T6PqQFBlHWoUWvvQ0N4
gsvlIVXkPcSeSasqQ7VKQTFTPgWITg6egO+LE0cs8X+Dr+4I0XrebeC3EuvsmjNpao4lhQYNno3j
ICP65itM03kC58Kx+OnXlky1wmzGYmO1NiNGBDZzrdsjtVEw813a1Ran4esEcBW6IwaGCpJ+7URc
/apKmt3kQZjC6lEqPaihbtzYBCD5rhlRAlqMBHFFxjSIC9vsTXWpHbmisRjfRrpemKWRh7YQkeOq
q4fD/9giZ9ghUAusWD265RIZxFuhJe26Q/wL46fj53SNtAl1uuTYCrv81oNheHkBRGT8FOLawZno
U1EUZqNnoJGa0EUac2mkfbdoybZD9dlm3cjrktfetgLz8Q/iqchAk/M4ki/0aQVWySJQMuXW+mca
AylJo4NU+ZW5sJx30SvvFAV1WdW2//+DyjXR76wfbuYL7qFfF53dun2pixK0UB3OjcMmQhj0J17r
WOMDdAk+l2m7yFdz2499Z+jjuflCEI3YNoYX6aO6PX/Wnpp6COZAxn1W8O1tN1ViXrU3aFH+Thb+
4/FFA5sVlDplJkvS5savfXd4nUbDIRPrf+NLmJK9WmMPMF0N5cg1t9F8eDUcS3V9ZEZCx10bO1YV
0Lr01lMYCNBkpk2S8MY7e32IG2nqMwkl5t208/GtKnIX/MfnfC2PSdDZbHHmM5sGfx6N0f16esVA
2Dun8p/k7904UHUfp2Z8h/7dqdbtDj4d7VhXz8H0cPUsj9ewupJS4lYAcYCgjlHUC25K9rRbwT8k
p9A1GkogjFt3Sk65Hm+zvuNZdz8VeBD8rJtMlJF2/W/a6fspWCPrApEQmKvOlg/OCE9FlkMgcde8
/wGNxuAwmg2wJmpyZLV/aiBBvfltPZPpB7bLimpfh9tqEbCLQlWDEbGx0b7HIAQ9cjfcrkASVTXF
E16VerU5SknxIHa5w+OJkBQr1sz4E1mbPBh//LoyuAWtf1FJbFEgWxA0uR8mWA3pSAXWesPJf5J5
wpgGhYeQ52v9tuiPAzNrFqF5V5eS9fJIlonGyVOTC2T2J+dJ/e0y+JeJXL3bhqgxg3dX0AMqCRrB
TUHTNoDgPV1sYZiYSEB0vSyAbTxb1dgB+F5RvJERBvY1qDQADBBnXKjEcFnexsJWhgiwu1r8RQNj
S0ELETph7fTX8IaFAHCdtFug+9Znzxe6P8shuwyzE43WhIH8VzgI8IWY7HvuQHq+ngnKNkyPiOch
6zASwARZCuU521wzkcF9IYybecc70IOvcTO3jixY/fq9JDbgGH61I5j5nIJxutJIo2CofUj0hD3W
N+A/FDnMhpWdx74yGU26t2HnFFjsNraMojRAM24+b9KricAFW/IxiypG02IIPQlrqIfEmvoP22qk
GaFcjhMvZ7BJjpDPpGv926U3Cy6l3K/sk1NQkXE7GsDK7BO/oC0d21qEnW2oi9VGMN63Dj4cUS4U
sg/iRFlgD6bl74yMR7GPMffAA7wpCskxgLGVMwtRkJ0B2RcMM3VQ4rCgX6OTRSN+IhtRApUEC2PE
Hle8scI5awUZXaKk5hLnAOnnIFWqrC9o19eP+15Z0dDc7jS+tDlUoX6utIGQFftFC5a294rvupmJ
tr2xC2FxM12UrjE3FfSeOSS+hR2gpSFbylF6Y4RZV24NQck5f9YRXizf7VIGdvE5EgQqXHPHuPX1
LVnDrvFNJbtgPsBURbwLBgcdx34iadmg/LwLMBHa00R77e9i8PSpMkQdoeDPRtp0DzJUeWeqOODE
zmY/JqFM17uiGStuBnwm9Scah0AegUw1lK+6VobQ7WPNeWULqUGjzGCSleVxV3TZWVWK/dXPqNew
1D0W0rstb8VuhnmZr07GrXmP+PhE9+92+jRFT94w+KLq2ONbc63qJlusUobFfGHZ1/bY4vCJGMop
dJK876UcolCmJtD2Mwpqq9UbyoiNdMQ3k2A4Nikqgg9aZ5F7GXo9TllPMo0j4K2JaiI3S8JiWR36
xw2pQuBAzZZbDj9Rmt7If4CQg/lOpG/t98JPfRqFvKPsHHZZtSxhX8/lEQnDicUl5g/ZObr00vBD
ttpN0Q6EZEuZ2+O71v93jZMm3avXXsmVTs0axPNgq0hq0zfAJQT/IbEq90RNBkeMyKkD32XVCvmX
YtOObsIUidC4/vP4dTxlGLt8RsaKrVIPzTpbj8s2Emnns+AR1drWyc7Wd04W6P8l1T/gUajUKLWP
+Wtm+xh9x55b/lgWGjKpi4luaF626MzACgaI6DH1+OJ5seMBAHCOGFkqNstfe/IobBKwAqS7f17M
Tk91+7K9sUB1yz1kbEbr1N05QU1FmeAj6q5Xfg9dcjphV9IzfWSUH06587PI7oP5328SSmQmfjHU
xaqqV1sah12B1QFyGv8gGuiDg+2UJtGpbSn/yyajjcLTil7kQUzU/oPlDIV8bgTtnbMaGcKeQrZt
w2X20rg7tqQiTTuamjmFzl/doQTtOAliiBKOFcFPQsBzqsCMkpKW75m7m26ImUn5uZ1KqZVkDTst
zxe1pDPRGRQVw3HVSDDdh0csAo/scr4JZtJKSVZ+6sXjwz5w1gW+W+rf5/F2IWIEmEaYmJPJPDcE
0HmNYGwITNrspTpqs+tyqsIotC4rluuN6wbMC+L0rynGaL3AY8w1aeKoZGBw8Win/RUVc9dkUl8Y
X9Mj4nP9vcKAGXqcqahVoxDdmNq7DZmn4qY+HWxCZac1pkr6eswGXX8e0EAHL6bKCrFglZYzC8jU
3BdFEIOKjEFzqaqQapVd1tBllx1h6+ToTK4sDHUFHG4I85ISd1WqCVALrzGySOCm8db8QWEk+nJV
eE15f2nCs7Nv9+5U++zwUNdf5/hH7Ce0Jg/PgAutLjd8Sq8pFBxCC9Swwwt/Vm5nj4fNhr3KxlLe
vYjI9mVrcYOsDlktzrEMN78WJMZBbQcNMvW9zCJBywaHupxzXa9T65sXuEqp92dNvikgHkFMUena
+zvIm+u8Zm8cPGL8g4+DfsNAggfhA6b6dKIIT5G/6ZxLcZbz1OoyFOezxMH1gkr5M+N22ddV8VzU
q6EfHyGD851TtULDOarw78K36FcvGx3kXHM3YKob6Igvqa4fHn01IWuCo/e2oWuE3TW0s5G30xdR
Ofo/f4I6+EdI69i1Q19RjlXbdsuh6Z0z1574sLZdlxiGejfnKFA11CW4q7H+w7Vjjz7eUAgljPbz
bdglZzEoUOVtObSplV63BB87OpXosHnEB0/nrm/N9eahsdXPJ38acy9GmePTL+Qt1xH1YVzJ7jBw
9OJZPMvaFSLd1xZojM/BhG0/GOaGTpSUJdTpZdbjUhJgDJocoDMHJNizsRvU5N99bMU16MUcQtXl
oPLWmDjpVft+sY5jR7ljMqQ5wBE4Z/X32gO931jVdS2svTSbgaf/RewR7tfZ7o0YhZCrEE7uLO9S
j2fuSU1yWF6F5Wne8gMi4NlPzOy3nbEcsnDtc0r1lSySfHcQRvxjIzZDc9X/9QFtBGy911VPHeqA
Vp5Z9YOWQaLvN+xOTX6HNjBAuXNHKFc1UzR7I+V4DrJQZMoo8aJfeM/ZbodfJSIPSWR5LLtqw2Jw
PkIskwZhTePA7YkE9IaEVTxLhxPIBlObutnyYRQ9ujSbjtyABH5UW6fgmsSS022DtsLc/lj62+GO
i9Th8rkqK/fV6LZlUDxt58BgzwG1qbybsHJQjjqt5vt4abowQ2RBQccZUrLnaoDmXkB0J9wg11ZW
AO5TSB46V6c7MUHkcNEMC+anCqOE+3ChId2WdAbZWsJCmZzGS/FNEuF8LCz26Mrde9RKrCCPi1WR
DPCG/R1kE16DQP36QfaoXFkaU4K2wJVPtZ52VcCo3lKHwDIzZuD/FXn/Ow9ZukQFou7p1OnEenKi
tb1v7rCzub0PO5sSVftfVOGwGBxiZY6GsyJPjFE59wQ+9k3eVNtgwT2f3fBwNK2EU8iA4rsRm1C5
2MGZ412PhASjZ5uHoAI776BxJMDGWB8yfmmxe1DAQVwlXZNJcoWiJ8WH67F8h8Ij/eREeqEV2Tqb
DZ88yYCqXOIPzIjq4BN3uu8lW5uE5pD3uJtlmBFyWmlEI1tLcly6M8WJVzvWIF6uolWBACSu1xL1
tZEViqPQ/IcXeE717QZJFVse2OocjxapNuIyOIL/wDyWDrm0XETlSwoF1XrCCfZZJ799fi4WqxL6
L1NB+naiTy0sFrbMmTJ4aLAB3bPX2RwXREbYjWV62LWVxWINo8AOSZe58pILtZOmstXC3rRpIgND
rbdArynEgaYHZVr2wcEV/XlflDTMwCPvzWqjKmbR/qbnJns9M2QArReOtuJDbhIp+TmygaHHE68v
MbMIzx7eJxT8ysjK2l3FSdFk88JGFU2M0y791bdwBXGl/EAFpNNt9PHgunpyxQ15KZVDqhu1hVFx
ZdI8zZGFCo+Cs/YycRu1W3g6FSajlqk3rAfkQf7AA4xIydP/jigNZBcHwFExznehNGBamQmA/wT0
N5agPhRvMGdatlccKk5TjsFA4j2NcYkYXPWRPccQV3L62gWDg93bjd1QIiXEnGY8tE2B/jU7GKEW
jGQ8GfV4mNheviQdbbUnCDM4AAbDR+5uBUcDGHNOBcdkyL7SF0ugQCjqXWaTj2pz9DG5q8dfXVvJ
4hP6XcZAeNLUm9ZIVOqVQRg60uD3q4j0aZDsSoxvRyS0KEOpgi3PjuClxe/uLDQnRspqvzlNtqAw
bixnmIYK2o2m7QkD0YY4j64YChVDd7cOhKkqZizm9O0MQbCEPQIsLLcq9HI6B4HtjddJSJ0l0JTb
JdsWyR0MNnRyLfem+UTrp6IfgbDPJPN5X/U1+STmrB9IDQkmoK9ITv5FYPb+v1rDhDAthUYgNjJP
xAAhhmEvCeCWOVEcxY5AycJvZ3rch2of/XoWLxjgRQP+HtXKEDfdVQxsHZENpVHQDaR8dCGkMVmk
0Tu4en9O0KUq1k9kwpgbRgx0HvTIzpCmD/+lzilAO9zcVdrfebNQhLN7jluDI6hLvo/e4RVrlyV2
uHWobL6a9jDoS4LEew3iSzOL9mO10f2Yle3FNhkyJi4Zmwc2r+rN/qPW2zCaHzcVH1KBr0f7IAx0
Lnb/mXOGHzASe6pC3fUyXaDzFdcZB9v5arX8HdumKjihNyZ5DDGG9dL3/zS8eOr0V/SDadhdWxF1
855AwBLm6H8JG2JivUsKuYij3OtjMsmOQVwNM0zQvxXatKSuXG1njinoVVgPn8cj0ZCgH46USuJ7
LhAFp/ACmVT5d4Ja1d3zmJCr99fqucViLMol+mUAsHVAakI69szP/aLqro3hD2zok/rXedMCrLJc
xAfjcuJYjM2K9H9FJVqc1xydgiFEorFl3A4l/BrS9r2gloEzx64VXg6d3VjtKAJ5oM+oVMGjQwVM
Lj+3DCtZ/p/vieW6s2WZPbPLAVaBKnJLZteu/mlcJgAXPbee3Ue30nhCJ0IQf1PbgeH/BVxC7OIH
Dv0VOSVZ+wCk0Ak8XKvi5Qr1V5DrHJqvA4xazAN6YH/oaGNI9sN32uOZh9819gdvjG1nyDLDh7Lz
8BpNOm9RlFG+FTNWNqFxw8Rv3NVtS2qsfc7RDJNg0NGgay2bQvqQCgQN6S+7J89zX1SlPJN6MXet
ZSHmhrX1svvAP3OPWU7hwAmI51Wa9z02y08emJvv0uSz1ME9YbOarAKhSnOBbKLb2vtJPF4EIYWZ
xVvvJmqojj9TJkeEF/e3Jkz/CwBryfFH0bc2AXiOuwrr5aBZ7sw7byxczQ2B+Kxx4yKXYTR/IdZR
MbLRd96eqDLpNvgRx76MqtTQDk78GGhfCkc5tZj3dw+BhCWhAZYv24rAbsHo/FeSc2VGcn/c2sBH
xZ4gVD4eNhznS4enhA13hAqXd4Fwpx4PHKh/vbu8kkpPmIrzBfj2IuCEt/IJ72BbImcCGhioAGEJ
tGaqsZnRGyqiKYyugayh+L0/G0uTarKU2hcHUQUDvXZemDmcYghRm8wy9F75ledSbvOumpDKNXs0
ctqq7il7r6XboMYtWlIm/rTpEuhDqxhPtmHS4D/vZYOtrVsXMbS6vTJJtU7dZeHFVIP8NY2YMJlz
ljdZE5z0ftjvzVevN2Wc++B1kp0zvkzNlL3hlDuDJxHZe9oG6FrGUC3eYDqJPBcWDwVI8YJr66kW
wAIEfAqtnYIl+3aqYEqpDIlgIIcs10hbKU4u5R8S2aiQ6AuyQl6Aad5VP0nZgsgx3Zh/KS7P8zYn
6Md1lMzi3N8GClSZYUjXBtcc/7hYyPmd6umrIUWtlCVXynhjiDgV6WKm1LQ/uVz57DteXAJiyFWH
ZUvRjFIC+y917xLKRKwH5z43JfTm+Z0rrZnKkM2y9QWdwfms16tNLNvSqCS/qdvRRR1tzc6CmwvL
vS1CnVafxG+WOXaiLInUGrBaoROPI5QdR17De0KS+lSbPw0iPZ5ez/HzjCehHQaoqRw+GfGwpp7W
1zi4uAdM2w+2L0CPGSpBiKB8EYEtvuM5dzwDYwW3kW3ZvJwt+o/12omun6SOWHn8BVdS4RnNWg/I
0uzGaSXDXqVgcpuj1Rzsysb/LV/FcBTprwvomPTgUf1H+EMf/00ZrpZTQuwNThaNmIGRLbA6ZpqH
+JHadztA/c2pnPSN52ue6Qq8IKDoCWuEYFx4rJQvpNqHMkQ24PWFuwmrR/qcjZRO4MB9jCnS3WTH
rBYpZL24HblLOiFbLTn7DfzCYIs6gUKtxAHz8SddeMClCYGKvH7SDEja0j5F5pEpvroIShdW+ZTF
avBtCB/VDIErIdXhfywaLCnLoDlzncEyJAV1WG1SN/quJJMKdwWe2GJg324rQ9LmBWiJoKAd5ZsO
eWJxzu0q3tMrgkhnf7Mei5Ww10VncaOPbt8vtBzbXwzBLUXukbOMXTGiDsch48mkwbSWynMSHqrE
Y8RtfpuqXeSJXosL0LNMVzdk7Mz9fnPKcR0z/Quzr801w2cZXrJ8e2QEeJGVsP6QdBkm5ck1fwgV
YbOO5LgH1Gli5OvtIuQ3+UvcQt5dVo6P5hi1jQslG7rWnpnM0bWVwtLzA9ekG3JvVVtwkGMKBtw0
44e6GvMXINwZgTy9/36WgOqIKwl0NW6VJtNI7cvT2PS87lP02krMk45hh1xKDXfIRtVGsl1CA/vQ
h0RrxPrXGKnBncLrWsN88iF7xsy2PAKQ+F97MM5rFJsyHxNvuAIZTcdry4Pdfs2q7TuUIdj9gx1c
UBsbkA34BAJlgGieJEXURwwfYlqDOh/MVJIhZYh/KSrS2wFWmWWh9qJeJvSigwY2aAgbNJbo9hSt
fZ+QZiKn51Qpu33f3fk2xJNrC6Gj5yy6PZgtlHu3BmNfd8mDoz+GLGHKhr+z+yFZuBOGCqejZ67O
rIgRqC/dOmDzIxPC3I3nbB6IrHNwxLSaX6WWJhbeuCRhmidwNeVIKiNu0vCI/+zL8J2MTnSQsPxP
iB4SiuZY0ygJSdD1esmJdE/srS47RT5KHUou/on2NbxAYtIvO7xTmMbfkHDmzyzdai+nzfZmjEW+
+BqdVY1qqGDxyiLx6jd38kqUMAI0s12sIeGa3c/vTTXlg8d42HHk3fmhe8SKof6bECiFY3iZZiGm
DFqoR4kKu1KdMyTWtSWUNi2R/Ozh2/qoBz/14XBlUNJ3WWKh3Dn+z/mAYhTpt2cn374OMw+9HIZQ
NMM+ZNZ+1/iArzYoBTe6tE78O2f/8ohhzrxfjIU9Q+Qp6LbP1oSgPvVUMqk2xkeRUPDxyMl4pLDg
Z9lff4p62Wi8PWkP5emhe4VU8lNPapysbiBGqy29sQHLrt15AISl/Jy1f57Ekoq2Cp2T4p5b2IfY
al3SbfAtlPUa0PmLOWOB81gyCIaRrLx4rSU6HoPjNru6JGIUA1OzZ7CtnOcznV5Vm0edb2UK+4aY
RgxUyOI70eZ55DSx4sStD1ktkzNIzUPOTYbOHtwUib3G3tpBVjth+Wf3USA3fnD7Vais+KaZ+cyR
zlPF2dNyFttUneb/5+fSu/UXxjBkJFYD+3GY85jqEd0Pqgg90wHcx0al93JokZNP7836k6bC72PI
QMs3askNn26XSvCg0dG15fjRX8zUbZuYRqM2+g2F55R5ZAMlI3hFugSaAdnOVHiRDILqYhL0KeEo
TONC4UBVpaecJl+I30Wfi/qHDk2oE4aHhP5FxoPQTFjA+1Hg9asEZje/rn21VAr+2XRv0b9wsM9v
r3vXJOApeJE6xFy8sYAn330a2S+hIO0n8kC0FvdQJghtSh3IsbJoylkQeO5Mlc3a67LCT3pXt6oS
GPVaIGNxYTZ4uMtbga6JQrELKvi79pBarRIoe5jKePEKcOFYJx3skAcSrC4naF4Sb+h66jGCslTm
qcWJ8wiPQah1hJvVdFy97eEuwOfzOXKUUbnb1OmKJyWQb0WDEWijtq1OXDX3Ksz8LpC8tfxap7Bj
0XIPVQfHglIDVc0wxunyHYZC6F5D63+USi1DGmGJBAp8C2Koc0YLDWaWwx/eyhEYUW8qtSAP5m2S
NvA24SSa2uiVflgS15Z7zfUOYM5eRkfW4rPHCYmJG6rEhAhCmp3A0b+Ts1/BMwiGs2Pi8phwFOrL
1+Dywaa2oMM/n3pw4TjTSZdqZ5mLw3xkMip+M+boyKIzc1Ujy1MrS0tkb6r75dhzCmqJJoMzJMIl
2llDPtqbdHOt9vzOocCxyE+dyFdnLIIGQvibMQqniC4MeyBK/k64RRodPHbt22RJ3RCIPMJLJiM/
eEX2HAEp3fBsa94AdmXRhBNOgbG0khRvEsfQr+57u/URb0QdVXk4zWe6Zhh6ouueOHP8D9OiF3h/
tL3hKihsVROwCvOV0gwwoAjGZ+lalxVZeXGW0taTvG4BBUDHYyaUWUopDTQ+lfL0nuaXLzuEyJG7
1r3FB1DMGJjidoaCSL3UvVW5pe6WK8MhFn11yCjTMeruvjzj80Ry21gk15dI2qZuTaf00VlMP++j
D3HjYpYIKSpDO0jXFJHMCOW+SOGk2g0RmgHsLwo0z4GxlMnW6hBPEaYSfjJ7zrke9Zhy56NrcDzF
OlFYp27o+q2TzSx/CL99OV/garGx6FK2ON+3Tp9qLB9tkxU74X7PbVbRmWq6FAiwFMahZn8dAdoj
pfPGX0eWdNNhhAtkz7Esi8Oxvr+Fhx7qh59W2Xo7VQYfOENjVgzGA17jADVJCUO1rdFQA3rq2yIy
5TV89YW8eHZKwr7AmvVcwN5r75e0bX1jgfMC6nRgmtAoEIv2EmvwldVqo0eb8XAtr2pQIWodH96E
TLGC8lAG8UhtTLe/c2vIJRCJwd7i45dEBZP7TqxU3qx7f8Bnnj0Hqn8GxLrND7AqNsbezluNmB3/
6d/ROj/9qDzYfzWqsU6l54NhVZyjmYWgMHLQwdArGJP3+Q4Cxf4KKH1GGiQhvYlBZGt8ffu1fmZQ
Qk9uvLEJ4s9fIN8fwj32n85+sLrFy7212wFWEJSOPVthpzAaF4tFjtvIz1TH5YAfJ+FolhysqOu3
+u8xasdnqT62kDWArT/dAUE3u3lzIP7FG5mZhJO3DzKTObUciowcRPEBIpMI8CEFYJadckWMxUWg
kQR17sYIFEpL/j/pPqoX5OhGvS8YA9W7QGNLY24ojfy97Z9+w/oYlceif/DoLE/Ed3/UJJkaOZH1
FuJb4Y7sPKaZBIGIDs+N5kfGJeHGhP0XYc8oOfYt0ZhPd8dmMfOTSqaGXDP+au4IiDD6r48pQi92
9gVnSPAJNzCp4uLuERWbIkQFYv/VmCpAsfOFsffVmjmyuZl/meLdr9zmuOFesESV1H0L1F8whgjt
sJ7VIFAvvEKGnfyJgiW6KDfLTsL0ltv5yytldA79xZ8Z9MPCo4hyufQMI3384vrAiIBV0zlQO6L/
Kz2loCxcZ8pkJ/Hf0AsWbMJ2CM6cp8DHUyiB6crrXnorNe+nRhpJ3I1TYrW3ZXPvWYb70MYyls7C
gIIj3Ecqltl9nKxccJrVY9eUs/eM00eZp194UYtLsDBz+qGrtX7MixF5A8Q9G9QFeMd6BGjVnDCp
1bZvYbrKjut400sAOnrXnWIy3ond77jV9DKd4jaih7OXo66BkhgYh6hrSzNrPnxVwYIEQi3/9nLP
QHH3rCNDsFz84q8HknWzfFZuMHDuStyQRNE1mZIjCeuGEtoq64Hv3ECroPtr9Wm10p1JeUUm+Chd
EbRZXbwoEpHC8kwB2GalWi/STmmAuH3TfsBYzOO++PswDUQ7mTH3vf56ZoZyNnC7LA/1nRfhvoIq
F7TrzZSk8sp3FATYsTPfJ+/hlYVQ8ELxj655i/VwW30h4cm1A44XxjUEHusgqCZXBFSs5ii5+0zC
Ly6FOYWW9/4/sVwFoJwUs1I2C8qcxz6JlAOmWixLsd3arAmaGaPFt7N9kNDlQUFjlcendabDbDDj
tGDtIUMPN5esT9JHex6LjcIT7YgUxD/lEcKV3r4Wqbm0SsFJ5OH8VN+wbftQX9CIuFX9L53n9WGV
NrcSz6cYGTXy+Ibndm70r+QMMUyJ5NKcMb9rlCtCbLiYsuPSMj/2uNe6+bB428S1PeUa6R0H3Eqo
LEjmwnBV5UdWF232ZgLcuRhwOzRN7JwyFWWUPEu9+khW3jk0V/urH2/OeKeoQtWUV1S83mq5Zdt7
y3XZxYRi5mlbEn1fIthTt6z+QiKcnriIu0rNi4iRc32sYXyDBfOUjf7j6TVNo6jHVVCfrXmNYA9k
4hzuJ01S8vQctId0MiUzFcbe8XdhdPSQQfZ0pueoHt17XZzj+ZgtsfkNpT92AF0pAzyNFDLnRanR
FG3VHHMA5gvctdmdXzRI6zXgfx4mSl5pi6RDCF+RcktYNdW1Pcy/y39UGr5Qm/yO0D6GbWHarkt0
K/cKyKgzfvsQZVPLI44htOpBJ7R87eELKcEs4G51kX26hlEKe9t8/XJ1V/cbmZ0Quf0JnkG1oX8V
phYus/XZ+WNuP+OH2ZKJzonyBXxy5fmUHWciD6/Vt7B7zgan/FYsbw1CtTT5bRHHuuWBfSLgxdHg
cB9MWB6j+sqqk5WgvqdUxSxr3z7mrOaHwfztFnrf0iSLZdREAGeQNerLYGbpiVBHNPthXIHE7joU
NryabM0P01/echWiW1YYyl5Oluau5vfA6HJJ8tsEbO/EFgR00fygWI6EAqxI9tFruohCiwFmF9Jz
HloPMfkwKTn4Bu11uKmwMnFakl6k+aN5lTmVOWREePRIEiHfTLOcs5KB/239k88oVhq+PU4jN2jz
8S1miqA5FTXCaKFCNm02/oGP1OEYnmHyxMLPXaam7pCIO5ikoEntqFUQ5+bD4RVcedGHd2t6bMDe
AGDN9dSg9gR8S942AbHMpeZcsaaiJF8EpWcbF44vd3b1HSm+ls8G6WAEr3fz9DZ90CVR0+0ZQn3o
XL+lgz+QIF1wdHJG4psNKRIB01f3v1LxBmgggW4K+tY3IM4wlrpOapDz3qy3mGbpc/zA9HjgQMUO
Z1PvB1qEuk69S6prTaaWjgjCECAgSLeOrbCDVKoYQk46svyFWirpYcYUDNGKTmNXBviHNWJrDoLB
gYWnA716PX2kiSA3U55bOUFlWpYSvAubGEC6wpZ0FNAY5Ppl/PmldgBqnaGLZJDiSW7TywwS5D5Q
2XkC94WQXmCXAt8/Vm1prrjodL105LnwdxqhZDJ7B8uLGGhS7NwU6d3AmRajs6u0i/6WFoQYz99N
+ElHb5C/vB+Oj2kjljMpaDsHmZUN+b6YCCkoAmKoLyVGyR3MbGvIwDOrGjU7cMaE7EHj91+5O1ea
GCbUKCXfTf1xzS9ztCsi1Po+xz10YedT64TA4y90BNNSed1xbAVCPjSDKOhu8ybsX9EwFjRzvtfa
Iy4d8waDSAqVqqCW4wht12pE03wnFIoDX5/CPO8KykoNkgqmiX6IDPDCZtfQx4P5mgnYUuW0FSpb
qTEaRzHQHecLkSCxAPJmk1I1RTOiWgt5Oq5NDIkyUJHeVYhXXGj+etMgJNW5SJw+YNjZXe6eD+0c
hSogZ6heX3tgPU501ZfuHIcTezblEmPrRp2yYZQLLghZDKC9yJeY5yXU8dIFEQ2mJQXzvyLwwA4D
RPGuVS7y2VPfaLEJZb2UGh2XhGvyS2piKkYVSSuORnXMcqF925mgj9s8Z0+ujWkJB2fnIVrbzsNs
g9HoVvae/r5lmGEIFcesyC95+21KQmqBWB0HJnmh+yefwz5OP6TXCwnXf+6p8QN5jRAEy8QiAXar
KtQUK7cFn58v+D0CrgefiYZh3CchgmY/Y8DPnkuCY8HfQ6ABbgD20d8S99RM+5Hz2RzFHjKq+WMy
J3VS3YLwSDKVtzeG0uuEihhaNOPQ1lQt9g1QBrcGqRDRiSouciN77Iy/d+X88lbXoQnhdtQpoZ7L
YYrusSuLpMtjq/NyGWhmtidjpKlXIahxI7HpCve02kDdj3Yvd/KmNUpGOgJBh6jFSBpG/IrdFNAl
EescRKn1FqdIn2D8f95tM064DH5r6exhjOq6CP3XIGLzKBvRdE1dnMrQCe4y68CYU8m9Q7njRlAg
NnlC0miVBQ7I7KhZgXZ4hLlHVVF9jaRQ0C1QDBXTlBdc39KOPjYKs0jAiJ78LnAkM17QinfA9wf6
l54EXM+dX97XwWewNY5JaxxDB1A7GSud8ru4rB7kdbfyYbaIlJ/VEzlhyMXPvhGetm8RE4t6qkK1
m5ZErP+Ohef0PaWbSAv4kCn6Tr8ItyNH3j33ExH7Nmjv3SPfY/Su5B0C+d+NRbxbYw/+q9OSLSxE
OHuQxB+cs/6DnmXBulIPOgvRm/LttVOHUSCs4dAmHimzWsNqK7InEJJEeo8aB6MAyrDOtOJwOf8Y
YSrBX8eVP5iv3gbAe5ogn6DztEYIY++0ydMVNZc7iRLoITvYIrnFstQLdVJn3I6pA9CKOmsYerFL
/+EECCQRn0/0IOmsFWVIZmVabKMThBaTJOeHOD6sXouREDQkjkorMNNOnxk98nbg3nVJvHA2rTeB
Uav4+HpDwn5YyH1EokPlvqVgjtpQBtz4t83OjuCvHI/45AL/kYvWXFSvxouMjDYsYli3dG0nmLkv
VR6EAeOG3VpnRtPDfxo8MBkks5Vhgh4rGbVgM4BvF0UOeRaGZ2hXNTjuf/U0/+NdMgsZ0u4j+82v
WB11vYs7pRv8ubHNkwpMiv9/BOjsjjD9Qi7IQJPoiACbgJxVUzQiJHmdB1i5phHZEVPGs/wknKwQ
PP7MddZOEiwvU+g+wLZLB+qvuzJ9KcuP8WeRsrL9KYVXDJFl89IOX5NGYCnECv7oX8iWO85y8EMw
/U1DtIOcF5t8e2AhWVNk2C8YC+1Ndy6YUK/jQYpWC1w1Z0hYaUt3L77v37NYAmoQ3mLCpOhoUk2O
zCU9YtmllyMSaEoErPQ4o1EOAlMDwmNqG7ST6kL+hePPu9oSigxgQMYTelpMOxP/tyTpOc1IUfrO
jLRf89XB66Hj15efeZ7ltNojwgPKZBojCpunixOPSQ5BvTlcgO34MjPWtJwJVabRnaXnN1jTj9el
V00MbkZfpveCaJAjxcWSFeoyTUv8ahpb1epeZzRriBGmDnN2BjzupP+kPfMlFBRG7ODzSlOB0urS
bbim9Ex5IA+O8+2J45wNr7lxNVdVNRYtc6xEz1dhaN72RjDWv0FyUwsMnHCfSjCDZ1NnM4PiQkPi
kY3BPozW7FEET3wf+KMw/OB8mrXn16jIGUiSvrEw69xuJXWCYlncvWZbs1wywJ9QnFFF/iStdWPC
Q/aUeDi2Ghe0xd4nVmd1LNGOwg92g3GsFnuvhBgc9gLu0EmdGunjjdDGOUKog4KhV0kK1a+QeBfS
I7/BSet5B7DQTgHDhIYg7cPpYh5TQ4zgGCTQOBG9j69aasEnhIvQpWTYfnHHrt38GPCsQpFdAa7r
yOy5TBcxgNBsK7qwmJ1TRVwQjGkjpPeFICvlBD7GQmnQ+PKz9K23htoydlYI+xENZpHPMWXkt0UH
IXwupFQQpGW64MSM2P3X6riLCEmcgQod1zX58uLtq1Bs6jgUYGmndIv3+B+T9c03DRRLgXSK7pS9
IDOdbt6tcDvM3j93run6pEg4KJOfrKDJZAVQK0a2NJQvc2ADuIVfKkyM9zGS3kcFPmhGtxd6QRyY
Y3IVDS3jPr2Yn+UgS23y6ejziXwsi0hy0Q/ClIHlYjQ+f4pqzYU7RQq82badk4r7zNXIMG9/M0rQ
DjBHinNn5RyM2v0OurD/5XSER9ycEWUjxZ1Z9TVP5Fl9fYTrbLY4U71+Swf9FGxRPdNB2J4TsInN
MtiekkBzCOKsocYcbkGaC33pGYQ8SN2Qc06B/yFC1wydzQ1efpHmCRScN/qIQC9klXnm5PmwPljE
5byVbuGEjVRzxbwnlqS6W/4tKnvDDlYIdK9P1+fgYuCyQwnw47zbltHEx9/ajHcWFvXeJkWRh/GM
FtaoIfmNY+FA5/+89YAtq1437duhCP8SJdOusYv+/vZ2zKdpcIAuIT0v4fW4ORE4oaFmBoJx5HwP
sn9NymwDjZPE9hqbB0rSIzmBsRxgFrdbpQNtlYfM8yFqUSQMH6Qu7tyOToJUhFIaOYobjVALeM8u
G8jHAe2TVU7n09WbXocrw8fy57/iOxyKa81oXG/azaY7rwnml5cJFm4bQSgWBXvY4lE9abgH98Yl
qYIRGf27dk+zNalF2+e52XvbQN7MnUMGDUHQHRUW/EcJO5hT4PEAyj7PkGwMFlkOCCDGDt0XobJm
1/GvcMegFMjsIZIG//edeKCrdQ8qnXQz2/st8SObnCsOL924CHyPCXZTL99A6ys9c1O8538nSur1
4lvU85c8BeS1Z0pFXWGVGpDWXDQB087TyyDkDUlAXRB4nmM8B6GY2f7zDKiYTa6rU4dlogD2aH/D
2wFHUT6DwSiloeziXOHku5D3dG0b74jd6+vtuRJNDAR23UBGuGykwGTw3si1nX6k+TmH3neWkaU+
b1tfx8mWr4PjspMpb3R9U9wKGJ9wjtHHF9v65TVomIldvUYMUxDNzzE9hScsqRq8q0pu0pCPxufB
H/0FbfWMqf/vpP9BE84nYup7gY6k8UZWwYp26i+FGvz/zgunLBewKtFlcE7dnIKYZWiredn5juP9
02AyrnJAK6RX+EkTjB/c+Fv9M7YlIJrBkEiKjdwoziBH3JPr3xYWAN4GuzWQZ+jPh1OdCs0+Veii
HpwDt4Lqrv84/O4lzSbXFtmkwcN1hOsKtm/a3RyPmB4RlzxOEvmsbspOhUvGg3nVmeH3HpRw5+3G
FcXREGTtaiRP8clWjNysGhXCFtNQczS2iFY84c8SQsD++OVQc0XuN0xxDs2b5apC8Qg8IpA+TqtS
7dNvBjVoE5DEDtmlllxKFh1Ap/pG4ecTCpQhWwIyrmwS5B9OH647nff0p4LIFh/dQq4BNh0fbSlR
ScjXIx7+PqgpsYt13s64+jxZP0nzb9YIfsZm2pye0m1z3XXcfHZ6qHnBrQCXmmKWIIZdejQzgCpc
9TE9Jt+pU+jfOyqHCEPuDtbxbEN+UsRXtLjrANFe2C6n+eOI2uGJarqmaCxyZQYSy/nj5ASte9KW
3b/rkMd/yWndCC75JfiKcbst+jE7OCSy1pgDRNfc0etB9f/Wm5FZx58ctWwV8nfYVGW20vcLyk7Q
GcJv3mjEju3ETe+mIOhBwVkIejIAK5GJV1EvkeM4NEAJ8daZYgi827OOixue77luq8c+QUWEqUj3
T3VUxh356bl9Cr1+9Xek+7Rp6v/GUEHZRtMzZsFZPhZN79VNKAWFFs7BFZWHV8UUe+3mjLWc3OhR
q+H3n5h+X9jpQKn1+XRxahpkwl8ztilHJ2cpDfAm88cwF21fl5ivq2cQAlHBQMbHS9nIoCNhly2z
uPpabvslgCeXoD5Bl4C/xcr4Ycd5TN4wyEvgVDQg6iQijB4v5l9Gd1FIpD7CJY3MWJvU8NjKV6vu
Tx4gWDYLYy2zhiv9EXClk0zCFeaoHJ8UXiqI3lKhM/yEAhG/Ulgd9B1RGHUvqIc+QYQ9nx3IuEtC
pQ3JVoXw9BwCgn7BBFhfPOZDRjxllWB20Xhs60XySCEtWNC8xP1cuEG5NjBrkcDS/X338pYMnEiy
sqbWnzASZm0et3bzMiW59i/kobOrn3wQC/ARpBksZPQzEN/5xM7WJsJtyXRSlrog48G83C/E3hiO
T0abF1qpufzz4w+T/QlbjxeDwVpPoJjuJHg3VUtG49dz8KBWUV4FLiNdLkSI/DeG1wO+oL2C/4V7
FQFoeDDQKoFc1PFGmLvcmj+EFroq2H0vaRd4+3E6HsGOleKu3S6GkxL3pyTimvqwxXaseKdsJy+s
cAYhiXbigPxdBb7ddtdTpC2u8CAOXAeya61HcA2UCo7D592gmZpb3Y5BFG9El/+/5Ga42ASxDb0B
uoJs654Jo/tye2bUdEkrRnjPKr7QKnxk6rmYym//jtlQzMWWvZz9mtPSlVnaGiwAO/10kv7nqjsG
83brtQzhEbPQfeAlo+KXvLgytSr6+BEzgxgHEknYkTSCFuzTh/BbwHTMuLLeVkXdOSIX1zGrH2mY
L2WCsu9ZV39hNI1x8Uy7c/4DPZ2gBJw4waZ0xvvYD7k6IphDbm64Ffm9tzzDcetZh/pHiYnXUET8
FceSwX0xrBrSP8H3WeblePwGBoqvAxrsX8SP5T9ktgMQiDo0MV/hF39Vdx5/Wfn+znF4Ps/0sFrT
zzW3c3VqQLYJ547tyxD4jMqZB6IEoF/u9t6LyjS09Z57uZJq9MX5tLnsYqulPuQqLlum2nxU9fRO
PD++9MD/1L3Q08geBd+gveyueq1uNvfeFq3z+fT1wGqKTHMi9otTCz1gj14ZVdOY++eB6kinbICa
y+gOvXjGktKoDjZnujHunN4xeNoNb5D+L/5GQdQf+0CYZrhrmuP6G0rZW/AafuVLAFc+97NYgNVd
QYtPddJswMteGk9KLWHK9A4JjVgV6zCo4qZMtjHqlkMXZ2KBirb+GVLahYMzLoLdbIP7FvWv/s51
WNumcyBtudOwr2V5jJ6LBb+ZqcfNJtSp2UvylSTwjAkfitcc+5Xui6cj9jV5BCkI6yQW2HJ5UakF
7YASKmBxCjz2AruTJNr0cPXW7/yzSqyUbmIgBqQDpcaK+/jjEoFaZ440XsFTWVO6LZ+ox4n0qoQg
EPIUSpHouvrCL8OeIIe3LvHZUUbeLqUiZApzzidKeRpKMd8fZLAQBearXqG/IGOCwnQUBMaENbvw
kJnkKkZ6JnXI9uza3LoH+h5tVFIRKivNS1xeVk8UIS7oW6LbTwlKGax8H937ZrHAkdgWPzWSukDH
tZHhySSUSS5iAIhMUpU0maau2khUAJcZ2n/v9Cb/uEjyLm6Q0VUgzSSaoylASvj04mq8AHI/dPo3
4WSpl9jnQlxZuUKkzOlEXVbleFj9aFxzTmxSWnqp8mM8gVUsE/Tl9ZNLFI3QHLcCrv1EyXAli5yF
1kaoo6bGvdbhb9vS8BnTXMKejvbaoytet70nBpBDGD8PWDU6Dq5mHDyew8k1ST6Jq8pIVDowdkfm
oR3Y6AZFE4Js5zYffN9kcXopKbRyzjIcair+3btCQAeOUORHkCGZO6ab+88Y+GbMUAkn7ApOYtZC
xjR3v2fEg7WzhbTJlCGh986ooZYPjJVA5Dk6z4FvejXP9lHCH4Dbl8uoYnekfBOS84U1xgqehLxy
EQunysSe1vCwXpGbtmr82ImpqEOrf4jKeO+hE0w4ph5HS+l+kvYT7klIyf3MjVE5bwmg2ypwFzpr
nd0ZwFb9ZCs9P3dFytBvqoGhCcBkxxXpeeOy75M9OV4B4jKR4jLHlMg5MOgZ/7wO/h6f3OyLjkjZ
DZfMhwlwdkbSA8N0ES/+e+vqQN1Xovi/59qM9qPR0DqmpyE80bqxCGwdRW7h2dWGNsaIxtX8Tdpd
BxmB7BaUNuFcqNu5xac8OD3Lbt7eIYYKa0xdK545CyMFdz4IucPpZKHYIu0VZrnHkD17wrHfFcYO
PnrEc6X+cW+IDH74IPs94uxeR6Os5gaQdQreXYuvSs+yK2SH5JRw+hnipLQMymQclYXd5VpOmUk0
rZAt/MXJk27F0pPeFpwdO7jaFIFV0P3zzJgS2C9R8z6MA4uJ+ybJ26oF+2w7xervN22a7M0+GRuj
nTfvdCchMmpz5MdYzN/bDJDgMPJXWqomb//lqALjifLUoXCax7Fmldf7YVXDNqLClrlLHRe6cpEK
7J0JeiBiYNunWRmhh6aI64ZygJA9M7GAi+UBBCXSJ+vwyUKE7RISbgfzht/dAT4eMvGO4GPzwdaG
xO2N76s2nTiJP/fOrT2RMwXB/8IXKw9S6SuZlBHOflD4o/DKP2qC3BuBwnmBseiX9Snux76CA92K
vhK0jwF9kjGriEK2bcUi3q7PeAPhcAMZLBPMQ20tpcR5mHT8jX9lrae0bO6CPkBoCfaGyviIHZS2
daNRFQkmKfizpGC1NaX5ejAo+yF7tJUsB7w55kwHxPxLBPs0hNLWsudkQC9Xs6Wjt6ATbmDoxSVZ
vMQR+SDe9LJZnXfmTD1T3Bt1KKQy0+JPYHeFwCT0CB2q+i5We+5onwTxUwwa3Gd0jIM2at2iB07y
JKowKGE5qhL3ZdVElR97PP2J4dyY/TOsi8asBfM+JgyOdLGHcUt2VnPTPwaQpVmIXL9kMmjuK4Yf
CfS6Al5J3TTzv0exTAPFXv6SjSdNtywIGW6SsEzB+khLQDgW6Vvv66q5L9NVhs7OLuDVM8VQFg8R
XeWcg9gfZ5SqvQzudaLNiLkm58ivRxIDnQxcGHpZKPdTf+QDIWXOk/od3bM6hU/x4f/xu3aQh7pt
FRRo5YykZxv+7JduoXizZUFhTdj6MayVLHPfBY8zPDO0XBWzCTiJwR+HeRuaQcfl+U2DQDXgUQ+3
YrPcL5mbZ19cyl2npVqxZJNoRtCoKNdZNxENYcP7YMYCApbB0i7B3o+fQ87PRmhKIQMujbymHYqo
S5CVXH1Q5EMOQX72pl3Ml/g5O2u05XoEautKBi/vIFPCIbOVDIYA97HhLHs8zyJmkD0oX2Jm3d3K
7JpttVUeRsOxbfi2qIHStjroTqcjXgvHzAYt6UJxJPRRlIBhfOCIJ/G5e34xvowW02rdHoN0Qqxb
S1yd2sPKBGrjCkgUrEtN1OmDnuZMRDwqcXRasopVrdAZ9NmPbSjmDExFSGZnOihm33Ff5eajZUSe
Ukoay4AKHWayrqbTbqgCxa0t8s95IAt/WXCZ3CUyl5+qdr9SCGCqXK1/D0mR+NqkXbhEH7BWRFtJ
0EW9drV78vZfJR6HI1MorVsIfj6zVR/paNj4AamY1cfNvjVnQ167pYqrD3sNlyRsOQt1EV4m6s+o
yweHZ2AeA2B//7A7NeQSk7FudL6he/pxPbCaZnc8me4t0xLui37AOXJuEo8xT9wlkBl7XO7hFKrT
RDkVoFuM05tPTMg42gF7lldfpjNXsOCK5YE0wVa408kZGrICQrOqsXHfGXOyatrhqiG+KP04TtOO
SvdSGSeuQBZXIjB4csp53tFk800jLcgTPqHtzrLylR3x1m+UCQ5x0Px1SvV2HOuOIVNvcMBwJ8we
3WgZ6AY0KWGbFM6LKTpOdvkAiyV2YJQs2T7W8TzrwS8UilrUoLdM2UBIvt7MlXplFLFl6sHm/wne
H2OKMIubjQvq6tsQF8oouKGJSw43cGmbIYJhSlsBHagPUr1zc2kOkEfs+b59OgwHYBc6lrYCj1kd
SM6DXok8pg8J1/eOnX9wltWMeMfOBwnSNlcHwAqaVs1dTcMm1KGH1VaBg5ZhnqLshtS8nZNSxP+e
dNeggCBnsArwvp7JGDSmfJbALwgxhoaCAa8FJTOg2SRnPzctDwPMD0Y5qQyaIUyjVUedGDcnjurZ
qSf+F+2gtBv21XiC4c0WXD2LUE6P4m8b0zOqFLOOdwWbubHNYIRHHZ2stD88cLM9kV6xQAXQw8AG
G1p67MF8QqXH7XMdYQfF2S301VT1skhucC+rzCl/oMgToQJRAyLccMSfr00cA0/8dypwDViLYg35
imInalFbxW2pOOBmcauCAsLOGbKwMzzGPvECftMz/XObTjKBKW6uc5EdhSUkUgCSOh/qdWyPKjvI
Y9vIppD4SYW6W9+CATFNii57T8AyMBv0C+p9nkxbCz3w4mDdi0keoBv3+4p9R1P2Jl00shP/F+Wg
YQvB+WGMlLo+T2GHPT72GAiF0Rh74FqtMDGxxyap1mYI3FBile4Qz0Qsuu+PrLu+AeE1XYtWmj/o
JA6ccNRkzjuMlFTUfi3dy5qjUzhT/Z343ny2IRYse6kyaOGPRKePfzQ14pm2DHO/JbNc1YH7KVU/
eE9F4S9HCIXZk/5bdYSEFqv1JNJ6m78BTFnn9E+4GOS+42+5NbpNB2ba/Foz5F3AtCroXGbhTva8
XI015DSXQ3BAvg1bhcI3bVsctG8hbIs+IbND6wGI5XF468IBOAUgxI4/WqrAp1U4U0VGljqwrr0T
oFvyoHMcS7FoQ968WMksXd4PZ9BzWxnZ9wAvr7i5YzFMu7NVYhtZKaWTnFfRBWskerORSZgp2vMa
cnc8XWA9KlMnpCOtZI53BSULcR/03TCsTkQm1PByYD97oYhbeOuJihje+NmmxVlUgRdIaCl7YQq9
cWHZ+24GTvYkbQxuUC9NKxZF5V/iCF9DzFjWenNDPFzLhrwb+wE/VHXwrOWtdNAOBSuyXPGEdT6z
LIypd2oJNiTrOyXBOOBCEtdZ8hld7LCi8mYJOSJe0kypP4J9IuyRvyb5SLnAfROvyhW9+nP02ivg
wT7obtcL52T7lHkEs5bhSH5mZ5AsKLPiu+JFuqLmvoRYUegyt6QLIr0vPUDukhF1oiXK9wiNPJ98
WxSIHXetzZR/4zcz3k6/ywU+cBob6Nku7z32URjdDAE2EFP13HR6is1F7Ll/qTcjDwFUNoiYYzFN
Z0DAy7kOeVrbtOMdoV5kVTf61uq0z7sBc+guLoP6aNvbjfCUMvcfOT8RHT9mf99TZT3aBv4iY/ni
vLkdQFW/3iw9Pe0Ue8uDZI9jJClsZnC72SEKM31qKP5oTHcP+mBM0N4WII+Evnv3b0DGrlM63xks
dBEriszN0csnpyydB44g1kRJRnpVs3t8sVSK4uR8+VgiNsY4DAzMDugB9t7QXqhR2D5h0zv0fyFL
fOPKjL7vIEx4EuoQ+6LdrZ0ZDEqFFQms5+N17Ys8gY8V3027OyCqzL2nDFFJnlFRdOx/Dq3DDpBu
7uw7YWeiS8BRi/ZUxnuEGvCkL9mcVWBk3MG7+X54YXw2UOmOgPcKO+a83w52JschHAQDt9bdWjP2
U2qOIJO16E403cEr/XB2k0DvJK4TqwftM5HsTmvvoMAKjB//8XuaQf7ahg9GTxVAg7G14KSEGF96
DNWinN6UAqZ0AWj3D/8YBFJpEyrhcSZt9wlFAFd5qJ5iS0sZ7b/18aaps/YA5Z8ZRquAbOtEBLTK
CkmW3aGYzdHEqljGRcqJ8qGBocSK9r7v/WHDkmHziulM9p9E/km+jv637WQ5oflqZdSO4Vkhv52g
F4272UUxxcDUzSvKR62cph9//Aj0p3WmS1Br5wQNXNu3xKLV79Di1ILWrqy+wocNp5BeFAqMeHYq
kt6upMVhQRvzocRo2462PE+lKHY5+M6nshZel+PM+srvVQvokxjf8MbYwb1QcFbh2Tkk+3BcO5ar
JlvSsnkvsKG2qLji6TLY2IOVgpUsAbLAf7i9OL6US4ualnNFWZ0RVfaoa8aQ71bRhZxna7W3TKrc
2luQOhW2xmsz30UdIWUk/QEMRqXhqP2VUdo8NICgVQlarNda0r95nkrWT6sBkjLMO4Wb5cp0rWxF
v3hL+SiFPo1Wp7PDbANccA8ij99efs7lkv7OpxML2Tu3M1qQMNsVKZuSSPYrGciMb20ikoTNX4zT
Bcv+/5JMvNb/mrXk1akVEDsJ43Rk5rM9EQxTaNNH1PhloBE2NASIuTSYnJNZuN7y0NNQ0rU4UoGl
VGHL/YtB+WD2LG51VTxjv2ApZKuLPwurcqTtBmvy/UUHaA9opBqoLFSYrhqZpL2OJ2HOrIgnn0tb
kpUnl3dmEmaoil1Gcbl9XHuGHMyd4ibpsPDL3G7N2ab8eVsIdUoQTHhdLgTPm8nfm1Le7AaYBF4r
8nphYP9r+wcq2lpwwf3CT9aMlUEAA+ArVcdUfAtu2Wod62eTcJCgoi3wmkLD+NfHDM3L+EiJEf/8
vNKbG8HRYD1yq+IicP2r93zlf2+Jsq3KoFDBxvXStJBIZ60ddZnx21cRwiYOg3PGo4zQTcpmW3zZ
OWHJX6NSXukjMnVFq1yaKDqgZOA/zfcswoyJj1ftALi+5xGHD9PhvKgB+7lW5OoPsuZUrUAnShWt
dK+d+59mklYIwct4Juj4v53+QXkrDEjrbnHzPo6QJW5tmBLfbioAJgSacCc2mhJuJoP1L3wbGK0Z
+C+aYFiV8p+LdK4AsYalt6wjykjXXOkny0OlOv8TMLJIzK79aG3NrVrufb3Jgt0mLCCwaACnCDj2
HNnlNN3JqM5iBN4u9tf3qwEyi61PaNRYmEdfpwcYg4PInX5WYCp5U/LYGJ+XSXf/UvidgWTaBmEC
Ulg3j2rDqq8iodke6HK8RV7E1Q81f/b3W3FJMp2jkIO/mmw/ZyKXg6zII58Rp9xQlASdJK/O5yeR
t+6wBqsAmwl5LjbFo1MdSIPN1szU2t6PrP8i28NfkYAkqvg3Mb2BMFK33Xvwm867yjI/q+q/5DRz
S5qik8XLAqCGajT9R5yfAvIRIEkRhXuBlM9baySx2hEfxy51BagdU+J7Nkm2fYxzbzGCmw8Hp+15
+BjPIMlqvzsKrTqxVi+jPW/UqfVIeFz72dOyWzU0IXuvupxNX7l88wWAr1NsDPaE1oz29UyunNng
RUJUTGS1xBp263HMNpdXLjEttk+ulHObLiC9bFQz39ynlgZqVLG19hTsxK0EVRAvhFbyGw9WaTdZ
dW0LrDiwPeluhlE7hjla6nS+HaYSNTREBnJ/cMzCbKl/81A2iHPoK85lrCuEEyiVFRjBomdBxzzx
gmYbmZ/o0rRFivlzVBOr8XcCnmLUxKI7qR4BRBeLvoq4i69i/jKli3QTsv/MUE+keijLqtwPDyu6
E8uDwXsrP4pjopi6KFTK+QOn9dijpnsZSwWT3zRJanP2MJaRp/OxaQ/JrivzAk/luovJacYLsS7t
oUR4GMVzI8vy+1DpU43GAELM2a3Of02pbPNyi1B78A92BEbyJyRHCN+j5FGnBqdGPCALvx/9wls3
q+jRByB7XAkJVB8AOoJz2LRhGhhaKn/vadpipBLeeDHH5fRYHOJbTO3yz0QsoPdOqdHHtJjuW4fe
5k/ocN7eKBkvDkuUPLizdrzzyG6DKiKQ02uMhARh7304dabkIRFHpfZ+twn4dGsOY0l+Y4AebkCv
3UH+TF+W3Rtj/myXvV6qcSUrbQzgwcrLsCjaCgXgBxvTEa95e1RNBnJRi6ikRZ63ZiTMzcnQImEs
Y1hAck//7hxL2YtU4N7SELJHDvaHzdOj3PIF/5P8E7wf+yshN5A3ypLMoDWMqYLNq7AkcC7vQyMx
sM/83geZaAEOTEfoSU1ckxLkJu9KkV84R6Ld/CamlCTwSppcrIElx0CxzLN2MEtwourfoiWLDDoO
8WXPW7x9Pub2oO2heinEuUo+tnNm1SiDjwcZekRdci+r7xUO2NbcruG4h+awePnBBRKwzfago6hd
ftZxVhUyY+e6BEpWgURPwgqyYdGiE/vNu46leZKTYcnVnoVDxCPzrJx+w88LND3aIDgUT4UZMbVZ
A9mlUe75sHaTw5r8VQlCsoXZntnft+SXF32txyM80JwHe/tWeq22d1F5n5OxFpvfnPZsJZe056rv
7d0n0GkSEM4vTmehWpY8TShUbwyasRPWHNRZIZM0nwi8dZvn/DTJ1c9ZzY2HH2vUjIO6Co8j9Gtu
nXtZMeOCNxEKemr2+goiv/zaRxdk3Uk7iAl8uAK4Jq5w6+7Z0PUrRozhWWNJbgfEC9KlZUn4IrRu
zOXbCdzoj1silgh3HSijULSuL+HGbFB3SV4So2FMMK3MW8OiOkt7DD/ObypCSAYKpL+tNTitN/rv
6oxZj/SJnjw2QRsPh1JwmR58pu5vYcGws+kEFZLTIQDktRofi+c3dRWfdQdVck1KLmTL3UC6p1oe
z00VSTQjDfxw6uSv6yYm2C08LX/43JaqxZvpKI4cg2oVK5XngGylwmOVOpsSKZ8Ul8xob6Qlr0qa
vM7EjPmmhksLe8wIlWeJIpwLRgI6aKpQWIME44RuHhm0WLkpZj7xfJwn1QbBPs7zjSHwv4AvF9C+
pH/hIvniffvSjc1RcZru/YXilT0HQUravd11ZZXplI/dY1RCjDzmAO4QOGNCebTD/agXQe6vaJv8
xcR9WUT/ShlfByz4L4GPTpwMdUwFyk7lLZq9CkHkrGudU3K8Ya/QGt3AUNWNz2M9qKSqOQ79FMAA
DxJ1bKufaJ1ZlvVBdynZf22hcQt1NwzzB513w0LNkLIHwiz5/qPveEXgNm8PFJUp/olcEpwWaZcD
IQvJp4fDJUeKZkj0kuSFH8I8WKSu72bx8dXHNiidpN88vcC/Sz734QxgZBzuTyJxR7iYrTToWG2W
LsoK/MZ6yfdGdpxDfG/RRaRpOPuiTrckXNkcEKRBO6plV2hOYeN7LdJff3Sgd1dt3LjFzzR2K0Li
CKrgLfZh5ZCnoEZmuwfEeMlrq5wc+6mno+xt3xyVaMfhUyinh6cw6WN+Akd1bfgVVGVsA8Jp45Mj
uv7T7loFB+IvREGdiBnz8Y5wkAjBJ4DnzwM93E0obGng70KqvAJs8VLKXKNxWY03FLVVvrJw+z0H
ITPxBaG9CIUDwahCm1sPyXT8mDhIRGo0YeD2x3J2IyvkE48l4NwKar6ldvcJ6nVv8ry3TTe5Ud+Q
G5BEDPb2yNYFq+Mnq8VZ3T3w2rtbDi8shgB5RpytXPkpuAGynTgZj8WMhkW2bX6ka2mRaqtQSndg
ewl11UY2eSPkBxePLoMYjJ414xX/KPt9N4Tc2QhPhi7RUY3JlfSqg7JAJm4zGW3ctQI3gZeHp0LZ
Gu403F/24DQvyZVyJKMrVxwjuRhvSrUKVi3g4EBKyg4GlqAAXxkx+85j2oWwwU8m0MStYuXSxozk
dUffZP5S3VvmWgljPFRqbZ9LcjxEvRYhpcsfW3ybgCsQmHTQ7yleAi2qmMHm1rL5iTRArrebpl+f
UlLTEufHccVR0a4g+PRzYE62hFlKnGPAdmqiq+YkOi01Fdn1iFAcvCBoO7QsUYZT0beZ+ZmsWWDo
DP34ayYvotKu2oYgMpD3BR8aSzE1cs6p+edB/7dWrmWCzidRG7kYnPWKf4dMRN7lqIXsVWDfmI9D
WGUKMLlJHU+zmvQnFmR0z335oAUE+0ENtDLmy06XRby8eT7zOEVjeCitaQVnvXuLIBTKekRfuV0e
fD1z1g6c2QwUGCVmxe47/7hv/IDpbEyveslXuV+Wf0erfhafIMwFWwMwwFoK4/JGYnCTioIjPuUF
ewOPkhh2uPFrz4oYa027ARnQhYUi+hJ5CMp0AiKu/XpvAT1atXBVtM65bcGl+7gEnz5ha810BUrv
WgGsmHePJpAu4vgFa/k90VwzB5t7KrQ3aKBEuyF835veglkOcHOgP1gewN3RyLzBnZGrTgMNz9lX
m4uFwVVoIGs4puqA4x87zlxfJXSZhsFmk7qcbD5/fzCbmPS+NA1YTO09TY8DuYEZS2t8mTpeW+nM
aB6rB6CIGWm1RegNCyTXe3ebFC1hGHR6l4rqISfu355YxzO6+MPXkBtdIqef9RLc/LXOUjlkjniK
w3RA7dDSV54MdPvphxvIUR0q3KkWxSnxNAEcEI8kF3ugoiKlCWFmOzyX4JFbINszEJXGRllYj3eb
+iug1kBdlHzIPEAi7hlT8R+r17sHVLAz++LntVtI+PpSeUuTb+da0rn5oCe7zrui/omEFGyHte81
Ovt0i1ioQEMzVtTUQJNi02kCekQ0sBtDokW6/3QKQxPV9dT+z+lvqJ85jcM8cUs71BwuZuX8fPHP
Tx3G2VZmAiziMzsV+mApvS7+Dkj7F/VdiY7dhggPoMw0rFsCyEv6rcu4E+PK00HIJS22i4KvmIgn
zqA5gpiow9mHsLvu9D5QQSZYezbWpzFH2vteoY8phyAJywBJMqQG4B23yamqAQqNU9aXZ+kwEdLi
IjmWk3St4rk4YF18CvfAwPVOF2e5hH7TO0lEi1rjnJ7dc2tKnXnWNNL6jofdz7m6jz+JiSFsLMMg
c4aNqy5nE/RQ6LWjpZgGpXPjTAew53C7gKFVJjurFvCLxwCjh8rX4LsgyC3gxWfLI8672DbDJkon
ywM/Vum+nVi/UmFkjqwBO7qy5h26bbbib6AnTss56rVRQCgFapmRotwr3BxSh7fXp6oCozKMRwdy
izyjavyDVenufvLth/bN2Uxl+C2cWXV+yWXtwK5iSTRDPtt48ZaTNtB7eaW60KwbfoTUA88N7W65
v6F7k0GL9gn6f96quFY+AVoewrivEveKcQwQ+lImuewFWHmjQ4CcUzO12dXJ/0+cAN9b9V288AX6
GN1hMKaOnlasEo1ghYMxPL5XTTcqVVIggMvejzOhsMUN9KqrjWpwOP9ZLgicRdRDPXVXitmt+fJW
yjgrEEN2f2IbEGREH1pCH8JMw/PrSWWw0r+kaTLqctF2dAY4fq9NiYdnEW0MKh7O6TzKGjd8Wlnp
zWOqEctWfH09W7GAApKkVfaTgIoGoHZvCXkWY5xzFQiajWYvIdDGRsaWclGi14rQwKwZs/Xzv67k
FCKeWAVqS2uEo2qaqm6HMjiv8S/3wNAFaTmjkryqhv9yrXu7LvW+QocijSVdzVZDok+e/Bbro94v
b39zSZ3MYFjzKoujpuXZeNPlCzKTw9B6gSNEN3GaawPnM6UM+ZoaJff4loxgyh3K39ncLZwjXUMs
699m2SHNPNkHinandaeNp3LwJZk0gz0bhQk2V81HhTDm4KwCB/9G82HqU5YBkTQ1GdCQ/QYFrtl1
Nj/uOTAOLegcq/Ql6GdQWmrt6DjxKzz5bp+WQwK1e7/7o0XixhkcWuXXMGnnPN8nxFHT9wlk7Iuf
5ox9u8ILHjD6ociC660jQITw0N0uUYBFqYRUIjJWBFzPFjBja23KMOLaJOqzAyGZzTdP/kbSbgWn
RVBMmkc9ECWe1uEGjo/HW6b8yC0A1Y9NdWoaW+VTMtfGGgrpyzxGC5y5sCSJDuLMt1sGMt75rV7H
mqNbEtEWEjf2ky/0+h02TLXsYUnWqyRW5ZRyJu3cngpSdHiTtmd17hQBDuL08Xw+N9DSJQDaYF5j
EL9yF7hRvXNt3KsIuxZ+HnDYKbPdc34v8OZpRjxjuMY7GQPO4bEzogf65CAES+wdBZwVAq8OUIZn
wr0T8FeJflYnLjxNxatELkcbJ3rvLgHHFLuAqBMK47fssqdpqxDWQIY7XxuyhWKC22Ao9HNS5MGI
N6jzZ1MSmiPJvf1HW/R2/Cd0WHU4o8wIc7zP/khPIbltHn36c7TglY4M+D2NU1ovGn0B4t2jOJiI
dvXxLPTVQIOvAp6axVabRQ0mLI+0BvFUdXG1KEM9dhb50yKiK09eHIQuihU+3MLAJr2SoixkfcA3
AJUZsyZljReI1a10jxIQAkZ5Zux3V5aVnCDArcFcr0iBs2Tc0GtQdf1gkJumUyDnfzunD3sUP96I
VTwTZ0j2fDg7MydTPn4W0cNuU/yHvMTO8KfUTTBKCF5wxpwBySHQ5oUdPSpRveS1HhUAaqgOw9Xm
4NYdAHRMa/ogMnItjp1WIMW6JdFZeOOVoNqJGkX/ru55R+c7ClKEzmGLZN9fnr3eqY7VPKTuND37
UHsp8YDM1+qfknqxoKcGGbNmFlf6Wz+MaObdGZB92LWFZ09FGBtR9g0s0AiCcfvrOeoN8Lz35asd
jJCV/6EgJv3Ip1en8kEUNKBIYk/1S+SWR9pD0zRciJlhPemqaKmSHiJVyTQNVM2e8lHHche4a8RF
b/8U5LtbOc86WidsvZFDiUcKRD6Gpak8ag8ZKZ/+ZMXBf6FBw6woG9+Uo2t+xiMWj1Fcj5zV/cL4
6xUWKgqMVwKoV6B30PpSsm+h0U7R6PjzViBETLzSM/BmIfWL3t8K5lBt1/QcoARoAb/X3nu+ynU+
5TN8XtOFMY4c+Mc6fbIufeg12jkZJYXmU88BG8v60WEBG9mIhSOxYRYhJUjs54PAYEX0SvUp8Y30
H//mQX9NlAO7sTfo36zq9OQJgBgpSh97MLpjoHIA7+jOYQnVqyvZejHdQF+MaWiUvcozL7CmJZVo
lm62fNTvc7YWYUWHLmDfptRPFxna3YZeC3WspMGyxoja/QEoofNpgia1J5gEgmsCfRSVZ/keTJDQ
4XrqklDPWYDaYeWbnUNjaURMiwAc9nW7pI8RqNvDUeuq0QlREwThv6RNxWp2ZTyo2c02QbLG9cyc
OB2+q3KI0B4Zox/Z2ilSvybpRUdLNWIiTJZo7GQUU13I/QdgCbeObLQgSX5+7zlssmO0korM0mfs
L7bBcL2smQzYeI96RZGsZkQRK/L2TovyrOQUyOfS/YS19EIZ9Ym1tWfTaypx8ZrIgghClNVJIqxS
g8o8CCZb6bnBLE6nQ99Gj6RC6Yv0JvAE0peHVPli8YvrAySPLAIjOcOfk310U9zc4/4fRJaXP0Pc
/TuvBjj5mAxIO2VIMV5mmpT1a/OXQ5s9B18aiQrCQr6P6lHHc+hw/i0PVIeJPc3EbnBrSAmBGvSS
jM7Rc4bpZjHPpJ7W/h5V86qdWL/tqu6Ng2jQXrUp9EiiGJb/WFHcoBsJ+C1pX3f9/+7BdVz9LJnN
7ojaxMRMbTMM6gJlyLCg1jw/Aab+bJsO1o7TjIqltYtXUdOibqhOhMbUhMj4iSF1Q8zHSfxm3r4Q
WImU6NpZruwwvVr7hv6Y3sCs6cs8x850JHripX+Xnh7vA/UqnIp7BDeWXsKf4hUieMI0FGHglzdP
eeJOkwCaX2UFYcLtvrp2dzuznV5kuUVawu8iQao5KS/MywBxUfMAo/BvBwKPgy7/cRz2iT2vVMpc
JixDZL8IU31NWpWbSlCp4E8EMHd5kSlR9Kz1FFtp9TLS1RTKByIZtZcDQErjmJ9I+QD1JM5gBgdA
2EbVYDo1hoDukNAkBj/Qp5Wj2C6+2xzfDDSCl2bTEozhjro9aowFdXTE21X30Wvzr51iz0F+zfNH
yJmMvWETABWd0DAqUR2N8dUEfdDqLXwU6Xp1WCLh5tzK6NuaYbnSZoWfaT58LEb3P0nN91PlSuNF
Pbe4JH+AaBHvoKP2F+OcY9wv/EshjIEdluxsaAdgDvBjznJu1rs70flrCzkt+Sg1YUaG+GFQQCoG
xoCfXsFQ8Q2PbSOGq0RLxmuoIGHYCzzO72k37h9ZNS+39n+QJWScdscHLkWIvKxAHfyfPoTSpFnL
J2JvsRTTysBbam7A4vJyfmQbIVJr+wct0638jrS8bV8sjSZwGu7kYruSSu55d0JQb/W/VHVe4rg9
7HCSQKTAmU66A6cyu3qqTW35j4SKy9ecQjJPNwgMMIwKmTYCE07F7oEkPrYSHC/GXdHy3E9LglAy
7aca7QxIFhbmiK/pnXBzSjsO+f/mQLYj0/GgQcKR11J8YT6MbIXkJU0fsEFu7VQPfXMq+wyRnJml
mTfG603ysxsNBFn4a1264kgsEL+OCN8XN/mh2vZO2NT8MQEgxakfD6Hj3yk05CtFtcnTqTrV4Jki
qkStltIxq4DONfsXy6W3vNggdZ3sRE0FWcI66vu6CLLts3I35W76g+/bJln3bG9sbk7BDdplXBuy
aFSQs1YZkB/60pmhU3GpmmZeeYkRBSNkbUz1Y5fZ/7HYBIoUEbfWjq2T5JKQOkBjXOavzWqSlSRt
W9cvpdzBwGa+pXVYZ7R0bx9yzIdoK56Tw63g/qKLstUjEP2s/73T1lYSVfIZUGRFyTR330GfLNmC
d2eCFnAru5Ztp32Y5QjJfRasbnQZ/bd4O6jUAPAj7Utn4D8qftZ5RsOukFHafjqhfVJwFbw2QDz/
MNHqlGPy5Cd9DlnSseMUyEs74fXZwtaELCw+6RrzFeOLHt9PyIMFvh33JN/Lq+fGMQ1TuWLE1UEP
noO+uJQkBVbcwU2MezZzxmWWiFoinAlkoQ2K0NZllMeYHoV3EvUX0OdRwG/fmfaVUkGi50KOuOZT
WUmaiEJw9Jrbra/dGkh7coTNuOnC6PvLMifg3qDNwxuFI6LRurOusw4JLO5Jy9ApgHqnBFNxLK7z
wep2E8g4k8A9rlxNI1YZc6i/LY334mctfg67eJlOilpQRuBcgLf/FGfPP48McMjEVX38fHXGyrTM
NWpwmmwgPMtnBBpqOnZjXtA2XeAAuJiySyLTAU+mHIBF731MhOpIKvNFxeh6Bq9HMkdW6uH+N6PR
Iuw+J5/APeedlB99XxA5S6HduSdJ7Wf/Pgmv4kIIkUDJhcnxs21M8t//j0yjsjpdc7FNOe6dFlRZ
nS3IiD60KXETJMxRRyTjWrfmiyTzoquVCEJlxNmprr0u72xfscgrI54kvO+NtHCBRougiwys5reZ
Wep64Eu9S0+eegT5E596vyMfhHKaZ5jmLprwH2dpzMGdMLwlJjw6GzO8peoBO6BiLbgRQ0zOtPzm
Ear+k8oJEVDeH36Zr28egi4UJ2c0mD72jvF5vRS3O3eUcO2Omf9A3u0wsDGwI7bVxUP8XfNhCNKT
MjGxEKiToW1UDybWuQvZucI+546eEICaVuR8pV/sTufKHGdOQWdWyi+fCE89p8uWnovU+U7DhoGZ
0C5ZnCYoi2hl97/TA3yb67dZeq9pJhtFFlZY6z+aYSyIGGYMDXUvNJu6UldVj3mDOUN0ace+0aHL
GT0qAUZncEc2YRZ5AVb+XeleXPXT6XL3QXxIdT3qEz7rOwVzGmSVfPZ0hE2aPpi8QeoAfN7UCqJN
lqXs0fJnESCoTHYMC9k1USbx+en7o1tjlgMYwH1Nzep4ncVsTBL8lSkoyOQNqoLwuq4zVcy7veIx
8aMCXkLgQY4C0hT0k39x4IjH12bOMlUJeN5lyDepsAk+VLEiMDX5bMQNATWjcYHpgxh17MEgiw5c
9Mz6VZYlLAGMcJKG03+AOZ+h/HiUHDz6lR85GYt00LE83gKOLFDDyYwwVT2YJnw1nZq0FB1C80QX
ikhIXXH0miLsXB3LODzdc2nnaQ8qQOI59zdjlnUBxcvWJcM+UWPsj9yLK51S6BMsZTY42ULdp6Rh
p4goVAsv7D928HnupFx2LuIbE8gzW7Z82mH8eQJG1qeeSXN/w5vUTjOO2YRklqWOCS9Zqb8a+qFh
YFxFbjOoxgcY42d2LEWYm3wdreQSYSsRdF3vphkXOQzFT10WhGRrXU5SI35eZNAVTxWDtmHIATL8
+5WEvU9pMZuILRSRhp8G643wz7WEruvvUxmS2ENf0dhmiWsePxwwdgGwGD1DAziPYLlTo9bPyFvy
o+2z+gAj7Hvu8SXPoLTKG8usQ3GEIGyMGUpOZF9uF1Ob6wvY6oCEvzzrGzhijzpoDKdUfdLoCpXR
h/q2YnPzYQHgoa0U6Hb93uYmrlalhCjJ6JzuXxGWdn1SKFfBouw8TDMDgV6ZRCZpdTT4H8kSFLDH
GCiTCyVTuyYIsmUYbdbJ8owhA4Yw4iRc9/aCpsPQ1AmnOLol1qYf8sVFBWI4d8O8syT3aTbecAMy
aJLlrZJABQGT2cLJal0DrprTfy/cgkR3mh7o6biYBfDfNKzSETsgI5c1poHiMTFRQc/pIUrzCA5f
sipMkUbpw8QfcVE7c0DYqgVI3bd+GNdfg2kZWl43FSsgYKzjwinhy2wN0T7IHyofJeh3caSwZlwq
95upLnTY4W/PHgVyzpA/uZH3VdsbxAbhYe1tK+IK/fxF81QtOOuS6Pofvu4ZzJaHw/N6t11U2ssl
/veUj2rEMoOP9bWpS0oJ+Qx54WBktwVx3sxpzop1GM+VnkIG+N5A8X10ymf2Fb8cPjIKfLJcPhvj
ES53WWO1OAi1OTP8bPQA7DS+UMg0Y1+jm37SCccyd7T3gABjilS3Xzg+GM3B3kW1tobvIMK+BDQg
NEnz4xqMOlOThvI+DgT0MZaDAUCZTwiKV4MSMvZ3k6Q9LT0lbj0xnrRvZ00RInQljmx2eLGfyU4v
hpo2xeI4MqzMGWbeKsbv8nh93sv6CKSM1oTYaPySlh3I8p+stfYoiPyst9ZMImr0p7Zrh03Y96bi
SWcmdpZ4VVABNa+xQll7tYr+BFDdJKSBL5Kg+2jeXD9fowjdes7NM+tNgfg2dfcn0p6JTu/vAS6P
ss1I2qggfva5srAbncJB7rfUj4QEwVIqRO7eL2LsTl/pRvY40duv6Ow5ypWCqh9LO+jmUUZWMQmT
hunTs40nlUsSH/Fsy7hDoLzJ9k40n+RYgC/cnaQKoGSOLR++oo6CyFHjyVK9nmyx8ZVV31epi0HD
hJwJ5lR/Gr5gdGpu3mMTeLANrbc7pXZ8W8q4d9BerYpzRIdzwIwhxOw1U5WswKd5w8JNK5WdrSup
45P+CAw6mh5DpsA26M8VGG3vtS2aGYOd27bJCJBnVPXNEK+2ZSDBPKT68RKxXGV64AA0tNii3CET
1nMSl+7AuJhylY0khNnyD4qiUVnq3f22jlQUGzawgAhP9Cl8yGSBc8LiIV7g1ERZpXzAUoP5qCyS
bjLcmcket5G8+8RPhiAQGjoxlzXhP1PLNh3ITCqrAChPHKrjy6fvTjD+34DekcK0KN05hoVhT4Zi
UnPLVyK9G65PZXt8OkTStukampkyZk+g9vhZ4UceA7+92eYtz4gTKtX3Ge5h8R8sbizkMbfnS1uf
SqyRVh2clNCACuHpqQg1EFLrYJByc9mwaRLhUNiS+96fZp+Wzr+YExyAea4JFr5dkTEpb88f6Aza
VbtSCXr2HKb5FD+m4DyI9AvAIjHiPHQskg2u2QJOjHQzTSeXfDlANSkXQKl8X97V98cHLIId0HXc
dmrzgFgx9uT8Ma+Y5ut2O+byKZm0+cXs3VMVJg4cuZML2Y+APRCcIgyJa6vhkZMSRq66x8LGDXeE
0EdmeJlpwI57hrmZ9C1v9Km3+LrY+2ylXUvfxgelHQycs8XK1IEcyKWoHYDNkMNJT9UnqEJsoS9e
KtJZn3d87+7Js1JAInMEOH2wJAYOCZwTUNcbD36oSGw+m73laQikga0yhmnDQtmobWG6xxBd588w
JYwNEn2/mo9yrlI/DZg64RDgmuyTitm1h2z1iLGt1NTvJcWTHTFRgHbAOYRbnWwO3Bom2Kqb2sLI
YuQc4RCOHMeIqbevsq+PYKO6slzW9dj0Nn1TLT37O45DhFBPeAjYbia7Kua/9E9IIU7gahyKVXKw
KxtlyypNY95BHmfePTfgbUxzYbisXDRmXlJ3ny7Tl8iENz6mazBbc5SaaWU8+X2ByOf6/2brRe5L
+B7Irc+vEQ/wgGluIAuXWlpjJJYve3VOnfRMUEKsNXIHZRyVMVRXQWEohNWMIp/HJL9nOeGIqE5y
tX4YwzHCCc6U0LIz9yqHckNR0+79TNpltz8TEvVsMDfYz5nD6BWrf724zPSIZjh/6ewTgru0tR9g
BWZkYPzQJfB/aXDKIW0eq/zpUeGNpD0XY7QvInGU/JALmzw7LA10FIgic9OKmfGhbLijTN47ONzK
K1vCixxqPY9miCv7THld01axkoZCzaDD10D42QlBcimmI+l3U4YbRGoJD4iboHtKI7vc3Ul4nwBS
+OzS/NJ6q/v3/qfz5BVBBkI662JfLybtOYnZlavS64vv6BI7etQ8R0kn0xjJDq0LTVOYKU7ygARs
JNG3mk/Vn7E9/6swyox/zAkJP0lUd1Up/Gm3yKz3qjFOBZFQBviks5lvutD4w7vhoAQup681t6bN
YZ9w6VXbmcrwbSKSN/2ufZG2iCpiMPl7SxpAxRuAPEl3VIQJqrhYyBjYoO0X3494DstPcx7TduSi
VIcQIyXU7IA4lbCU04Slvb0xknJiV3SdDCRw4DBvbmUK6seyZICy6wqjO92Xhts3XAWoL+VJIrJb
u0XxD/fyKFEoc+DbO4PQoZP6QLGQDEFW66aAhAWlE/efqSKquqenQW2B6dUUiIImeqxXmBbasUQK
o3yfh0p1i8hKGaF1ajoBpaI9hdJ8KiSJBG4s2JDBIHrWkIYct2ls/unieNmbKmbIAwzOI3VxE7FE
4TZ/+16pXpRs1B7rFagsDJsvPBnDMGjAt9we3ZWX0x8nr4g+TQQXxpwMcVJs8/F2m+1tk/J5jGDo
DbrndgZNOnl475IEwqjikp1k9IPP7yiY8y6NQzCJV2vIIJtrXyngBsrP/1DfHolbvGIhuhtpa5Gn
mS8GcDd6xNGrWEY+T0eaCtH7l5QXzgRrQJuKi+clGG/Eg4Pb3+WzYMB2BG5rT4UoAWyVAuE/mdN/
KVwn9cNzR5q0GT5jBHWCTo8TWP80xtxeo04iscaXWLd1q9oDXrR/1M6UB5c4BlW71ESiHYcy+sVA
7prjeMaftudo7BINeQG8lLcpFMzNPQ5XbpSKG6vVK8APVAmVBJEE539WKUXRNisCiUXP3/F6epjv
YEsET2+pDxvdAPwnoxZN/NidTbsWXj4BhnVtIfdWr43R0s4EGi3QRsG04W9L5GtmAyxvA1Lgk5Uo
81w7Yg6lAZxMFfb831/6jGd0Hdtp7eaWlHMAZflL0WDw8SKEUpDabW2hLpTuIasppl9fuhG+Dibf
5VhRHWYaqC9veYsZUWzIWaARpNmjq4C5gziWW193AXxaapHRoGSiMz5uq9an7h2PcHfFhru/ITkC
H1P7oxxQsithYweWxJpnqcZlTWkEF3GfeCNsW3PqnCNeA8Ie2IWBlTERcHM4UAENzTq87K8Rqwgj
heJ+/rW2Qb9q8EGhxG+sRm8KTBKg9zaRxrhlLphZw2hqtF9I0ZLc1p77hDxJl9aK3Eu9jiH/hlMh
XI86tFYm2y/kdkqMJSA4rCLh4CJtkPu4DHjj+df7ANixBtpryc0kMIxFfcNllQzKKO2/yny7owi1
gdn15uPJH3wi5hUVYpQIE8DSGU3F142hHgPc6XiRBmsD3GFiAGT+dKK52sXhgSnQihcNZxzYXr67
RxvDWKNquckfbgBPkfMWQegQkbT3BN93gB4fy8Z55O+xSxnDqdZzT8pSXBPf6Lgq5toavL7i3CNS
OEr7Qzel1ngTNutRctno3+EE7eVJumZ1u1joA6Y3XgkMdTGqVtm1d+bZmoxOIRbEEWRpYUy+jUJg
IHtOFNB+ZYmqF80LGebfpm4C/UW+/GtdIFKLLAQZgAmTz6rugtIof6g3wUjNx4qE/vGj+e+pmsyP
WczK14DTxulII37dIpmQTM5tMyx31pvP5B8s7MBZl70mUM6fqIz7xeBsyprrpLEc9pcDtSV2YKoA
cSBJGY0LvK5gMfX+YFHcMBYaVrCv64Zzi3Ad5h4QfKvFYkPC+i+Tx8+mOAwEubFH6c9yX4HJ7y2j
LJkwwQeXsuwvkWUGjIL+gCRcEQdNyQLP4YY2aMhA12g3x3zoK8p4oMPV0mDtzk3PgbJbONem5kFY
XURwRkjjx2kWQ/pOmYFtigARS+Tl53ThpOqRKIvxrl97/DVNH3iANZlV3XanpqwfI4Y5weBu+VvZ
cmFpR9cN8oTK6VOy2yIzEyPxdZhQ220XiwMj3xS0NzftFal3rSyHRgYP7uLDrlmst5QCiLEJq5M8
lKfwJOIm5v1G+kJdz0mnvq69KOer9xG5k0ijzO0VxdKjXLCPH3spPNrCbi0HNt1A9BKtDEwCy+92
zZw7T5/Tnrm3T2WnU2pRKlfu/IDqnEKEOoPkcCLPXwtwjn5YQYpjZFjNoR1r0fSt0WL4+BulLAf2
38fS4ksZkJiQZIr1V6eWobi8yDuWX0fpGQDkVMXbLFPctp7VLcRNTYPF6w+2K8QpK2SdEnFV+SKb
UkZ+DVRVCk+A91/4oyeXbXa8AUdxD/4rN9DWLmjljXSD64+j/w3A7+VIqXIphwtJBdaORkGsySWY
5StIlGmB0TBYR+FxQpPFc6UfGM2c81swpHb1aVpgxBLthE1JKDoBfpElA2OB0CA0Bz2Jie6jLfe6
R+u0Y0yATfx03NKSo1qVie9KTjCkZd1qbL0gyhNTFhdyctXWsOzD0p6u9yF+0jLnltTBwfnjJD/j
U1/CZjkXtwzZofkwt4Lg8UP3pCPVxU0qFwSSON6n8tLFHCdGpUOBb+ttdxQdrDJt6ogFwz4F27nw
+RCOA/BK+Hujs3CC7dvpK/9su4aWVWkvacpTypzmNWdq7fkXQ1wB3EGw2GcHZlPzCnqzIbAYJbGX
3IghUkt6FUYhm0auPTNPNSHxIzdl3h/AJPksFc9kc8OnMIGsfDn5mNtZW+WFnjq4/QLBbr0ni7oq
IiCjIf5ucLhpqTyTsLf5cska65JWQlRt4MRg2bv0DvPYt8iIjJHGNnmep0r2FZvYAl5vAUwxR/tb
FZ2csSfTOyHYeQo28zSJ9VvM0dh2iP2YPfOgOxGwIH93fCSWZaihuYTtObjNT1RnWnD3qdrqenKj
dfxS9PlpCxx4jDK0goKvLuSjzHpDyYWpvPJaFN/u3anmyiitx6wZ4qmwwe2s1Gv++hdjOXJlcXrV
qGuBTnQH9+/kd0JvAaNjiZAoetiuE9Gy5tHMk4jG9WMxM0Fe771Aq/nbrDr8DKGr2rLjxesuMoaA
+d2LNb7cDS/Lpoah7WbV+mkGXd7h1dVvcdz45irAdcKgb8LhkJhFGKhEpkulPwZsSNZFOuzenhLA
H5sYQfGXY2AUOMlTQAqHDiwMqSMyDkXoRlw8ojmPDcmwVVwojEjt/EYGrnRO9rn85TGJbgyLZ2AD
p9b+kKUKDPMKLUFR19nTM2/GcVT7Q7MH+21DfYrvF9tKoeauzOBJ8NgAkc/dk5dhSaVek08Z4W+P
Z6aNrAK8O0k/OlZDKJeRu8gTMeK0AkcHKAk8qW/sN//cgQiWOxz3IFneefpF2ZHZ+6xG1LwHJ+Yu
1R1IdmvZTNY8TczLp4cHQLohnLKH/S45jsFk7Yb+L3hk9cEgZKCTLBDiYfc4q6JZN/VgAyXmdjik
0/sBybFSdQoQaolrTstC1kPEJE0yLO9pUOlRH+NVDc7/6JOp8fm9CkBgwht3ou3Lab8PANEBEZVE
MXdKXjHxeyUy9nYmYY+5KINGgbprv6kPdEwQhXesB+9bbfeTebJOLomIcl+4aoaJ1EHsf+tocD79
hX+7RhCnp3SBIDN4+V2ANd6fUpk6Cb2TKCpi+fABCqnRVng8Qf3UDRpj+vdmvQsOt+wdjY/k/VN3
Mq41sZS4UfTmXbBxyJuRkz3CzkpuuX66FCDH+fRxdkX65fusdGejSaz5LaP/D4zcTo1pTOVIZ+r2
DTcjksInfS8yilJGDtqrCjO+OLWmm42m0CWc+89C0YqoVaeYNZ9AF+sfqYW3IEF4j7Vr3MF9ou+3
inrpt+jnV6+FYDuj4//TR62yo20+vTBgLSa897RMv5/mN0SZlF4gaG4u2PJTiNHraPkoXhu8VxyU
Mcoyhck1BCWR8x/HnNlUCkvzwXyrjEhzFUI9gv/RAGagC78IgKdPqT7aLrAkid5Ej2pS+mMGow/D
Gt4RZEJYF3ikZn/voanYuhT55wSKHXz/aFZRNFPJvBJ07VZ8Dsu64PWzPDoprgZlSi1CFZUiNkgR
sOwPWLbPi+37b1kNXuT8MQu+IHbKZemgU2sGXMdzAAYmZa0b0fLlhTidTkMLTqeyElFdFNpPs/gG
/lUtwsLjlTRtr8wgCJ9/tukZ5k1nta8hdMKkM6P8DF7Ddzw/QTNW0t8x1KHlewD6r/ruZE6l57Cc
XUZG2dfuSv0ahYLh/x2wFvGqxytplkHVVR3x/CvKEmUcPmaic0Mq355tO2HY1JZ8DYvhtdWUrU60
g26W2TIYJUX1A+OvDMyhSmhzyVyHXn9v4t3FsFwikz9Fd1z7R38f1IX/Dyysieti6KCK5grELryq
l6aeAlTNmka3+BPNGp4OHr3OHS9aX/JX7ovEuRJ+R0jU4coeHlN03EhKPv/DjAoebh6qvJ5NZWVU
NrreAe1rU0E9rWd/LwKgfynlWo3z788hRFq/8BqCviwDVUN19r8SY35gdQvEPZm12sEZtLfun3Io
E1V2vPbmwsOnVnaZneXmP92UWMeE7O6uHnLGUKynueWB9aRtjxgPN0dwxR/tWgPF5RjimEVrgGKM
K+ZEfM8EqdLVxi8hKrLFSrOyPUekCQQlrDSh5/8AGg1XBiVu6lT4z80+r1P2cyLHv3A35wjqEcJI
YXE1TsWxcT6aY6zrHncpCYmlQB/Q17vJM9jJYvoK5ZKUTSGbUfuNYBMtvkD/Am318zx5ZhWhx1aq
IaNKDW9FVXbOzSDGKGFgl9jKO3jVdXyBSE7wL+3GLCFDcNqhqkz2hEu841Zpeh+vVgzo81Li+jM9
oHulSxy4kctqfSV3MmSWN9sRabFheKJOxV/tCFcu+2IcFP9vjMZF35wmzM20VzSvLgN+b4LHkas5
WcIjE9DIP/CrctenRZgCZ/igZyZhaiqVHu0y2dYCmwzWKCBAMYAfDLs8FO7PDeo1C54VcvHGIGhQ
l0yEweR841PQrYXho8AQfXuthwVpatLp29jfoE6PygTxOXZtiy/kYoq6NIept7qlgQa+XaacM4FY
Dv9FW3v37m7zaDZJikwoDibIuo7LWATSopf41SUClaexbeNstSyvhqfGl48ccZh97TvLs01VVC7O
zd2aaJe/6nwHZCH/D+Xwux0yOjqre7qU5UwUkI9y0+Ckvm28m3D0KnE6fswLh50GwntyAVgWNGxG
BoFZ7DbFPq8AhYaK23hswJCXRMpCB485ZkZ5pgFng5cm7ojuIAKsjRLQaByGacXpCZYVRR99THB+
BwV6il+EUvulxPQOFjiDXcjLYIfJdT5AvHJlvOlKn/RiHOkeg1ZwS8byNCt8yy/UfIBT4aIHUJLl
ubrcn+9sy85BbQJO9AyyRj0fRyMlov6nJ8vgfk3OKqyJcva9rtdowDxb5yMx4K/FuQOMr6prC5xi
aFWXMLPpj8gazeG7KqoFp+e77ZObRUubcMYsNFIE94uHuziSwW4PGK9FR2ubb76sLBnd2YP5DZlL
UYUmmistgs9U2LgddcQbP82pDmZhVCGNe9DXHKJGwTCTGdI163pG5JDIyfiNEghHC18MOnXSt5Tl
F93a543iRZsrJWso04X7+nsJSfW4V5vQL1AWiheZJwcJolajbnNX/LJRrbs9dDHbh5yybyJYSs++
wCrFK1vvAvC4J5UMF2c5xhojgCfsRrfyrrn7eMIGq/1unaPbCMssy6mFIBfhUa1ZV8KPeP5Vy8PN
hDXIOiKf7Th8I7pD88L/Ja7wsp3t4gyN9er3wqLtqAcqCLcCxCT6JsUpLyLbG+ckgnjMetudmcbO
QC9kFUUcguWX5Yq66/efJDPA2ZzOLkpeqvP9O98ljxpHdWD+RVVrXovJ5XVNRaXsPNrBiYjLI5AA
sLWTlnYAzQFZ9YR+tnih3To1Nkyabkzp/mhrHXSJt7WYbTgO5IggN7JSWNxWuuplZfleM850d3d1
q+63wp8cOpFGBpNIOOBk+GyrP4Frf8VYZyhEd/aRTudLgbHTe3hMrl8h/dO3KWRDzZw39SfHEdki
Iiao4M3K/GHyjJy7qs2atAhn76X+nGFfrjtjGjcEwrVEyJ5N5U9a2KCTqhRa2hTzbqa1Jp//LgGV
7xsx59222HCNDMO5C2YsafhV7jc2/ZGRbZuZ+uwYQyHw1WuB2YZtUpLzM2slDKtX7P/viVTb1Fgb
ve/5lWEyXZRqLEP3k+qzBQwBHV4oKf/FGSEYRLdtxX4LzqPt8JGGP06fP0MEWELJmdVaPubzM49t
vR3mu+JiOVygZWOuEMAl/+/oOUxQoJ4ypgsbKVokwUftU06szamP3FF2WgNSNRJG4aWN3AiMHpyP
FChQhcXzY2N8PB6+MuyZiydiG5tlMaVthwR6Fq+j2i+Pv8hMj2Fl6cOXRCYGUYY3QT6acVwXy1Sf
3+xANmFyrImCWHiyldXqCsE2cOktReHCB1sbIOfVW2KNPV8Srz/wd4OOgwHj+wFYoo7twD2T3XJh
tDjfWfsBbFd+jq4jdqBsK2+6fXsAIeJFTj7SaoVQcuBbQVUhv7dVGOluvY5RdRS37n6EOAVOrNNU
AgEosoLVUNeeJlsecjSBnS4NhRi04ml3pymOk0jntX/UU0JIFY6aEGzyMOWgDn3yccj1rZlKnDCw
anMcn07IOn4CpyA9TU48SEzl2hf91fpQjFUkuJVMrYA5WWKrHQnx2aLWTObSqvGLAmvTgAQprpC1
x9DKhafvF1jGP8iE6SjWcQZYudm4aJTg6Sl7YMZfOj5NDKuSnmbNLNZTPzaeAsjwSw6guj4Fp5tL
RFc2/EGt5uPYtwrjM9FvROLlkHSxBa4ZCvHZYw6B5w5/FojwKnQH7bTBn8RrNbu28r7j7LXrai6L
rTy7rA81t7NETxSPpdRtSyjCvkyqi+5ZKLxOH3HHRQkuGY/qEftExhFl6B23evNVvmCUt4XKIJaN
YOFGvj4MtlpVrQLgDJo5dWJOVgsgYqvy0Lh2pxXURpOg0oC7+whIm+YDKCtu2TFP5HauNQ5dyJVL
jfoj5yvRNHCoOA7oSruX8KIaPWHGWskloH3W2er6ETUbRQJghOX/0s24tXoRyhjHFV5FmcOMAkz7
Zdy8z/5GbhFgxYe6FTBmZyvJgiWK5yQCoXhk+f4kxIRBECeeOevBsXEAPeFY0PNfw7fRtYvtlswF
1YziSJxlb9EVeOiZXrN7hpFSrN6NUhZojlHIgFo9MF5ZfNBBVNnxNKbTErWcXRjfs5a+9uYkVlX5
rILV9M01i3LcWtzwkFaF6m0HIzoM0Cb+pEKRzbEkBNXUsnZvBQLr8fHPoo2oFynaLetj1ZTvJ24L
Ho21kC2WYSCHDGyqjzytV1byjHbe8LLFAb2Ql4Tm8ffHO/NUjF4U7SddD6EprbW6UTAR/0NnWIhQ
pzj+UxMFkY6UZVBIPF72rmzuZq7pYRPn65QKrPPYmktNHcELiSFCSEyMtiXWEBFE056rUtt4kC/P
yenV4dOJ3a5I/0eaPOiJDJ68PI2NeZxDOsw+JEpglb80DmuGZ0yXUwXhk7/D+la7gLLYdlkgnOdb
lA7A4pFOSfSvUH2mwMiA1dOkKk7rTfV++izNAJfNy1qooWIXCqOXQP/9G4VjTDUUtesFBeseA2W1
GhNldJvGsWHAEunTP99xyU+q12Rp8hRKHgigZjpN8Ph4OXjVIzO9W1zdOMKWiiOHrpo8S2E4MXP4
yWJ6leT7mfjYhH5KgvcMuMrYsIjnRQ11HrClgnvlia4OoCSJDPrH639uRQmgYaAHv/m0zNWk1Jzy
kqZVd/8IkoU/9PyL52RhMHAqGvlc9rLipnEmGhBZaYAcO9JauTQAAieqRhek+9jJ4x2jy+l6OnxT
ofP1+avZjKgPoA8xzTn4cUBE4i8KzeKi68tRe2oVFKB/Crfo7lv5dg3aKUy0GGMXkn6cq4mBqCJF
aYbEycIm6ulD4jDxv/SxK2nvtlJDnXGfhXIXsXkL802kSAVMisp8ujM+g/RL2Sz5Dq4ZJhwa75NC
ka2IbRSCU6ZC35AKH5gDnw+d7OG46jSlSmlBhYqti1+0LhGefjss/xhHhgDw+rwgWro2r8V6PDjV
i1ylN10BMoLqCDjhKfWrHAfo87u5CEyrPStW0XRKDTu3xSyqd1bRtzQQnNasJOZ9aGC6JrdxsOBV
CJN1f/y2oPHDy9ej6VgFqPDWkhd9zySq9sbD5LXvHwnGa7F9UjlmlCQdth9LURACMsOrctlZP0Fj
q8flezuQgHhKlb3eOjoCxvqrhphz0Gs7rXo0VWt7iUKgUn4Vo6wfcDxjsLBx3E8x9mfrfTDq0f/d
gL8YZclHAx+8GkXgcjVr7qPCwQu+Oc+9a7TuyQUnTEraWgXiNW15SrB2T/OQUGw+g4qGrWrgG/pC
dk6ROANFv0S7gYod0E4QYbMMfVeE04z1oKrGikDifAmRSXUKhzv2skeS5Nq/a01oLRTdNsJXrfE6
shfDoOVFG+2Ncp+P6/WOTW2ulyLXWB6GyHO8x5QRm4LfYK14F1hoNjepqX3TSSzn7qOjz6/eYCpz
ptK2ttp+jnpWW7WbceY1EsAXBaE/Hn3H/hMUQ0XEDzC4CU9SkX8vKMZLHmNNPm2pBkeiZGUopzFB
QYBbkmgKSoNjJoNDLuW3CsjfabRbFi3TIFFMEgj8OkljNhaKPlR+oDrOHhYuABRZdGS2Ehhs7eWP
Gx1RpDvi9tLtYWJbwztJzG+VoZfh1PLxxFcphK4dCbOwimgQaKJ0O6u/sRdoUj70hQ309k/QtQoE
vSaMqoTBEzUr4McOLSkWBWspC/vpEbIpKx82kAKSgKtwSWngCzkdy2G/i3MWH+p/N5soTM243JzA
CqA6QFatwNbriwQJfCJ2m6KyEtAwYZ8AxJMyX6h9QMDYrddTrIBTk5NhHw7RRjQK+Bx6zzOZLbUw
ygkmbYNBYR3/UohCLR0Fyi9aG5amXmvVmsrFcOHJH36Apj8gTGCmqxsIE4UGSyL32//w0BQ4w9O3
gZODd+xxrsbDcSggXo20YDgZK+Mlsp65MpR2KoI9N7oo15alUCvM1+RwjtgufnwQU/dG4SNJA4jj
QiVX4/bM2HOCqrl3AQ556xnHy1bphKsppWtYCekYOOTANFsAgIvSJ9m/b/4I8yjzMOlWoOhBQIaQ
7too3e0vMQB7msQr8bdzu+cYt7yi6jHNDl7oXRVtmodwKJ7WLsfQ2gDpJItcNQRuaNqTJvxLZpuJ
TiNn633PveM7un1tlKSPG5zMwyuYqu1klI4yCBgUw3dqWwiYzGuD4qcFUscormPhA4uOoxSVM711
8QhO2sCfHyH3rHOqqnfmKUZyyfhEc7TgpSt0VxDSxzmgQ9u8xja/0BIhlXIXSj8BJDw8jEB5sfaZ
HLbSC8Ss4a8X6lT+HZCthE1xBEwyPqZNCQQGKCHCm6h5yR6cQrNiqsfsnMgFfh2p0YYCwN1dC2Nf
FAN2yK2dymFMB5HSbCvOLPpluDuFITtHX+aFwNSY6l54I5xcSZztS+ccsu/QsENzvuR0uGTcVnZA
3oOgCpCm/EI4nWet1VpPo1Ny6yJje6BMQlw+/FWz68NFWw8RuropJ5ofMEqgagE5/U2Z9QeTqbDK
WyouBKZaQ/MBsM1DihtERJxaeKn64qIZcbh7m38hA+RZJrz96cBNPNJZzsbi0hbBBdy+7XcwNDiv
7K9/K/nzaOf59gktPylNlwqvxRPAZbgmFLLWqix9X6DEE/ezjpN4yWHNLlLYr1Am6qziB95miFmT
OY8ZRo4mm1AtxuL1Se0jkKrqlckNCW0/NDxGLfFwmb76ek6OeROHtDuwnNG0RV/R0R5w3OPzgCS7
vam3vX8NYH5iF3qUotU3qL1FO27SdpdnP/K7SxjNd4lZWjx+qn5BW7ipk24O+BwKXK4gMvqDrwWW
L6bEF1eeCkm/JrH6kj0g0WJ/bC95ua0RC9zaUSzujqqs59Zojf0f2DzBL9IVU6HUJLSN0QRs2UuK
TvivSU/mYaP5xDo24GwwnIvNt/hP6AxnyCPkE9HR70L1EAzWLF5uQSszNTYZ8KAQREQ/H5vZ7+z4
/IySe2c+Hw/tx9v3KNhtm7dbTASjQNZsGmg7jNZlgjoCk/lNw6dS/eoQzmjZC/3BTcY+2TH1iLOB
nJWoMBD+uyNdbewlzj6cp7ysV9Ux3g31d0ifIPfr1712RyUhpsdocYyOydH/nshct9mOQyDCdpzu
FtA/zrRhVfnkg50hwZICxqPiJ6526JXWCwBOT8IWslXa1DhrQzW4itGs4xN4fbm+21uyrlqfBXhU
L7LnRMoR2rVykkTGcVc9/2rdXrrlyZYzQ3HnhFbqOkzfBq8r+qxWiCmzUIZn+Ns1n/WRAHyjNI0g
TwrOYHDWF+Ea+/RnEMgR82O8iwF/oUwAuQk8sZO/rebGjMj+5k7xm62e+3FsQYOsI7jQxcISm5C5
suylmVYJ/JsX0ZJiA9lEP3QPwLEvTojrN3MjnQPPeDARwVcWmKfpafqN5jHNviUy/Rt2KkzTwL9Y
zA047vOEmms0hWADkJd/z8TYDnkVutMRItt4oc08fC3tzcLQjxC97Qwnel8uwvXGJiPh2a7jAbQL
msEXV2FmgJ/Mc825DvGoQT0wVGyXjzK28Gvs0BM5Kur17tYntRVDdxH1DaYKW/mfstoBh97YMbPr
/ecDmdYea/HrdPdrWYV1C5YIs+DeSBE0iD4rElQOGLe49/7jEiofb9ZjmZ8ypkzeSvwat0BAaMiC
A6lE54pjn1YlGJs1xZkkHMufrJctOY7/iV2BlShNbbJ8ou4AbGqYdhAdLOp0KXED0IV26JvatwZo
y28qWHre1f9V5DYi1S0t9Gtqojw40Lg3Mb+TXQM0vYHUMO268a8kem/ESQPTA5ziS8ZnXny0cQSu
VL6Xy9ZsbVMfGrzpzk4w523ZZl20RUu3kdzOesGX3xi8Np1kcd4r+cntGAdZPPZSKZVz3bQXa0IT
bZnsw8fpW26l6evlR4QmRTrQREe1X/2Lfqh9INUa6KZ7yUSpOFfMX2nQJXTWsRuq77x51kUEF9rg
24i5kUDtTlEzYQv1CQrw4iGVWDgbxKDXk5S/fPvo3yj5Snc7gzk+mqHrDOVZ/WkypEjWDfTkhguB
cGH9kN9qjEovKDvWGodsXnWZ6KUqCxJkjDA9R2Lxpi5UEU8LL8ZakqzFKjs+6KNGuqtYN0sD4cfP
bU/KaBldm6hFxZOm6Yg3N7+SH2sLreLK3fTdhuLdOWPytY/hQET+ANgiQj9O88G1AqNyHNWX0yUh
xLmMUGFS7kTYMxKVDHrC8Ykc1/bRZxDHZRXHTDkLwzf1+VcFfqCq/LYBGb/f515aBhRYii0kTtVb
iIe1Fbsj4maBXPcn/+qz6gRLYYeSnmJrgKhNKjsU3xTn6RbaGBRO1Oj8kxuivXauZGtqenuXwtH2
KvJvf4/Rn8wMpIk8WQf97mARctMnZPv1paLt8z2GiWB/tgJ0nA6Cgn68ZKPGnWdyIKttO4N2xyGD
DdlYUSnkFjhABNyYqpPbnNA0QDXd+SQWrtrB6elBn1i+o8TL81KgEWPZDDqhCNQu4oVdDebyvhCS
bZjFnk3u7iBHu6GPyhnKUBsDvld4W+uS74ilscHHMzcqH36vCypc5tg1f5hnHHsvs1LPS9krRHZA
vk0/7iQP+K4oRzMy31CDkRaUdQ0i0EU0ig75qbKI1ih5VA4XF9QksqUFei0VouLbnDbnVtHyyt5C
UKXxbi+EfexP3hXILzWx2GAapnxkZgf7X9yKO8/PaPQqF7f1/1NT5Xd1xYcDeVBYVOFVZiVnCl0d
mnk1VTn1KkA6U4pVlFWYRR5QNwLeJ00yn8hdfhhysnyIvOdnp8EDOCUsM3E68o9OPAccOKq7G9fv
NjjE+/sg9Y2RWEfKApf35KsFOdOUlUZQkfDn2pLZDLVQmn05e4/OXJ1E/HsNsDnKfExRuosnwMJy
7ZtmvsYw7Uu828nwwDS9qZoqzIqFmahN/NTjgi+wBjP5wwmn3u/pKmxS2d46bO63LEt29ZC9+1Cj
DpsBM1QpHwBJKi6knAwlg1FxkeY2FZQM6fHZclluwd3SRhWRGlbi4tf8/gDyumGazG+QPOtrG6Jp
Yy8V6F4EkJLVRozdr2NjQncIjeS7f8vnc2ynHV+mIgi3y/RydJXwhhJtWaNYf7fV4yCUK/18Aw7e
sfIhnaT8WXVNi6WpPmLIWWiBRx8rrs6ATF0pYrTq8y23GFNCBqS83LrR9/W0vW8vJMTx0epdOII/
cCFeF33c645hs/emsOVSdZpVl6OgoPYim3QkIJueD5IBBI8GaDWal4h0dC448yQPYp8At6xfnoDs
xaj45QmP6/jHnl7Dv2zE7lGnZMNjX+irJpZ37ugRaR77MwArGAY9rm/mfQEycYIQXkkAV4xKR2Ly
pqBch98fAZH4kw+xG6Urh80osElUThyDRRVmoOkt8e4H4z+X9LvXfD1FiqNIaYogFRLsWokucHKN
JOYPoMOlzTsLoenmH1d4dQQrAWxg38s3vD5rZKjwbx2ckUmkxCCOkNiJTjx+FF5lgMtIpbLy2fp3
gFMTr+NrPonUZtiMxEkn923h5sJnqHZMVinZiIWf+BDe8O1yHEWBj+u62ygLzNb2distUtKxDipw
+/zRbElohEyypJDYCkDoN5HamkUT8dEd0T/ujjWyE+MQxJp8OTteUCVRXvj2TId9D94t0EYBr4DR
AlGkzZOe+GvqWcCRmQUnAw2GwBaLnKnNHBPXoB5tO3nfSDeibxNOrRQBotjkxIlZFay86qUTusmF
JFSlMyvho1HDPSfklhiKcPaOLq/aEbT7hEuRtnvJgadsCkcyRtjCS8He5uBGnGqRHM7mZ1yy3OGN
GNECD1kS8b2j2GFe19xrD1dp3BX7PjcNDd2tyQF3rcUQxT9UuDy2XjgE+3jUbBRlokGE+YwguoOl
nSV7Si5Z7LK7cYmG5iWg8CNcKDlxc+E50jZNyk0GKFb8ahCwUdlfkpTFjKKTHK4hsi0ifw7GdIX4
SHE+cHDR4M8k/rZ5OO0IIDM8F/Gb17x8Qng/J44LfHSW11vLQd7PAHm37YvcPDlccnhKPA6jZ9Pc
HpbdbVe4FPA3ypADNJ2bUaWNbj1jFqVbcWa+jIchDxHH/ly1nHlKHqSmjak6ROa1es+TYQMseQ+V
rWinG7dDyj+BQ0P9NR1XoBg/7ZEFuv3MwmnCh+0v35UK8lOVFwz2jgW5N/6dJSquyL3JPVVl2L0Q
fD2F7lFTEyZi/xF47+ybTi8D/F5mkmoHukIKmKFSvsRlJBWTAxwcNmOzhIufJr4HkyPfQM2W8P+4
KOP3vTOMr62LNz5fhZdpjhjacvHR093T1ogAxxpBrHFJNXQ8wtjQojGvVPanMA+ipbdET2xUneIz
y1iVqphhCBCur8g9RQLZ5v04xQJd7lItRxR+KThZGA2ybGx3DcesA6n/XEj9/96smpMOvXW5cWoK
RrnM6qFEenrgA8CdxGqAs1YeUCGlZESbYIC8Snwo9rWKktNYMr6NcMkXwodaRWQ+9I0ESF3YliQe
m+gQYYtn22bAmPjxNqYoJo4F+VO0592PB0V+7ZFvHoc/HNE2cDRLhtL0UmBBA8VM6/tkfN8dSzu4
yOsxAewgOa79y6Aap+uGmX191IHNG0m2QX8AS3xCAYQGkjl95iKuzQBdX5O+5kSVLqzvWa2wE8+M
t0u5u2sbAjE65kqnN6/mr+5UAuprsr8V/Jphb/0ar2tTjZCuy8J39+4/Y4O17LtnkDKdNj/abNNT
cAikQn2kDZOujoETpHjCUxPEaUPhxzq/ypnn76Xcrs/AmlSryUPaa4uFnFEapkr3KyVuSiQnbsgg
o6JI6ux1kNGmHomAlSOU3abYgu3AvxBDejlf+Z1Tt1XgwF13A1SsJDc1aunuUawY4+gqjwcE7i4u
Rjbsufi3tzYKtHWOoYEvh4HpiZvFLnL7nKTm60GDize5Btt1xAFLf8if+N6sCS5aK6pNEboV7xuc
kXAyto4RZOq/eHnYlcbZrH+Bd2JnSA171NkfFnKNy13ho79ie4PiEaR7dPj7K0bBxdAvDZX84wK6
q0iWMzM3xNPzpSDhHMOORJEiHDs9onmh/kaObEtIU4ICk4FR47zVrCMwftenF+DTEV0A3qCp6tKV
V2jyKLsKlzipKtwheuvOnWQRWIkY88Tdf93fhKb9wJqnansR8vNdgojSLeTMGrwGG/V+8ozGBxx4
92UxdiWLatBKjW2gWbJAQDQRRSkNsbCGPdtGqwR7CYLAlzO/0Dm8vUmmp0demLXK8ORgox2DTPZn
c2IOsPMWRvsylmzfxeistEvWh9ySgG2wH3J55YiG4XDDi7uFufSg5GFj4L2D08rr0L0oanNQFqCt
RYWQ2uxdFO/LftdkUT3Bp3DqbO0uduaJ18o9W22HDpmULB6st91dgpqyv4iSr80Xg51InvwfwEnK
W+GtGcY+5FN8HaQQcsAeFlMb3Qy3t3YLCm4qRGKn+B3oa2C+NM1whxFE3Z9dTH4H3vsNLODHxeCW
KyoJrQPoaAPzGwEjwhyRzh9CxhcOWot2yDU0zR1+Oa70/3wU2EF49vlaZc1+6MPgIlvapbMbU7An
sstTMGeWK+VGr8Ic6Y9UMabYRY6/LqKTXO8jTUanhw/qKEYYEbSa9WAlwCHIFcLOvctWSjLXXnto
2oFT7t+uA6AC1yBmJ96tNLiMFdrU7AXbEyztZKK305i5hp4rWHquzim9pwvPHn/AhSQgU4cbjH5j
xS4ebEEo8tCaokat9ylVJrtSR56PLLK94Zm/rKD31mV8Q2sfgjStohbPNyzfHRvCigaoRme/iz+B
seh8E1BCXwkZQ8L7RMJAq7RM2Pf1aflrjJ9bt1DNQtn/RSGvQH3kfA2CdX1X0Y+HzZljr7v1LHNO
KlOdKo+sdf12E5RvqDVGLBndh1acmI2smZR+RKgH93yJGAv0j+YuRoPETYn8j3kJrj1M5j+GRlOZ
Es/JJOtIJwmye290RiPgweA5aQytc3IkhkyMqnnJ9+2HHI8cvm9XDR+991lw30J4p72Q8Hzi0iNy
XFGNL8rc6dGiDgP0KnGgaRBSiA1PhhH27PWg7Ineg7IF/KXneoX+uhIz2WF5e0d0wqdjygKWY2Nb
vlkkWsNTEvS7UWC2a7ITOUPdKNIyNVEz2btWAhfLlJp1/Mjv6Q4Qeheqymx43py23v+tP89xSzH1
AvYnlXIhAZhWgpSsdM/E63Yu159FYMgpmarPaBh94kirrSjYri23Z/bqxVuUgdZVWJn0hw957r4l
UZcWbL3IcVQdG5pvLQvSrA4l+atIGklcO52c959LWbUQtVaKQNjWlgDhx5SLT5jPsvJnp6ENxLCD
kBvsBYWMYkBU++qTIQOueUtMQF0Y7fYZZEh39i7SFI22hUoeEHXIPw8QIwwhON13qdgwv1doGEAy
ZWdLYIukaya+QcyVsAvNFSNixFBawQbRunoGCJOEK3RAXFfGOoY3QVnY/AqMDk5pXIZ5b/pKAdd0
q76PdjGFpJbHcQTR9L20HG5r7m5FLjg9FrPhjyjNrgdyX7ZqaHOE8oZbOUZWh6Sw4GlTaC92QOrv
VGhfAgB2m9VjtMcC/LX2exCL/bmNDW2+UwlgOmWQiKmJ6M31slM38FEEt/m27U/REl0xWa1dg8F7
obcr57A2cvdZzdE1+WPO4u2K+0+J3KlFOYF/d1GrN4Qi7lfA7hiTeXKe4+u66NqDEE65jg3e3Q1N
xtqjJHcLue1749tIiCbwntvrj+zcFwcctWRdkk63haOsxx9v4YAG/wZlg8/Ab0R5q10upPM8WqtA
ptPqhFTCjrnbZVH2QmdIMXNBxj5D/HYJ/Hkh1ldpnFk7qiM/goHmtU6hmv+BD/ebHXx00tCmgrpT
KWArWLDiVFRsNZOAUl/uiJfnkLR0B8i5oWFy3RbpdRQuO76HePTvFSKvb7a8gimkuk+V1CU4uGW7
I5c8HiFDH2tMuxRhmBmrQ4Lv+zSUeKgQWe6Dgp/I4vPiY2/lCPzcPI6b/Q2xwlt5fDh8PxpKiqym
h+gEomkkuOhoMvyoG+i98Hoq+31HpBsoEOIPZzHwEE5wZrYoAPoOmp/C+XUOqef/DpurxmwGhhZu
9Ax2ENh4c+EbyQX38TXKf8aFg/HDFqClL2idZ2ie3a/Cgn1sjAnpIeLHS5Nc7pNvQF1ny3mxosp6
8zVfCO/Nr7zXePbgUuilX5C/rOznLnm/sFHkaemy/edYAE67ePJmZeBccazGrEQ2GZZ4c3gU0KHR
mbYgsl9eMSP/ZZl2spuYn3bHQLtDw+b1OuhcFugoa6LKkW357h5jY78n6qpZnx0jdYvI8ClEFGAR
wbzsxt0YeLfq6LShPF/umbGyM4RKZC4j7J/4DeBDrnboV1ryzloKueMYkLB8kn6NZ91DUPlBtVlz
Eiiqmd/MeY0w22VaMD8/Ccnm0DM33lWaYtfkVz2GeikI5lXUOOyuNbGWdOQx24STbin/xmstUfm3
0vwqbsPXBGADgCAT9VKyBNUoX1BjnFthYYpCYQ0/YIz1Tg8jiEw9iHqmgNy6KHy/EMmdk2LW3hVD
PZO/AWVYH4eZdgbWfq8SQqFyA6E/Qtgh6iUUFBzxTikdXho4tx8OK0gleXVsokMg2J2OHzciJRGs
/YEgoQS0GURh3imhmFiZkJTZ7KfTWLqdqbIZHkUhHTWtJtAfd9dtiQn7y+bRwrgWrkadrgbb8aeU
T3qnhdtlcssi7X01LQxZLsn6dEneV2awaeLxj1Kt31/gO5BqMB4I1/RWAoXQxEq//VAiK5g/5/kw
SfThrpORo1odWikXQ1yJKu6+Dl2o5KayGk3mcgwpJWyZbKh9q4Tn9FrGF/GRbQGjHjD6c7ILyA/y
oUwkHuY1M0USahPPjIWIpwWeKmdSZDjvNsZuVO73GJeqWCyp1YWld7K99LNVxKTHWYTNLYiGAkt5
dt/QQjrDk2XMmja8P5CLCMvTUKAo8fTfds0lVRbsesIevcZkcsgjr6Tq2zUT71Gb1n4rN03I87BE
vZFz1r3yWsb0XZ/me9GlxqMD9NbIV47OrJJG40WStfS09kOHNkCDCtOjoZc+FQDZyz0kegfwtpIL
3WLS7d6QvjsuisTi2TNDXYzgm2FYZYS3IMkQQV/uJGk67PCWVKpt0eJuAnmEJSbivSxHr0Jb5bMA
pItWiqz/jFXBH+fUCkUqWwbbHfUEdEmLjW6mgPM6V2JvInx+zFxyy7YEZ/dndXx8p4PXrJ2JbAkW
JcvtTDnaFrE4gDMU42u9HSpUUj97d++kVNj1u+w5rASm75JIe7ZZ6Pi2hX68CVmL4V8M0ht2SonG
HjeHoMYru/8/tZC67oBgLqImCVsWnKIIW1LnwPSJhPu3uAGu77WJRvqHOsJdUuoq43dCU1DTS4hh
sgpQZxNNsM707byJ6u7DI0Ow3iPg3LKiBAZWUy9oKeq3mdHzDacebhzVVAwdheXIQdG/GdQcR0dU
6ggNtXH60C4vdYFyN4P9G/gNefAYPXlxCiCZ+RP0YbXxA+JDL8/k42ThQabY/W0bLOmLk7nOuNKs
ZZYaduFuytqF0ptKscIQINxIeVfq7Tb39aun2e3+uacjkdL0GI/UcJ36uRZfKdXCY+2TwqRWELDp
WUEjgDGxA5+9n0HIV5PzTKN+wr7e0UuBbPuTlP9CXJvTrhbaeL/bjaXsP0xtzpVRsqN8GItnbCu9
eqsZlYajMTKO9bm3iUJeyYQ+mXS4rW+Vpaw6bgqFtlCUaEe80lIpVE4jogIBy2/yGG/hiO+Sydl8
yE7dnIc4purmxdQ5Bq4MXVdU0CfiGunHGsA3RDFP+SDSc07WGBdzDHnOaWCMi9P24oM4Co4utkkA
dMiW9POZL9XajmDygzR8dL46q/dUQmDWWh4KPFUJqydkwDj/GVr6ALd2/z4Zbie9QUr+PhuQx7Vr
SomKN0OpGEZxDO9Xv+r5ces4VsXn+Ebqf3qs9cIv+bZl5Qnj6AMbWflhmqizqdyrXz8uwF1julAg
SbewAKg6Fx3AKhNQ6MS81IbegAbLilDLi2qKSzbrR83/mVSpNj36GoSlRPLwxzMsPQLHG7bntor6
AbTuiuLNBYdk5iGqvFjVjTiQ/siX7P2DV9j5PceTfmndP2zCxT2c8IJ8Rhk6dZywSo4dF5/V57C2
9KROXN6EdabrDwMPeeJxV8uToCmgtq/6tgIfxBcz6Jhz9vaAFGPxxA+1eMQnvyeuwoAKjJqjqfsX
+6aa+8mX8w9R7b2k7cZlCzhiLkg8m6nXjCRgBB2LnmnWRqL2c1xXxNoH6R5Fac4hIkQ5BaYwyMIF
azgjZGV91EmyFS8JqJgro3x31seaHIZ6KLw+ESjAka7L5+bnbJ/nOxehOdwSlsj/QnAAPU61R6C0
XWrZuIvYYw7RUt6WyWAm1WzIXJRnjn4htm/Bhr5S4Edge8Ph/Wy7iOkfftxj9XQNTKjP/B4/63xp
nr4gpB4EsVpMptJo3/j0R/U6YSaCFeORpJwMkuxVe1RbpIGuIUPhcNZeE/z03LnaDhTxSfY3/aQL
yUXfYJmiUOC3GzVJdeyycMvFr6CLy26tVGmuIBAm3l9P51zcPwqM7KfTrGjpltQSbbBtT97uQOEQ
WWO0i24yMUOfrWKeouWYTcTtKmWyNTLdhHsFSiNARAsltOcDyPumckqObuRXgPypOFnO2X+A2U0r
3by+PT2L/hx7IYYiM8ICrX9HAtImmsSBniQPAnhhdOxLQvttMeYfh7tUUKxD6wvya6XYIf/Jlj+c
XE2I8la1rpuMckAR77vLG1y11DV0zA98PGxl2hOggSxM78U9yCkvpSRQNtRlwZAaMabvOW3S/iwe
Cc59ZvpNXBXhcJ8iXbPyi13kSBTtJqIozTqzi9V/HsZLxP0MtmDbKIcYmukt+6+gTvLdm07l6R29
/dWYwp1ZqRs7ibfebskZdmoh6GwhY6Z1gzgpvKj5ym2mcd48CJRrJ8ssUbY0VByFin/PFdnmgdg4
6K/4ArkUfug/RrCzPOQh9VVHfx16lBbWXeW7rqmtXj4AZuUEcZRqecgLB1uNHfbYQFMtXB5tzICa
B4EfCAEKnWLelZQrWRO8gbX+E/lvc1rvKkZQy528OdTU42Q+gp4LMqWR9e2QmDgRx4Umlw0a6qWG
Ieyis+RFs1wtTNjxLsuibg9TJMECyt2EgyUYe8kkwZRvkKHS1gxvl/PjX5ZT/SjVn4C7+G7ueE1k
EHk1NDFAqmiWo76QuG2mMb6EviqvY5Kh2NPRa+vjincyT7zBEuR6jZhenj+5jzi1F7vj2WR/3e7U
wNXMO1K6UaUtFEviGxx2Vs+99HqdlypylzxVw0WE7nQ15Td3tUH+7o9Fg3jCUcNtXFPI5X78NQgg
yC3MmjfBHfwxAvBFOf8WiZm441vk+ANTPqVENYguwT3J5IJIr5jNgk7N7UY/0xjGljRaPVZ8iWvg
QY+NvKr/k1oIPbj8wibmv8f7/W0qCHn8+kazmSkAdQvIl0WeH7CE7AYDv5L97haQnPrU+aW6f/bN
V4PncTuqD1XoRXkY5YsMSkpk5O8ltf3py94bxsLHjDSeI3yxVmIEn1kBYUN/VnI/XCo8EBzeFaHv
ONRnt+Fu+wlV16GdiFU+Am7WS17++P9rB4Z2WS5EwG1/n8ijz4iZnpCi1vEwHW5kftWjkYhmMHm2
HSzQjFYO4e+G+a5Vl2vQQ1abRXy84bPxqKCtfMHFNSDmRRp9Ta7KAIsfNv1LgHAEj9mCvM+AiBlN
fWvW5iUooNKUhWsrXv+0wUhpsbGio3tKVeUry+12F2S8D2AyHLMZTZ/1EDyKPYYAzbW13Ud/551b
JBzCZC3F9fMMP0ws/+GxMNxczqGMc/4lfWwy5TR3k31LD/ib7PRAV5yXgor77UyhlnY8UCnhTNbw
A9tvoX58ru0QURBIyGT8/CdQtTOB/yyQGLMg93E+ZSVEQUvgUegu1M08+XzsbhIFLwGrmEX6aEH9
Jx3nApD9GRS3MEDfcUD8HxB9ke1PD1SSbVrO7MdqsW6k8DIn+iqCATkc0JpaSKNdTR84ouZZeL1Y
5ei1WLXKkYMw8HaFIafqa4wY91WqZjnhfpESMKXWK3zkn8MBoGOVFwOpf9yAzpjwkPIOZdwiMoqI
9xJFxutffC6aW7gZHqYVxMoXROK9Wm92VkAXATERELxVn/nqXldzcRM6WDHUchSP9RKhJNRvwesQ
greUHpE8CSMBYi9dkKfEIKPSLROCNKiKrdPLtBSpypkOXrmkFwufWKo2G6aF/7jgRwK4lXfvE/rq
QkCmCT7ZL+K4wCODYSoH/yGWtI4nZ0L1GXEQiPIWTa5NGSDSfas38iKAXScw/zBOrmORpbQzy8vr
4APzRQ2i1G1EyQscfAievaiq3VO7mFkhCvGafdSSU3NHn0V2DwmGx3hHqaP8LqhPD1NEwRyRroRd
Cc8Oh+Pq8EQ4qJLRGaIYwUFtRTLwBnQ86uFGFhBApzY1r1RbRK/sYb+dQYReRGAbn4hiOUhsuwux
lENazI8DhlqK++RoiWaBm9Uu4Q02Y2iqa6RFO76hSql/UaTb49K6z2pjybhOn6wuTCDEC21t89Le
Js8u2eyGC42PVzMj1ojt5cTMTK9gu2wlTcPElrS8PHspHiGiA9ReShjw8ARW3vHtKb0IDWpYqOyL
SDyBaUGBTBfYREeEBdiHOtLxheZgtoANetKDdRa5ER4r8+z+7Zgf/UYZ9LN0m7pX0jp5oh86u8JW
pdmYKoG6ZnEmfN3Vnvs5eCKZ+QCI/XGSWZb7upX/ksfyzQIE5KMJMS4OpH6gTOxQiJcAOMYAuhpl
xi7XlwkZYPSMXYeAHF9kqsGlYyThBIMRQsSqdJqvP7zbtut1QVOu0LKLftbdZTNgjTs9Guvlv4X4
F5y9cZ93HR7g3ILUUztzQbt7rQh1cc9zjKmzEfqWIKg3FEuctsMDY5ViaBRxU+hREcy52Irf9qsU
2QHOFWKJVrKcrf/IrZDFJMPfkobk+NyP9qpDALflo+u+lM67bqAYg6JT6eROQxi4+y9jQ+5qYmfh
+sN4RTc0jjFojCB/4iibMkEva3egUBAK/MXWCiS7fqPvDHm0/bTPNMgYKDbvpGNkDZJg8mG97mx3
vDOmc2sCW6ch4vSjSbdOsZlUp2sVZ2bZKGsIYPfNxQ0yBU07Tetpjk3sJM5A1Zh7VGehATY2M4mY
lEm9aU12Inwl8C1jtuTfpMlfn4xWd1y07lOaiAWwt+JnpaGXjkJnXPgBWsOSn1x1E9lDWGjAAU72
hCsH+nYLnvvzg5R1x+D5awwqPsooj4VPD6UCML1+3+gnV/VjjyOwz9tg4Pu1oHvobFm0McDqTDU9
2WWlnAWVP7lZB4YdFdNohgMpNjF1ISWGudR7fAm6hCJENU9drSlKD0Z2nKM6y695uVNDx3qQNVSU
Q4X5vBaXwZfLJcPvkEyTb9oYaPMR1GbW2/BklTIVAsPIg/d6GL3IpXGhURmRsQ9OHmMWa4xsFswQ
wFp8y3BcH/FVLgwE1rkh0dRpFB0sHNLLHSqowCjO48iOfovYKDK58LzA9j62D7EjzQkf8hqfLYGw
J1+VkVHVuTExEDEkzjQ705szD9QZvmlqpAdWKRhGJPdHNB44hz80R0V0Q7VHJ9ZjwXFH840D7BU2
N9H9r6J4b4w69a9tkH3rV3LK9ed35Jmjo1Z1/JRB712zPol/asufgkaAXypIWWTw/yZ7Fot66wej
MqP5AautvElpyCTjVkNIbYKvVTVGk6K6wixCqkHpT3u/JC/5kPxmDP3eNdJL//5h8JYDe+6aM/s1
e1eE22MQTTysHzUCw+UyKM24sb7LesLS85+NGQ4Rdhp2N/aPHzyLcX0cEtWHjeIzxbjfgl+eqBLa
7BG4R/HaHZdHbsQvWDGVf3P7zYG06Sa79Yn7f8o8L17eZV1164JzKcbB4MaHSvbnUkJLG/SWm4qA
oWhRZCgGU9t9leckqdg3Lf6IevXde7bfyySNepY1hobhoIktYNY8zsQZ/I5eGkG+pR3s4b6LrHLo
UznApKMvZHhKa5lI44jQ9H4k2Ze1XVAN58JyMgNtnvDggNqmCdMfj3HbjEVhgOtPLrTAC6GGQ/6F
8CBWXS6TCZNDLmZPPDhyPyKzjWBmMW3KL8sowGYJNL39IopiDZLpCWL+6l7D08boavmL8teUqivU
QmpNOS5jmQGLDrLYA8d5igT8naNKcrw6RZCOL9C3dcQ0wI/gmAIQshJZ/SXaXFujzTBTpZXaojyj
cZVScamlUYk3o7iJDjwB8Pd8dMClAvKCTRSO7FSpQPXPvpzkJWQG7T81Yu/gPtyoAzWV7m2thO3z
psE4ymGrXOp5+WBf/knHmYehGxPZKwrA6ricwEWhg75eXKdYoLRJrECA1cyzOncU/s5/uVSKVey5
uU4pR/JqTH5jrGUb8VE20NjHWavI3v+o3Era/tpX56M/mxv2fKRF0sixWix04TTPSbFpGYJikqBt
fSxkZRXl39f3mxwEbXNla9klA1Gpq+JF18/jUSdj8CPSmua4vkUwGyEc43TIUmL88ahnwnFiIPjK
rO5CIIx1/zfOYJxG7KVK+1MEuei8U+YXB3DgWiGX+Y0IHOJBeIpI6OjsvUl+7Ejq1HaYXvGIY4NR
7KqARvD0UHxN6lweauw4P0+pDpqwC0dCBUiAJTR0zGmvgR7T/iEsoI82PIopWmIBGjjSoecD/fl9
TRvihqvzXR88lTMuesW5kvcHDxRD59Bqj+4J2EomyX6/gUJSNdSkVByp0+KwEwTwMpjP+MUYygKN
nkJrjLe0euCaj5tcRW8TeQJDoDn1SBggiCpGPfxN/lGvuXge/1ELM1yldmK3wPf3FQdyCJrT0ifS
zB8N2eEOMqYMNpjHcSHvQzv+G8SuPByH4L8gyxKtLceRudkmbuyTc6zNjiMC4cdclG/fM/TkTCjH
DxhMUWv4PP//pV04W9L4kipmIQ0N1nrnSqxFwaF/cLc4KiYfQtpoaYEvKMUBr1wSvqFcLwwPQWnH
YbVOU5utmMidKR5DM4IMcVDHXMpCYXrr/9zEElp4rhchkynZujayaJKMxg+H5DO+dwUXl4Xe2oWi
O+LeNKl+SJXY+uwQHQfDjyzXImV5EnjWczwetlnRcNxmM0bgE+BsYvVyHjCluEziD4jk14H384BN
z62r9EeVA5EWyHD1Df7qg+lXyA0+XtVBHkEdBvFOb/sX6TTeLLPd8lvfuTJes4ytaMEpLfIoTQ2M
wXhTK0LO7xzGuR12dwPFFLAtJU7a1NzLLU7kDvvATSRJYC897JnoriqOhM2rfjcesCzSA8uOk0Lb
xwii2+rd6LmqTxlEOkAhBh9m34jutvSTkEa8SyCAnjByVE5Rgi+mft4en6EvBk8LD27Iu2RxRiSk
oDho2trr1YWOnfd8x/6AGDrp9leOPvog+TobjCdhr0W/eLxS+o0AXtySe/UP1G8UEnWi+FbWFoxB
NyEkjW2/0RhDeWME/Tc8MWQXwkiVAOcIZPRF8JTbd+blvrniJv+OSl23CRjryaRpt72mAFLJeIXT
hqwccpAUavRcsbEY5Jc0HJr+EkBrPKy0XOShK074trfiKL6J0CPnKlE5mDPoEOwTWNz7G6jbULAC
hH/1WAkhItfxuPr4IieQiErQ9xTe0gYmYaDzQZFolazFFUFH9pnvn34y/radZAK1TNL21MWRqKle
nP9SbpMi7pp5gD4MmDEDKarjklCU/hMWdb4f44Z2kfrwKPBEwlvQ95aZrK/jzDv7qH8Q15JTH5dG
wHtArudyxArwrAAi0bz8jKpaF+zQ4aOVBAJJwhmVS8L+7B/637LK90pQJo9IP5QtIP/PrOivEOk1
Kj4aYj1j9vyuNmiTpuZMeij3uCEnIpZ6HvosG9pCg+UmH9Zgq13U69UH/OaM1e5um0b+CpU6yTfe
ZgmQwVIDiuyb3nvIfLU/lU/cCsy+dKzB3K/n1cNMaf6vbvA7VbHPJYljaMe9PQ7uJ4xxQ+VPSzl3
czdbNZBb4uK2Ib6d2PXHG/3sn6mEe/6ppecFJkXGuO/gXJYlVJBpD/eVQT979qOftuaoE98Rz6zh
1gAEs2KfFfb1kRyghh9WNdASKTrm/2HnZaNJduCpzxd0E69rqZNSeZLNvnttfHm4QGPC976x9Ra7
7KPBNruyolrHdtP6WN8WP7y6v89RV8hDjSfSZGOSH8yT4mBqi2/IZN5KfqGTNemhltJGq3G5SYfV
OG6Z0JfYV1Bil+9G6d09wLLf8+4DSSf9I0svAYlMe6jPd968bv5NNCRqGpEqYslCc35DU/iGfwK4
Jqk6uVrwRs5lr7EfjZLP66iPRtftUfuPfLvg7ydGpJ0HGaBCCKQ8z9yOgvg+5ZN7/JwYRKt1Fu43
John8aFkw//ZLBiqZvlmK5xhU0AUxHQmZ6/IDy2BOLopng09Rhs5cRlFEmq+W2Wg54NOcWwt22ta
0lL86dthTgykO705Tear7qUNXlJfZEQAbnENKwgHswiGwGeKZIr+hn3YMRRxy3JNbGRR/zQUFC6u
vbBAnM/HDNI90GRK7J74C2yvD9dD7shMdf/s/WwuKihqGhwsqLtPwfjSZhQDDFVZgOtZfhDnQWyV
ynuja6OIs/UHz9lmCe1Mr916XdI1dkBuJhcwDGdxcQyL1GD+Tbrfn5Sdve09DXDs1g2TVzE6ThF4
f1xewUMDDi/Fy4JtSpFawKNlBl+Xev3MEA9j833KvJbQxqmZ35XgjeT5KqS7HDmirT9WELkTkGUP
J64AgrFbnWm39UzKjo98uLZKKrEQfavngNT4N8e9rWQ6kyWMVLVpL5pBNyysvAxJ56Avw9dwvYtt
jSRwtHniE4Eyu/VngMEXfUlFvb1otzcHBeTWw/3zoL0e9q5dVee9Uf/By931ZTmCg0yJ5JCDudCI
TBnpUn0dsqpXkT2oqO2BY1zLkrNDgKpV+MbMyV48rJRcJ60gsyvw3ZfqUZm2eE4PcpVb9JLf8xmc
nFMDiv7QDeBaXaE8z1FmMM839HWPx0pCzOOsVYyhfn7TKJuC29T3eJfkc5++PlG/uDG98fPOuACs
HXpZMzdVWOT2VlYbAId5gH2UHGmeFHODqHjXOtjVrjEaBBXPjZ6XTiWKttxAHawNE+2gf1XaOBgW
spKQijGrb3LC8V3UjrN6zip6RcD3BrbDX+8lCqRHcuP7GY4ufo+IkQ63DN/L2VQ69ezJVhGfCk+J
3N0m/QeGn6KU1MaBCRjZpxG1qtM8kRRZsYWjG+A+v/S/PWskrNthr3YWngVLNcdvN/Pp7u1Gf0k1
0Kvu5nSrHzVx6Vtn05W499dxjbyLOOZ0auQ2qgmarjPNxB4HffPF9vyF0tclzOlMXSbhNJY2JhKm
KoarolwicBmi/IcQNSdtQRTadeuCc+iAlhTtinQvraP+pKLsAkrDEIhWtxextT11hNEKWDC0dLsw
UrKaT0oDRbHx1iESoVGzSMSbz5+mBE0Bz4ie7tTZZCJma55KXrl6giOKgxgUab+Tk9MRUBe0+OHF
79UNqDA9jSOF3l1rc7+9eJ9InOa8Q62cY9d/zsnsrwRSe9WafQOWsqRhYeTK20qeH5DS5EpG6DdF
XFvU1Zudvpu3O9KpCI7yVSk6ZeYEzargIhE3wSpaiXILq6Y6iLetdNg5cC6CEj11k2cqj62FEIqC
aUi7XxfHTDslQF3TAL9bm7nBidFF4qcuyP7ngPO1xOAOPK3O8z0hwqI+h830IWu8fv7FYoocPxf9
uN1RuqMergexNkCTV8L7jbWCNLdr7acDRSSlcCISuB1XwM1htPRVHu1F5aD7l32uwjLfeUgIQrIu
VZ7ivbuhcrYI2nE9VE/c4vwnYTWzNZSNDB+bzAtoIGTzgLHZdpXELtKDXpUZ1giRjXiY7m9qczOP
gGjXri/8MMC3PRvoLAqe/LoOQdCgn+uCAjw4w07BM3t7MxqWzASWfnuXBLrnAfv/GZRvH1lflvsP
Jivq4rXxvdIuJzLvoBylP+jdl/+D5hylR6A+wOjV5eT94Ixtjem/7nW3pLcpZyS64PqrJG9pl7BM
Bcm6McFbwxzA047qlTkwnoxwjacXX6LI6rx0jsjB9vNKfzOuT2UGfgluzIWvIaH93xXtRmcSsygL
WuI7oAhsciE+Mrxe9LIThigeYs9OZxvMqWI3O/P1f8vcC5bWbsTLu8SxJF/i8v1tmAC4MUUuXofn
OXRhGyQXVy4ZkJLF5Pt4dxi4CTyui3diolKqFVDo9sPV9n7ecdRJ931ZjipvAHi1BWk1TZJNQiJv
gRrrRtWrfe/RMxyhxQLAZMtITNW3NIAgOJZvzdlaAVScsTZhBur/uA0Bc9blzBaehfDnxOHvUXym
TBu5lFgbyABQxXaVv6FtUda8vFgNfvmSc4LPQMsJWRL3MffPltXjb5gWiBwQ/vLz84dBXM7/6+dH
7b6qpdqq71UwCXeEQP5FNx8YyLtDm8axwuLGRHeNqZ2g3MTU4LDwo50Q6/Gn2mWNFdbBV3EVz5JO
xjjtFgt2qBM3piYE2QcfZcm2I7OkeTO9N9a33EXCIFsE7CBCp8asdNReiTtC3WbHxCR0nQ8cZgZK
EEnHifGINcsPAtqdqjuxspcMxvzlA9eRXsNft9PM6U3g+XUTSPIHDlDFe4d/S9OI699s2xjl74u1
wKEDOzgGW6PsdXUprk9H/LHvPT6ZwQLsfbGOZQbrrjTIY8RquJIHmjMGJRKHJ8uFYZuakqOoXUa2
zmrPTqh5bHsVQTD1rnVKu2tWUceEZdd7rbVBtzsSpa8c3/fKwhiYV4sn3TkpmnyWAhl1ppZ0EUlC
kfhqqwSkqyZqnah2QgWIsbSEX+k8LOm7U2PE8BJPFqOwlXym2RyLU00O7IfVB0e+5MFHQJg8pnFX
Y0fV6vajwNxFaX+o3wo9iVDXvAjJNsVSQ2JlF0yxuQO+if6asgQ8i5Cy3+K78LIpCC9S9oZlIv9V
++HbCctpsknD48Bv1PR0inKpXPdLhv1s9foUJ1R4rTxh9IU3ykIeT+TRlyhuRncv1BNhuAhmnMFx
XH0qXNr4jsi8jzZsG2NnS8R1/iZVC4jKbhNd2ymyz2N/oGWmLZHtbNfEHxwc11s6ROV5xcFiW+hs
9Wd8v6cnhGx1R9bK3ScguXtwxVgDm7Hs8SS9Yujqbg1xbFWQbcdC1vSiNr8KnXcvfD63E4djjFgX
OQCzuvqL7TVEBSDgZbP2b/9//IIvXdobwlP3fksaQ5MdtlCvkiosRdjnsyiaZiKVpDMUs+NBhNcE
LISfviHpX71yg4xbSo3TAHf9DA7pjl/vTNtLg5PiaRM9Ai2QVJa6dAwmeiZNTBmxwn9zKJ+hJTTM
JmHjrp21xb4huctXHLhWy8yGOpbyLaBnDFoTbm6tQQ3pS1NYuZ7cTSKWJbr5Zqi5qj/pxQ8J3cUv
6ZFb/dQ+VPCvuZ1g2vi2iVRuuusHYwd6ZWPTMb3cssy3zlV92BNT34bG5CYDD4qo75l2z+UxRuf3
xNBm/SzeO4caRwm0xT4HkF4BucCkH+rPPfy51ziGv5CzqHOql1L1559vxS8cUlEdo45ma3wkyXYc
OLBRNZn/OaHMlWz1xFpKioGVouXR3E5GFB96g/SaLHr3upvjTBMfpH8LLbO2JKA7qqfCjOEqq63q
sFO6FUcG7Q9UUyzx2QahrLkFQjvmJ62qFBVLH+LtjiMX+NZj9UIQyXrb8ikjHQ+kl6uZ6/ewMrq1
mShUl7b0Xqn9jJ1/jo0AeUCMIbQ+q1ZqPn8qJZJAJkCMALpjL2Lu6qiWiUfyJxTv7RvH/RHDU4fw
oyikQVsP+Frd1hF0PFtBcJ86s5MESpz4x174XMTL9E3DxwLaL4i7GOiYiTMPIoE9Zfd54uEbj30R
s1zpnEM4QAA+vcQLsVYLqMZjslPoM6JzeNmVZbCmGdWU2oVXOrdzvbns5m1H57N8AjwtDq+bghJ5
IsnBmvb9wVpijjo3GTep3cmgT3UE67LA0O/qTRbnnPPP5ECkNseGJ436tQGjrj8zc2/o19rqcbpI
r/fYa1UvHOMzUFmWUKCW1G29+bdtzjZelyzvWGlePH84y4AU1ELHUlR/rvgo37lfTOF/XhRJbYYB
HRbprtDruwKS2gXMbblbyJd7a5NW5hYe7/0g5qSoQRHss+sEPLFlETNlO9XyOj7V/RyPj5VB2x9T
OCVcUQR95XQo/Uo5C0P2aeiljAudVTSlxItaen3RKZxGUOhsQ2y6hKEqPuxlXkQwsUnpC5PLbb9P
rmDPyGsAG7UQNxLUIGZ61Npb5YR+i4N2kb5f6npkRI2znItzwP7iH55/Rcs1SZeHooFLMHQMRc4P
wxOD5IexEAAxpHmao/6EW058H84me1YHsXLj9H2oGoPrndhkhN734JHl37kulC/Dx4KnLF95sIUi
TkdJAhaQb9svS7B1hUVwKRQ/kClJXtEzQ0mY0svsZLtOEbCLFoxjZ9EvWJP/NtMuRYYbUj6J1VP3
G0u89MZR+wCm7slJsgf6BCuIAi9DDj0rknGxtIFx59X9PwAFF5WXGWHN8IcnPmP0HAxLmF0syGNY
us9cxgvIZGz5JAeqX2oFjCG8Lx0g9tTgvOueFyYdklNt22wLK+SW+ZD92EqSqS9BJazfbw5ZYZES
pOywZTDTMs4j4Z+sd3pNM5x/zC3M9XUHLVumbUU8SvytkQySiwzFcCs1LjBv4IYO3f2obSS3tFtd
dU/CSjAw7ZIFxjB0wofsP3PZyZrYUOA/k/kKF6yjCpHcEatuFzUqbJo+dZsyQPtZWF8tfXaYyhlS
NDWsNsURKVhBrW4YFCNDpx+NP7zW74sFM0hTxdB0rbaP4+M+qbGhiG5e1S/GDeEKiVdbek+c9ecA
A3h5TZjtI4lq4+IA3HOOmC4x/2FdFjWj7FAlNLkOQknaTcxjx87nv+YY4g0p5/Mzd3X2pHW7bZRC
ZErboJ6/uqGrI4FUwNGdswr4lCQNNATmrBV3mTnVq7kmssK9hJkZ9oCALOLA2hPu/Fg7td6qjMBU
7sYK1uGGY4CfIxKRN9uQriH3sR8VYVgsz+o2IjrD54y0UuK3MX5Ld0rnCJp6fgTcwzyEUL+lIGRe
DtBpk/XwF8Flf2nyT5liktEZuw1jQPJvEMFipIlUZxtjBQul/3dgTt1QWDVEF6etoybbzVwMsbOR
d4s3k9crCJ4/Sf3BScdqRspeaRJig36Ul04d8fjPNF4tOTqMRKb9weCu94Q8t2hMFxSGKw4qrw84
1JGyeo0wCFzGIs7e6qYEjOlHLEqle43Ek37frTFA9kaXYsrMVGB6dNx/Y5z28c39tk9LRW0P6P1x
JBIS9vX9JIVYhO6N2O1+YM+m0iDb/95u/FrsQ9rZUid+uviQkgjQlzX6okvdZm78VMk/XEGQYHK+
ahsht9GfQpszM14GWxoWaEeruhHr/ogvXmqqrA/Rv7Ws8x3SH8PFwaVYVMS2kCIfR6vQF4txu5i2
tXmNMEmKtoEHhu32v3SX5XHgGMdwbSVhWI9e7QwcxCd06G+K1SWh3UCOa1uOmutbaBQqlEMdh8l0
yh+GEzEuRgylLVzNNhmZucKBoD+ulrJtjWrbz/MaZAir8z8zYbWpDjbo/xrzwLhmz37XS6nCTHZS
fSfZKAsSDvbg9J6qi6iYOyDzDMszJUrdl4rQc+3niFTNJb5tNRabrjK8YQk8e3Hda9f6HiCdKTiU
RCoa1fGQXdpNWidUwupB7HnCPkYhDpuFyVEJfLs2K+Ire13klJrQYqzi4Zq0b6mhDYre/0UnuRYI
fLXJbc4fz5tNr0wmvx4P8wHecUj9Cxkp8KdZNcDkVpYxBYzgrvRTjVd2NN+S9mPN+355G6QEiq5V
8HJ6LpxnI+ezpbgwOIwXbiN/fNplzjOIp9VVVTnOS5imnk7f4mVmCwpi/r6pHtkT0vWIcujdxf43
1xUFmsXwFPywdBX9XYTsl/CrDAhKQyT6Dpz6GO2DA23nbPhTva/+16v0yELcgUmU6L2RjmODliXg
TmaFvcoeKhcn3rTO1MhmjZZgfrzvqousD65bW6joh3WmRYogguaf3yhirLtpVjg+HAnVFEEOmdjF
Qmn1ft7qi19c9wDmQL5uULqa53cXQFyc6TF/uWXtc7u/tdLt+RSBSWKh8f+hxUpvBMg4QG5BSUti
JRO7miLB8/Dk7f9Z9SLpmhi2Kf1xgEcI0ncA/zsh8A4XpkplaDbY3COxWVGZQ1KX5visLo2/Ah4B
RGBF5Mq0xN4UDFHy8jN1gMJ6qHvdy6Iw0t56Ubr/GEeC5Ck86vDx9HevI/hryYP194r8prtMMDoo
/Xo1BjqUAOJ7KO9rvoAf10lBit7JhOE5h59zeOpZAkOg/cOhU8jnGSogUbUAuCneUZ06k/ATX4dT
Gxn4EU89g9qJxYGuFhdfLiSvpKSmAG7r6P5WHrl80lS1fMTvqKt78cNZtWJdsDmuYgYMlo891wqT
YR5uacBIN6mRcoeTn2hPG6OWlJLxAlra+yX97ar5gg5pNgRDXUcINLBi4CT9IWeLE9PLfbA8h19k
E2Rnh+IRzOkQm7/sE507o0LSyroHAmN8RkczaCNTnxdcqHnh4jUWBVv1MFvs+xH5sbWPws+x8PPf
8VS5a1caAkLSFDoExIbRmxXKS2m82bDS3EY+Hr1hJKANkKaME2HZRucPvQVvLqjd43U73Zt3IB7W
7OuXPmbZD7GqHFjgyAYW2Z0lOeQwv5PaJe3tmoeOLjdkShqwN2Exx4ekBDixR8McbhxYhZOZWVhT
0KX2VsymJexcUSTGILgAY+qLHzyEwRncBS/lLsa4eKNW+LYm5UotJtoi+lZMsq3P/qj1k/SiwF9k
QjFYL0MI8y8vl8SnGpqPMyG5sHwUfUUhUtnttbkeG/UoivcsxqxvPWE1F8HwhrZvKUK+puNG+vNX
LG4DStPmjmdaN/m6gvnKQVmfu+kRHKfamZaQsoSIAoZaElSa3f7PUfzhv+WhXVNi5TgHvEuuSQpD
z7QbV9cIBj8q2Dvlt9KT69mRU3lSLAY7TbZnfZIowkhuuVLCNFukvuNCazBq8/4cVQ287BjAYkoF
BQWZvbAHF3CCVv7hDxlpjlfO+FJ0OTqneSSJfl2t0rhr4DD8an+rEqCxCsjt7r5u2PlwNL5gZIov
qqUfxapwPnBy8a2hOLWjV88DsgJ9i+n5iX9uXDbYdUB1G+ofGRGEEfcVYFYyJHemAs8uFCkKEpQg
n8U7jF2tVCgjUddjcpRaemGj+wuVBUyw7v5rT0yY5N+ZuVvSsrLXmKLoLc9YkzUwe0OPhapTRrFz
Rq8OmLJkQPzP7edrzzLkyCy2u6W5qbifSnsOJ0g6EQ15lVKAPRQVyp3hIMACJFrSr33tK5yabKGi
hbfYJ+IzWvdkBnhqTFL04iVuCAhlCFA4RLjnKfq4OnRAGtVP7BdfMKqnnuOHZiO7/iris7zyBGds
Lb0WmAb7qOBW1pYSRKpF2n7tOI02hT8p4Q4cKuyd4rHwQS/x3yGbHMhCpkiQT/Bb0eWJ62KCMZYL
wduiUEBkdvqOhq0wpB/txMrgEasfBrNKWeirrBXxmriwAglcpVM8/tgqD5kki04WI6sAHmaug91e
sExcYgeDOtbuocseV7kEClw2XafoICcbK/tT0Z2yUrPTpD5g2CRVVs/VSoMdUz6yw4/8bEnXr7nA
2Vw9vdMpujYaumljaIQuSjcsPfderDxWnwcaNDaTcXSyv3245V+ScAdy7u4j2t6KZxOoXfkqj6HQ
L6/Ex5STeRv0zbie1edHkQCOb0wRHEgLDZL+ZaiGKFFhBZ78Up4RBYdRYXx+F9s1w/q7AAn0VSUH
8oO9w/msYjfzCWJ1lBF0a9wUhVYUsAAqJ+2FLX6x+XhJ38wYVtaWMJwnZt7pAfJltZFa9vPR1ohR
7pqkA8aRKUTswQaKhUc9/TYwifMLGqhJPaPPXqbAvf3VzRPAPrAzpF1Dxh3FF8mWDQcaxmloh1Al
O7L5Ue83N70I8B1x5OihN+T6R+3GKSuTGdvqwD1dbcPxgEXX9MB4DZgYgCncQUMAdhC9JFjG1nLQ
sD12qjgkfr9eWbt2LcWzmPpacEUCs/0i/2orHtmAogdMKLlA8Czc8wCehLZfxhfqK8rY7yKoBOtS
D0NhYXV4/Qp+hev0Qvih03z7m6df0A9f3xAn2F9/++9n5XNoIcUMD+D5CYIfpL18hNOzTWJXyWIE
HUppf2EkP8uKTcVvDVka/85Ghs9abXAXqHM6snB1k1vRYtxwa73vbjZf+WSubF8FgmAnxHG5iVxR
Lk5WwIRgvC7y1nfChOemDp0YAkaN7iUEaqZkS/8USWKBYnfvepY65DDqZGPS8YqF/64kPdwp8ECi
uRk5i3d07yGvxTH+Qc0H/mbSVbddnsP3R7dBUyEJLJcGzs46IT3WZdBPPJFF3jGcqszXjy7lc3Y2
XpCPzcF1Eu5eYBpnwCteUbr+aWA9QOn3EIoXUznAz5qU2kdyx6Dhgpt1/LNHYME6YEBVezfSY2X/
gtWP98s7werlbgN5hYMUq1YfSUez2q5Gq7dDTP2AV0fZX2w9vhBE2YIetonbMJuR8vai0k0sffl+
qBOLDg9KRX7fDoI+F62hdsyvxxpDWbuNI7FspSIsMvdzhTbKMAIzATdjxxjfDWX/QTSSj+PeQ8CU
T3iXzuyCDCHlfP3BqCvDRKBa1ogI6IY65KlgB52sLPKDiP+edNY48y0EPXDxGpxEyJ7TFFa4PSCi
I8QDOuiaLlRjgpENVHhoXE24SADrhoq7sUogzw8BaQtv84j7+6exDR3CdUEk0efO9ZgkWubUCcvK
VOpxeCRU7mgSqsKpTXsn717wQS5RRlC16vB2Oh/Dhagp9+8X7YuaPK0hdNHcBtd/1wbR781tUGgA
pDPw/QsR9LqOZ9TkwDo6JOCGGLKOj3Bqi5WHPOf1q0WsY6lepedElIj361oLwTvNXPtQla5gsN3u
cVRu4tQOGFTXlbMcsyFqgtSMWr8d4OIqys72eDdr5/yzjowivGKFuka/JR+a7Ob4vXMt0PanYrj7
Ow+/nHPUEam1IQIvdrTB/QvKa+AVnHf4BC1gdAFqQR3J7sRYNg7vcqtcZue7zBFAd1tjaYEo9Nk+
Ztv26nPg27qm9FN1TVtI2yXjsFeYEwdQmjcsWpn6H6aUz3nFeRBKGt4ZclMAiUKCxfn4v22WcAXQ
BMUMF8U8natZ5jQF5XzteAK35IqfhKx/Z4s31BYHVv2pXF+7l6Gl6havBzPqXqJGDrDyhCbCiymw
8ebH1Xjemee075bBRwB098Gtzcyk2RYX4p4OePFZqhbRujqk3GfuauTmtkFYo/l1b25XuhB1pVZR
r38J7fyeyCaaM38P6mV4NbOaUcI863w/vOFtxqQhG1bcqicOanticm0gq/pi/sscOD9RaIX4Ntho
m3TQGG9wB4jsqDbK9z1PDbVr7sMRJ+6To0f5dHQ8WxmcW6IoWT1kCmdPUb4Nd30fslM8tL08CM70
/soceO34NTijpiCqb7GLzcrtqq6rfXXAqlj8eU5l9CfSqb3usExIE8GUgRPaYb0IGq5tCrcp26QP
BB5+Rb+z2Iq6aXyqP+uiLY3ZmJAchOKxKdmM2VZQZaYsdDh77Me+kBnKBwnVhryRJFj443Ep0tGV
np0Iztmz9/Sm9PJsyCrHe7dy+qfYV/5G1p+mrrbHvPNI5MV3fi8FLeoiyMOIwVAfi9Zcmc0Zf3CN
23ysjw/FF84SyiHUio8DO6w0TH1MXI+yzrIw8+jHrsixFAZbnuiAHO2wHBa1p4rJA944m1WHq0Aa
pRJAFlc8uRpRwDEK2og78vxoLY+KPMV7E7jFNQt5UCGWd6w8gwSZ/pTJgQsGPjIbVAaXtgi8T6ZT
CzIbg0R7hqyRhpKu2C5CYOPNuxjgeRYQ4pGHc/k4PDyeY4BCMuPfJdOhDYYEYQBnm27C0Psdr1Aj
gcdHcypTnRdM/T1+QfAerUUeOvdJGD2lRfIZg/cLHGGO9olOUG7A0Aa590OBaouAKiO8vU6aZSNU
69fLqM+exJk3+M+5bupDJMS7zzdfGDfK62waDmjVLLhJAC7ZLD3E4P8cFPG5OZwO0lmMZIUqvs2t
IjX/olPVFiraDgrLt88QQqjMS3gWbBdAfET6AVpAGuhPjcfo9LeVmm2AlFAqLzA0wKfrfTXteStM
yEnzfoSU0t6vCiqm5mzjURTl8gWnTr0E+jGlpFwuHvOqWsGk0ZoIGsLTDhq9Da64mPitpIlWXWE9
4iyPAPgvg61oGEUPVfrGnKSmhKPlWclILXffUH8dmHnUAaLN3IupXOF5AP3v3NvuQckPSJa+hQLg
b5usnEwdyBXXeZZry/CSM75u64OU08UmYKJZdtRedTgQGCi16VRWbM7hK8kga6T2I0RQqYUkMZK9
mnr34gAgDHzkxFM9oSdXUlvUz19xTt5BQHOdrnYLH3RCt3U2ETbTBsvlnCOU0oi/DdlFnZfG6Tle
FXI8FudGC06nlB+mNjL3VL/MDOZzDKOY4Rl8w88DlVPzqvJ2XgywIWHMqJpduptwYVdYhIryZSlz
s9RxjSDzxA5zyhN12WKcG5evVdia92M56t8jlQiy+AmMqynBXQo4L31/kAb03reRFwnz6ReOFiPv
b/C/BSsqUikpX+Oxxk7RscjBR1PjYp8J9HFvFZykZzICZGx5blwN2Iz/qACu9CMLVynY4xbdr2v7
DuaFnklSytjh32nT0RIycv8eAxAAB7CY9fg3mFZLe0s9IxSEVgDcusW4C8dyjFgKDRCcDsTi1wJE
siS7YWFS8W0k3dw1nUePkyeXCYHHLrlhq7a6wpHvB5MnDlCeIu2JaduOIZ7rGsmwvV5papwVJdtv
fehaxnF3FFHbJqx5FrrPpufgsgiG8ed9rypZkxuV22zaKVr8yVTvdXgKkJMhiEplEMynNzUm3WZy
oYp2eEIlaaQ6Bk47QkDVayDRN4MWagOBXGV1OpjroVwermYCbYezFy7lEVOvG7lrZUV/JlEDeQhk
7PPwaBXAtHg+53UliK+dHSA4j8jkx1diCWISNu0mX3lqrTyjOLfOnMAdilLOdQGIysZWzI/Fske9
EKCSTzm85gQ2nhOQHKlR68V9jRNb+VmF9UxOscX+w1VizrHQk2hltDzOtRsKG9rbFIE/cFqyH2nw
XzD/yhheiocCKQldnbwAhJJWFmSIthpugtirDK+QX+L/0PmgmnLzZDXKW1juQlt2Rb8tWsD0oaZd
OTCwzIFw7BmHP0xNRIU4nYeOt2M/Kd6fnEn7dqMAq/wI6xnzJriTxW5yCVCRszeQJPXLVdBHj5RQ
8mnZNaqlS8zx4JVWN+EJzv+GBrv2oseEqUOio52I8nv4n9LpWIrxzPk69spXrOmUmnPAK5gGORLZ
sp9dtLsgrZJf+kcWUX9iVC2nI/w7MguZ8MyFvQ4TrGYh7tj//rJ+4IqWey/RCLpcxk8lj9UDgWyz
RJalzgBozVcd2QPh9iz9nBIUkfUFSI0Pym5s4/8ve+0+wTxBJij4BJ+5t18Zx1W1tOpZk6H+KH7s
UTlpUGiVjrZe+sxSUhOco0Qp16tmeb4KksyZ2YqbbZwgAq+WGvDhiPK2Xcg5xEzhZ00yrejIu3UA
qU2yO41BDyCgYdIk3Vaz8NPahErk2WBPVUPg/j8qHKqAiVJ/iOqdEoOQProsPWZdb9qTRzjMbFYX
K3vEPgw9wbdPaSRXR1xPWx1iXnuGxY6Pq73/n43DY+cEenh38PCqlZlGPJZ1OHynqhqaiaY/bd5a
Hm1kXKKTdG4acutHUB4Kc/xQi1FZng0R68ZOgJRL6bG0TNxncEe6iMIcuwUROTa2xbO+s5dCDGic
z2muVGs7f7/lBRRqNzXKp2LlZrN3P/4uSW2cRf7XcivcrmDCEGTABjIdUdBe7NDeP9Rznh4+FgnC
cecjCBHaTnikSzKscCQ3B54+i5+IsJYihH+Sec76PBs4GmMjldMxbUDaddi3e2PJ7BZAzB9hz5rs
VMBpEt50rSLOrF5IpYjI0KafB4BsWc0/yM//LH+MT9310dF3sdHBm9WDPWPTHNHqdoi0HM53ptbH
L7gKI8m8Ixm7kE7+ywbIbtVDqXqXCH26DdhTAgGxSE8DFnSZUe9V4p5ab5lXOojD6ZkXqT4rIHzn
DtQgFL26i+CD4ZsNp6K+hFJHVQE8NV04rlhp4RkLe6IdeI5sUKFy6uViTGODu1bgfA9J7X4SyBoS
x1Mnfmi3MhBwkdZHMFuy169j16rEEhjbFdPwBudMLaQ+4yZZRs55sDoj0tqtIUQ153T+WKZRWHGO
eJThu3fq/w5+TO7bVBqH2mo5HVfkWzp6VRG/CxgMTxelDcljHNuSpkAsNXuvtcMYWZyhw2HCTmFa
tiaD35mB+TEKRfV9d/e5b2x10fBQEpj01xnWbg8weqInvEibAnC0LHPgsSoW7+W67mCan5e37vQ+
gwqTMiYtGIIB0J3qVVpjcIeXy0XL3VnsxUkAapjOMK0jzVjXBbPOV3KAv5DCjutnmADjO8VJG26b
7auE/eQyNrxbSNAXuwSX4s1I/cKGzEmYJH0ilz/FoX5KzoO3KEjy2bX33U4I1CdUAHATSVrdVo3A
q8+EtNF9tD2ZfPxqmhzi9uJ8Af5RwH/wxp/nPlxfNFEVMd5rgHf23YcWn/Bkssd7BiHAjtpeDW9r
ztPG2DLRwbvStbR7Zp0lkYUQNV8rz2a/DMCW2IvnzrCLBKhSPLzop9/DtZb9Mu5uljUlMwnDq4JV
G6uLdn/3aLpSnvxN0afDJ7txJuvHf3QfGYsuPd17JKP0P4RODoLJeUOhRSJoz0nexoEqJrH5Oe9I
BCied0GHpJqQ0MSzKaQNYzjx2UGKaKu9n2BUIw7e1Yv60j3hzONBTpxRc5ml1vwrrtseKaYea3ec
o9Ro/eL4NUb40XYDTUYDSdisfF+qPRcSPNzCbSoBiPcwvMOxfTfQpJld8xVpOVYqhaWHwXfoWf1G
1WMoIba95rYE6Skfh72V50emvzfIMiG6HMJD1xFYFWziymQG4wr6y9YQ0C09yG540FP8AaMqOZaW
1etcAGBNzCdXH3iPzk/kfavTxOlzvSI32zGCVLewRjv9vyfKU4SKngW7PwPGFK00N3+0IyJWKXnc
v+nd1Jk7f9B6qTF4t7dvduArY6jkN32Aj0BIc5oyFj0txWjU6VPDjM8V815c+0AvYwKyD7OnRFE3
BYmzsnhq56tCBPVgrEcfPSI6cYcMNOsqjbDfR+4bEjgUR81mqtYcyr9MDo2O7ua2AgWUUvtO5Q/a
XyVKTFz4VPnCaf48cIvskl8NUopGoXjYiEyiM0ReEjgqlK7DUTnsUV9dRJwS9DGfENatmD7G43k5
iACtersc9Pyj5RCUn/2lC7kVr4MAVTEjnoy+G1TTBL5cTFZOK6M1Mvei4fFXwiXp/pmWv3F8q46A
IjMC1KTzsYd7FbkNkHnprTPnQi6vELkUl/6j6FHuudweAn9HRrsnxthDCZOolJ6iWr9TJ33SmKdI
HHK7PTrjpbMlJtPIEohZN/UNXk/PO9npF6Y0ihpjsLybRUWrWToT8IDUW/+gRV/fSvg29UUv0EX1
+hqtnrgPedTJUsuX0DV1sjoyX1sPYc5k5Pzj682GdIScU3i364uob5ZWbPcGXyEmsWxHwv3VHQnK
CarWqIjevUFuiJeIFne/aA1xgEqLA9UOfr+rfof+fipXY88pZE6hv9nkEeLCX/I/GWcbJK5Z/An6
9nUR2plQdHG0r4gQebWrIKUIg75TH51DtwG9kO3Z3GGCtq1aawgsrEk8VQUIMhkdewfGjytqw6aA
d11q484ku4nAjD9zxPo4GkPZNfZ7bn2hZlQ+movr6fJfZwhMIDvSQwdYgXq72l3ct33nedakZm7O
nHG70nyN9qd0xjgWLpaA4DdvkvOrDnANki3vZGvXwYKRbMY573eWiF99o42NhoVd9sUWJsY0Uu0B
DcS3Hwv9vu/fSAQCy1iohQJEh/Jsu0n3YKhNVdqO3ZrtLRgNb/p0us7LSHF+uhyOih5xcE9C5jdL
/4+wLDdlxkEMaWqXCwjwXoFbqfHEjgsKu2Aqc9NzrsEyiXiJUQ0ys7mnRcePnWf7wHhUQABgk8vb
nYLcDIjdp1+8mjIa9vTslRR8JZj9miFEK70eUILm84Ocs/ByUti48rfTIEyfqSjtgtqsf/rIkgEG
AbKWI0lxdpnjEoSbD/sO+WvuSb5RJ5QTIKsyEGkHigvxuKL/NGdXP7ZBExNdy6D+0ZQfmCMIsKFT
IJD3YjGq7wLN/Mve41kGfF64HXmEiDT05EN74d1sUvSt36If7w6jjQ6UaJHK1qeojXkoM1CxzSa4
0jBQNiNQM3SzRPqEEb2HwZyTp3/9hY64S2yd/r7pyD69K5wTZw5kSNpiKBaNrwP4JuEHOSWbhw3/
Ospr24VYI8zmUAA0uIuTSZzUXDMQ0DDr8V+ZuPR+fo+JMllotqgJdkGkb+GsBfYXAbvRInUXpJM9
gLLlWic0+Hag75LF4b5xdTKQkRDzGGgF4964sW13Pp78sxweCNMlRy2mWwMSFuncH/51p59yAXw/
bgigFyDsrSILysCdtPxPnakMxIrHbb2lPlf792NoHwqNHFKvkBW4P1iL5ZhV0wn4rT6VPuEO9HXv
7MOimob/L6Jh7dys3WNvrvrmxMdHJY3gO27qNm+REAv1qZc9MMrTAhBaR90Uy3ZeWjwmsfzdEh0E
FWDHc7DJETEaQl3utMHLXY+VDgJZvLD3GvFXs6xnEzly6Ei5M/RwLKoUP+JhCLEJmlgi1luNV5Jf
d+kfZvgDMagKsGFjDImI2G8MTVprDw/52gIBCgI2vEMAGbBwfWXjeOVNX6wyPMD4J7jZBzvOdSDY
EVKsLEJ/ewSFy3eItdM2dUjmDUa36EcgMfwMX3ulp736c/Dq24v1DGcbKq7sHGBay6DWqKCGx78s
mKu+JIYMIxn5COcXGsJHLOpSOXIpmPW4z3AemRDiIcheeJmkEDsFj6mViFj4eFVT/yC1gePvBRSJ
3XnZiP3Gr6xfDyYpW/mbee97O0CQprEuchdS8q4nFtqDNGVDU2War2cOQjUCYwmfQNCB7F77E40r
nH7RiBcisKyGtMU3lurka/GpgpHA+a6D9Sv2O+t02PZcRMpjbwDwWkDoDRjpz2EqizrWrYgjazo0
pBf3X3MOO5dipfypzRNuF6fVBIFBthAhVwC7AHZYNLrvzxY6ZOrwB69e7NwaQuDBcdAyGu0xpyM4
fXj7EWvxK6O2Wfc2SW5NojsY8hms2Z83pRdteFc64ozbK3DMK6qi7zFfZV4qscEWRWFsjDhbR83g
vds6JECzenYZbok8PGew/hZ5TEKDFhBwWu4ySOFtBKO5RB3aIIR9WW0d5OhAXYm704IBsECq/o+Q
MYytWAlsdnkckSA1dWyHquYaVHjtqZf2n/DdBI9LJzykLf4Z92MShqj/lQksZfY73v5pEiB8Owqx
W7KqLs6Q6haPBRcFjZWQO0JRdGfVmIL/HKneDHv0h540zv8ndqku+Fnk5DYjyMhm8Ez4CA3duwZN
botNgAAPgRkEym25agJxsOgt79noB9NIQG9mvACGU95LyZnmcqCgCQUphlxyUTBHduFy3QH6q+ff
neWYM10iuVIZ7bkSl3E82eP9PxrwJpWlKbwpyMrsuWIdArthq9eX6Z/4iLMsijvOQfTf3r5r+WFC
l6KFnQRKER/PbzA5nxBcnUXKgotLnv3dLu72CnaGqta9IIbvR2w/zeG1Nn/POrJkh2W9HZvzWFwu
UJWjOkVXL+NG14XC9R8w4XnXSlIPr5HuT5amdFSPPQp4BdyqE/BTVe0L8Le6leefW8PxC8NRAPGk
ONzR93WQaSrJaqqpk88nfJF7ti8WZJw90g7a3VJJr9vsvoH+nG41jMTxuMDISVGlFTGQz9gbG6Jr
AbQ7xXyS6RUFoWlTNyT/mLowznrJyqHrZIdlhqQ9YDb/QieAt+0QaLqV55ScmjypNVBqgstMQWe7
Y9mup4JIQ/2eT9PjF/TUgBPUJ7kDQ6Do4HvmX9f2A9Mcbm+YlOvgtWw8CmCClt8+DKQn3kus4Bsd
oUAT0i4Ekgc5KTuw4ruvs6S3rI6dD5tMqnZSYjhsuNA4Jqq7Iq8FwdMUUpwcvlC2O1sBihyXcyFp
gbRQU8yxSZtxjqwprIZsc4YGwpFBGGtArM/gcO4CabqkZTWXA4rxb+GxaJlT0sxm+lDa6X/0J2gz
gLa432iznf0ntW9goIpxjSyPH5TAnUq9ptEpxZOYNobS3IOMwmmqoFEwdpy6bgYzTzJ2JLXUtYdj
pH8ClcSW0/phuM9zPGRoxs4fqGtvplUYUnTcovWYGjCweNj9pnwWdMArSoYiEIvRnujPjaaa3Jcb
QcaSL9/ZYQ3ZzhL1lUbUmYcZ5qF44gnPJyMSY80o0CItjAyYxqYz64VXU1xozaAanHQiWCtf3JgU
XvmOZOg0F4n4gQRhe//mjL6wBKTyYuKZlNQSuRolhPPm+n9ZLG1Tvrs9le5/h5A1gynIurztoa3Q
ZT7zZJWX9pPum/Oc/G4bHEjEp4d3Nk/uVdtyVWERdkIWtykIqCSNVkgfRw8mKwBvLB3h34ado19a
obQ1zP8v3+4/JVcM3mi+BUlR4wF4zN+/dwz7ORPh5j3tD2ciCSdDPuEbIx2u7MAeVq8ko2U896FW
4srjk+ntVC0B+MmW531oVKEhKzyXcB7ebLYkhJh+ATjY+qxrW1gMrVBl4vNHH6Q9jHyj4/jsBSg6
lUfsCSW9gZ+n/AYW4RTtWP9iK0WC5KDEdUohFVvWOZr2bBVhJxSfHqEHH/AsGTrlf0JsgbFeQuUC
T48eCcnxJAyx+6m6zbgjTHVmIEdv5XoVe4k6+Xl6wmXyrxpJ8DGzbqA1KPXtjgbfBIS776ZBgeb2
ekWecI2B59uplrcV0NQntZx6pWHhXIpgntjnnorRgKjjK9NqlZ82srn56HI2Z3BdElZnKUqhqJMz
8MGQOEJU/xoxhn3CnuRSADLZg3ozEhsk+ygxXH6W11/YIYpaX07m0FJelltOCoa0wasX1krwKKao
zGPOfajACL6zdHJovFiRlt+wM5jwHLMmei7xeQSrxWsDUNzcFFfdz9/HNoPoqGPo/ELJJq5FP/gK
p0P8VIGhXhM3H8+T1u2LuEj9sku9XGNpVw2BflgG5stELS02b9H8wv+pM376EOihFEixLrEHKKYP
3LDze2Pue8GzcAai25HmFjW8Eq0q8R0BBx3fx3ujG5qsKjmR2xpmcCmEcTE7vpZVHmnAy8jwxdqu
fWqcO9NOM9783W41nRWbLcdBv4gD1+8YC74DpGpV3mYh1XZQ8LHmT3W5i0iKttp+oCKX9R96Bmhf
B8XBEo1yFarbUJxLASOg/9S98xTv8oEh9dChqiNZK7LQCtqoFPVBlU6rAXsRFjx5+pj//P9tmtb5
6Tx7cXBnZgA9Qlb6ktodqlEjjKvEdVuu6C5EDAUJzoB7TN8S0QBI9wGCwtyDN9a84PXOwwqXjy31
ZqgIFidSG1YFbckY8DS9BVEnuJJTYAA58ZLVgJvuhtOQypaxYNWoR7jczMsYEvTYH6rTFqjwvKsw
Q4fAqhWx9c7NrO8vKk4B6RZ8rYlrKQTYUfsbZ7FXDZiSRlcKf2P0uOSIzeCIKuXL9ozSKFOuRPAy
LTfkVgmkpSpE6heLIJitm2hSJ/FFXpk5Nn4UHop9XJ+jGAZSeN/wHVq4eeiGbwWXueTLOUYqtPzB
WcmZO99pRcblJwZoBr3Y+zLrdtwHu5S8I41k5l5T0jN0uzgQ85uYD/a35HuvtUBJB0oeWxfEka6Z
6p7cna1OPehQ/LWG5hqqCgETrHsouSOCIzamTrZkWu2hAIZFcD8u9PeARB/prXpFT/vHYQDcTOMm
qUGTNbUR84qZX2uLj+1nj/ow/yGji4OK8AG0hzX51Tl7XEYpxIWth++H8duwA63eWdaZcbrZUGAe
WykpTq/zfenZqtM5vUhbhQ44czVPRCQItLZKLsvZIq7z+tj80r646gIU0bSFMSSTUm1lkxzOmJfd
tw3M3sowLxIZ7PqYiM2aGXIFrXtfhD2Ac8dWskWtPNV5xRVTRZs2MSl4cxvL501UY76DIgg7ygHy
phOvaL2Hvg1P/1O2cpk8W3UW21+5HUcGFtAGYu9lqVhiXZpB7GBReWgXBAWvkiyPecR0L40jmGMu
uT7mWXjQRD3BuQyQWt+jUR3Uh7ToDr88R4WIAfAAe/803zxWyBlglZnSkwo906fo5XJnKClQ0vni
Mmmtdaozad+Pu7BPEXhDLZhAEDgij7g3BHGQQ7wLraLCh5fenG11fGSqJnuYAMDVReeAxMV3BVOz
2iZUT2fkgpBZ7Yy0Z75nARrq5o2WWw+dzYnVeguIXK9gJU5iQ9xIAJHLX7R1P/6GAWRGKKt69YMQ
5/25j2fcOOLukmaGdabOtxFAFCROeJV4t+sv736L8fXCWORVrCWBYfrz4eweSXBx5zXL0sT3h/be
dhnZ7JFY6yENhffj+2Jey1opruNYcYi047gtQRE79CZqH89ajjwx00M257LQmrtunwHYZvRUjYXi
xnKuljrfGaU4viNqhLOlUCVDQwSDLrwPk0ZElE72Gr118bsR/v9w1d/bvtMLlQACSyyOPyalctGw
m1hWLDCirSGrMGN6dyhCSBVZ2vZNaViraMytBDQKjHtmpB6pcrtjV/u0GZZCsoSVJ2c6QUYH1Oqu
N7L+Pv//WcfZa3TQPcTOJSaRw/JptktEJegXZfmpYUFaYx5KV2JXDcMDmEiPrvSEXAnO0b9IA5Im
04EBYarBtCUTamKLsSePQn9lemtPIMI1AJQd7BA+u1KX7sOPLXJ4ndCMHsqH51ltvXVd6N6PhOIJ
QEFocDdXT9nODoQauD38v6cdrrIALej4TA1rEIknkjEmFqSpD6qHezOBYYdUtt4OhoCNJMIlVrF9
RrWVnjpEYHgz/YCxRvghzG+IL5C/WxlM29wn4PHSi2oqktCp62SDfjqCijQK/Nvu3kyB0X0ue5yh
KehuLRCgZXeB90ss9Cxizpf3qYL1us5wJjdZicVoCTZnBPPWYMsZjgEPDTqrTa1hpuBE38HF6Vo9
YnHVHyYyJv1+Uwql/s9LY8yrM4ug4pvg6WCUNAp0VcDcspONlk7P8YqU7cBcMgQbJxcl/KCavyVe
8NMA8GyYZ1L3tyC8dTAX1AvwDzBLCgAc1cQVZPfQLl0FlKVP711gD5MKvZ/dTvZqqw000rUar85d
H6wxrbbnUeauhuQ9cF7V023MoUOxH4wNKZvr0PsXVS3Q1PBFAFG53ZMXVQbpCFNTajGvYqmHMw9R
q9yBcvXwGcSe3ILYEtTdlvGee9DtchrYq1HlJ2eLYtXGMetIOHefKvQLu2Nlq+tCyxYcGoGyA4Kj
g4QJli43tKk9Jx8fRnuKU9+KDCQCquAy53RGyz6QTKmjc4gghyaxbvPn13bag+pZyHulMYRm5Ls9
Jf06XiVVUDeIJp7jeOjiKoT0MWzYaQZ1eyU7cJgeT13e7dOCeJgFDF0bXXnf9bPMKRQF6sk9OISy
16eZ7UeTOsQvkPodjguUQPKUKtr32fFW2SwfUlbAZ9Fr6vQycDPaZ7gRrWHy9th0ZNLB1BahJh0F
nX1C9V5fRIKee8EdNXxpkRQ6Hf9EGqPRvew9Y2mHg+ckhe/l6/1lbodIBNuPXIpn7FCBPdY9gKgK
XYAFooBD1mcOCDSBgqo7laGbBQ09I93tsXt/SYb4cqCHLuhm5eun9HcKIpkE4JNq4TcZzYU0X+u0
5SbV/5Q9im2/KQh6/8R9NHzZz61ShkdIpPSgxM8aDq96ckuNMjMXr/LVkpxDXEzj2ZG+1d6QZvv9
JdTVLBOH7NmfaFYzEKNMM9aSWBbMoLqN4CcIUiLnCUKzp9Jprb4P5mtLsetjHJ0smyxY+24KcRPg
5ZyQ+46/TqVJJq8qqW9PbRAxGNH0UWittPWCILrIsMqfLQWnJCwBxbI+RDFURen7C0JogJE1jxuM
9KjcI71BAVV9jlbYZrBHpjXVw3PTL9gBscxfGJDxRWtVhXzUwABHIWdFomMkFwgLCyb3PatPR8jZ
Yrg6WTFcWLMYfnkbZkuTvWBR5tMUIIoL9BX5ifJa0PPc5Zoc7+0gRr3Dbx9W0GMb6q0sRRliypfz
GKycccgw0jdpRXjYmwuQ5sEu5hKw3bqe8WiPMTRofd0z4SBgrlW1t3dlXHYsfNbaUImHvI74nDZh
SsIfMr+ZUEAY3Z7tJmtYn7gIph7tNwsBiHZc5yyzXu0nsKis3mc01DZTAYxfewmPgF3i5l9Ega2D
KaqR4krOLnXgg8mLViZmGlNgoxv4kVZLX6QsJD4QoCwZGEJdIYmWZ8PF2XJlX2op91OoeV3ZXM/x
N8hadzYfEcJEyzXeb3w8P75QzRtbs6r/uvPZwsesaFtvw9R9CWGi4OH36x7XkqJnxc8YYdl6wvaA
R25BrgYcWAmcM0vocLcHU2XwPNt3JqmVs/mE6BFHGQYQkAlcmckXfD3GQugiLAIlVoEaCQCY0yFu
dUITNKbgST2zUWCWH2XZmE0HVUKNyeX9zMH2P8W0pCA0DXJrtYezlijSCB6wwnpzLI0h4hbrGpq5
PbCUE3MvzqBLC5aVLELUnrQCZeizqSAininIAOepAsbhllpBi0R6hcvChaghQ3ikE8rUtHzG3/iQ
IdVhAN5msZMLMk1TawV9Ue44bPxSMhFt9Zx0YR8ScUJ7b+DYfITrBza77D5pZijPOtYeY2nsG9JM
9xz5HIZeEXIR0fMzkrcFOPJX4KWfHei2YukIaqb1KLw0ppdu19WWJyxhvlTiiV3/AMT392393bIF
wKl2c9uTgaFIbEAONnBtdJHq1oskoNmHL6tSOb45zVMKd0Q3JCGImXPP6fsO8jpquBuGxxzJe9LX
56QfrscQX0bgu8DhPzn55B8Xk7g2woMM+javN4U3G/bEGnQAKF9wGvAdtZ2OWVYRbpxdIqZpJEa3
VGX8MmDMTG7Ll4TzpqgQpK0aV+GrkMPm/4Tf1W4VHecS+vjVfY1ikD8m07pUKGTEC05NYxc9lPSo
hvAjwxBj7HJiKX6TEzBEDunizfh6BYQiVynInuIE5+Mf2z5Kaqd2MdvdKaKuBJktfU9cbzHspGWT
sYi+tbYDagQo70WJ9SD8q2wVdfZKPAOmlqNjDAhP/bD+6XpUlA4qXelI4ZFJ/m3RNqLvUb4O0Ybl
Emtpux4oBnDwqR8tmUqgBXAtqCuuh0ymWCADGu+3Y+qEToMI4L5KMjDXwt9I2t4UPvYBosHmc4s5
E1a6MC+z6INjHQAWQEsF33bt2W3ZYU605QmrbvRYlsk+1etMD2t0nnGpyw+7CfQ8fizEsMzpDXIb
0AFCXhXha6bkzC8vLYdAbLh47on0+pLTE2jKjs5gI3k6aYA3zTuP71elc3pTG82t/3cgYVFs0va5
5YzemeurXHa5ERzuxnnlDXJ4gKFaoJbJAXw80jBQwExq8loKKJMWVJlTZQOSBfNAdklLNHfJ5HnB
dpvyjdW0hQhNl6S/uAZlEle5IG2h6/AN1EVtgWHDcBIt3v4+Jgbmz5l35520hZBM4UBipr2s4JWG
4Bta3ATTRyZ84yIFHdLZuUTc9PV9yyl1AzDntfMg+3/u6T0v6QMG1tLwCIKYAXq0V9wgeryvVX+B
Q9og5nLu8lZKza3JiJTzWK76n+i/GU9F1Qhswm32QP/aubflyaFkG5qrsZF391wV4H4TU7DSPZMs
6uRyeaQSmzx/o+WnAPYL1qcYCur66ihMd32g/Kwc1YEYg3WvHTnRxhvdgMz5MUs15qlVuZlaQU80
QlREKby0RdH7GvMJ80orIWFTsCCQmkRlgE6IL8ZhxYUKO67UY+FClH/p+J98Lg+DfefdgtwMBD3F
Mquh7+dBVoPfDVE8eHIKbkcBdFovRrerNgBK9PgjZS9mAEfGdSYY0T8htgOInAGRWXQ84eIUdwrF
mRA9d+SqsEs+uLQL+AnrCu0D6Dv87facopZAjM1ZIwte7ZBdepO8NtDj8ygXg0Ii4hi3Lhc0z4qS
TEaTZmSDfkqWxE8yZf+ynxTQOGtRzfOmK99icDMWDs/W1uK/T9Fo7DVoN1e0rMq6sOAryIIL+rJP
c2ANDXFWygkRQ+6/3N9jZI0DwC54KlsOjaqoEBWSPPCFcD+iR7ufjSAHPwnnP89Edkaw5GszaSfh
oWVspcayNCtSHpQdGQXcFIOd5t0bSKeyN2WaSSw0tPeywd61N/EaMGwkA/g9ujyPrhuhW0hbHmaI
p09g3QoWRnExK7gEl7d3RTBASgrLmqy9TW7ctIusq55i49XMI3v3fBXyPfCXVsyXAQNJGcOOGOjV
6k72zTjRKdI25dJ46HTn795OFOckYBjAyxX92i5rYx0V3FbqS2NRwA/GCm13CsclTUZqwWegLf3+
Wi0wTpAiJCpPoX0ip5egG7X9y162J7VvZJ5tUZn9C7RnhkScMN+f0UOpgrFTG/es7WNGx5v1FjKE
1Z/GBI5SvER9yXagKkj/ermx1fx98Cg4eos+Fmbaa1G7+f5pn9UbsnMMBn+K/UG2BnJA8DHl6+rv
lDuNN8eP5soH6Z1zabVWaUlh7zocBKNKgNcAuqVel+EwvPWFLOs4W/xCYnjWaP2aeXvreuClouCb
uIqTgwGRUeDQmiR6Om1FiEgo0gMIxI0jr2Rl4s4rWFqKpGTKBNp9PXT6LRcBCdSzKdeBxEe/0a9j
kzZdwvB5xBJscCgu7QfW2c3UNjuJDcHSc1sBBnWcMCR7kdycbpBtyp1BSLxCvL1NLKG2HJi5xxKR
eb2zBl6wZwOnKmWioko1z+gZokfYu+OgZzYdDFyR0c9hZBKdJBtQdBzXj5hGtyK7r+Y6vYC+fdrC
u4OU8WSqF3v97kV+MUaw7g3DieXbTxfRx6YDClxzNZ2QuFb0cmnL9KRR7FONWhYZDchUNJmnbTZ9
Tk28gexWRVv6/bXZOQcRIIIXqPhxSpFWwCDP0SoeAGSWWOiBdNbPgq9GhAc8B0Z1Wu9Zsd2Er/2g
Wk6BzdrBnOOKDWLWhVznis6JxEay/HzX8tdS8RFs8YaezAbHz8TNf0J7XMCcEZsUt09lelHVHjM9
w8+VirRSJ17hnQPWOd1sZ7dsiyKGT4smEV6lqzatESddRJlScty8TpNRCjiCu2OX4FVB5h3F0SBE
ie4stRWuUdJy7zt5EzQck6Jx42INpMm66WF8Js3owgmp2QuzzQc48XXNDGjtyMdQlX4t7MOONdu4
5xi12a8FPI3oRQMIycwwNCuaeM9vg+IZgGsUE9aK3ewuqHgC2X320vHhcMi7IHDp/PbQjiuQzRNA
kQlAPwQQn/m6ZN+HvwXndl91HcEWtlE+1oAeVM2uTyzF29kd4K11demQoHsy3caUOB5zqK8qHAWS
mW6BD2GOX6JlzdUf5w51Qne2tchNasnzfKL0MnRc0qfW63y9/bDI9yGLmp2DG/hbjwyfEXZSYaJs
3KEhnmpYy3VX/cf5XMLpivTxcRpOdaw8NmqQr+zIsitGuWniHik5xXsf1GQ/eB0xX6XeMWmLC7D5
rjKEbUMDuvLCGNxdPvQjwsGVEkYTsi4hi9Yc9ycqrde8g3d8iYf9LaZ026HpwxvnLLBruTjDuzHI
LCT9iH3fhVbe3rMjK3MOHlxK2sE/AwHayoWtGrKL+TM3LE704Nk7P8s08C09u92tLdkckTOHRrWb
Fuc7cCVlcLuT/78FIz2548V0hgIZ6TphHbeUvDdkkyjmNxrwPfgWGHL7fAWMSzGQITVEvTh5uqPV
Ez4w/qtAetPcr3i9mNvSDvy82iTvZqlNbtwkn9KQtrTK3NuQpa1w+zGG0T1W4qyQXU6DXTeyRf+I
uDcsySPs0LI4/Gic1JAlGo8U1pSs4CjLlxYPNnivP24H2uWn6IMDHINo9s6I3+nOZwHf+ty3Ms4K
eTvvLl6lzhzdcKgI8jsiTt1OUlEM5aFVXPIMGF1ykHVAO32CYnaEWEnMw9HzK2cg7gEHSDZR2HAy
PaxiuxM4WS5SeVrtlbx/RggRQdnYx0hRhr6oyVzIvSPbf+BD1QYH8en1Z9yoS8sgJrawwuCzgF20
a/QQMbk9KgQhgKLSt2c4y7X3qjpw17UC4R/rgf0lCF4zzoaoTazth3C20b9fDj7e7lrYdMW36qDy
ddyXsenCrR2j7XWsw971i4Hl01unpXr07Db1oFLSnJtAiOR603lsTtLBN3GWR8euaAJyOXZ93bgv
DQewu1sCS8b8EPs8efqx9GhHtRm9PJOczwQP8oJo5dkxc6YCAPqkti2n34yIaviFjVYaaQzz+hZQ
CWf1cJTIex9Uurc5o2C5AvgqMulX809v85ZIGbdItU3nFmHK5Kx1yy88Xk21X+q3WJJ4QFxvAwKu
G6yQAskX7PG9NSLr/FVI/NkwY9MKrut4S0dtUaEBAlNIrC/AAqRcfnqLL0n262hhCJvpDcJ7UKCs
VO024vgKRG4Ys49v8OTwQHax9vnGD3S9QjsT6nnFRFyv77jYEh8K8Vy5aLffKEsVyb+9LAcdD3pL
BRJr1L+zxXFkVEtLM28mFlxty+/U6rVXKgTsZ7eoijl2Iqy1LP5czVC5VNagBf17cnQzQ5hjvXsH
yNstWVH/4jRqAvPgNaRajXRoWdO8ez4ZbASYPlBnRcAbT3Xqh+ZiD7vt+lZn8i0TYcaRm6bSd+0M
5WT1FQJ+GuRiZGD2aeee7cUEvqJsCOzDKR2RqVtTZXASM1nE0Rpknde4XYfNgzysZTSURT2x2eSw
3TnA5FIfFGb869E3S7sYBN0sKdduN6kPYfXgUR0KofMZbGgvqLd+vkPkvqyLiieMybmLfTq2fe5M
feyxLXapcOgytLfTQ0TBY6xcWn46CUsA67bJuMvj5jFqusAclE4ugymULZ3WBFfBitztzBFYWvB7
b7+4SHxOm1ZbjJ2PbDiX6OzD+cHMyLGR084iZiCnNUQekOZzjOURebaOdu3YQB15gdy0armIzHod
Ax/0fTreF7hbp6I/c+hQnukf51h4QpqN3Ssf7P744XtxR+oOnZv1vGeaj1aBbxfvMzul4sBpJR/h
iPicdggNB0vNxudCmwHmYVs6bF9xwIHzdzuC6eakx67SJIxwDnXkZ0HLjjou3lt7RCcl5N94zOJ5
x1Zt193QlXP+SNO1mIVc/ebkkyEpX9B2cLwHOqUCkzrcpLXx6Hma9U3Y/wIh1D38vBsfQUMAFAMM
QKUs1gdoeXs3gvySNoeRyWXtqV0C1mUcmkIWM/co6nU+PEZueHp2O8P4nwMwDtQ1vUw35rJt514e
OgLyyU4wnOQFTs2riAmZn4erK6cJCOtkIqJA4f1/hpDJbWYlq1GOwdSEUxzf3TURrVaZMI7hHRoS
KpQJmdIJVD+UvnWEoiCgZd8A3o6SWeS7qkeMNO63N4sqvdPLEazD3bUVV0CFHxj58rHFb2sWYsnk
TeuZ/qG4i5JuNp37Tq48XIAsbZe1mE+1nt1prc1jNHo+Qx0oI5zUy3w/+L1geKKD+CqXXip8o9WV
uuDpj2hLk5sMkDmbnibWB67oZiFNIo0nj09upCeHJnQjvMx+OwbXcNjUY9+I+lRqLaPx/arzD4Sp
6PemQ9fc+OhFPQdmfbEoVSzl5frQF/TQkmJjFDotFXWR3uY2clbtyXDz+NfaT+XxDYuoD/eHgn4I
jXtrMPleSbxducPlCksyKbcR2ihTzVDDA2+SmocMLs4GiO6+d6X5nK8WEndPfnk2yQYDPo7z9hVR
aCKlGNzRduPylPvvecUBex72mIjVXSJUOufMff1Q2mXuNno0nFouX81EipzP2S524jHgnMndzaFC
2FXKaNocMQDzl89vNpBsGMxAkmbvBsDQRsF3ryYCDrNUcuL/C4eKM6fVQ6fRAvI9QnJzUdWRSeiF
6+Zcp+OhQGF2mORakQUVydUuLZbGi595SU2Bj4ALfPr0ztEt+AF812PUvqfZ2d77nmspojB87+xl
0C5jCwQJjX6hKchhKHJIZiszsAouUALyl76sQT565ZEr7St7wIZReqIqnb8U+vNqJw17NMDoms6U
/lxzuLRdtg1RVYirmfVZNjUd84n/B+2uhcIh5geZnjpHePfw2IAGRun9dktLoSmsOo9qLV6W5dx8
zF5txtmbV2nGYfRuv2tOykw4bgCiQglckTEEDYmggr4BRfdsPtrrLUlb6VqdCfp4B7xRE5BV2lIe
xDeotNW39cIgNN5V7hUlkc4xQw6R6xrq6v3cGqPBLjVIVfgoWpd5VN26FAskdryDKRCnmiVXU7sL
+HNwnDRtwSYnJDU94vW2OTF3kspGQKCUQKjgL+E2dizKXU/k/j2juvp6rYj9t8T9kUHUz/PxVmv8
fY5Tt9/XskwwoZ2Pj2rvNsqZW8MnOI3APAPfvgm9pYaRhPkJbXmvHAeqX4wBCdnNiGZdRI8iuC7h
bUXOWc/dT+lx4ReElLDOTYdlVN/OnWBTlC1RQACj3rwr+w7uL3tmrh6lvlN3sRxxy4JkiIqX3Zyl
V/6dfJmtZ2s6Xc3Je5jescEM/Xw2a0pPtJCbI+re59EWyAf0GA7Buba2MrSGiVe7WPWXnOq6G1Kn
919fcs4LoqGeFuZkK7kv3yEL8KVt0LO8TgXWd9ZrgBiJsknoeiPdgffTZ9i3Nck8Pwo8WriFSHu5
VssrU1U5nFLpSKOoZbOrPFlGWEIuxmctyUxbTHahpfojBM9lnJco7dLFHIBzl16SwoHxeXNkI1yT
H+C6/j9KR38WvVj8WlR2BC73GWftBF1y81rYVo1RYGP+KZKNSpfnOnAQevIPEZmVTKg/X2y6Q371
e05MAcGjX7ZC/LaBFCV677mXdJTd98UzrK/CqbzpSkDgnH9i1J7C5PxJU92VN9Z/y5kw9Btxky9D
EA5PwiRNiTVD5WtH2neo+YmJGxIrCmD2CnjHjyZCjpU9weBXsSAfDNflpQI760BSoxCpjmMApLB+
RzZeQ3xCRREjot1wpszl8pb1RO17K740C++f7EuxoUVRaCrGBqlMaYCzzVmkMv44cxEBT9uTlNAZ
GfLn//wuO7SNMMF7K7/3TVsHhFUOFNrcfvSpSrnURbJwF5FsG115deYnco2H6cqw1r1Q7+RHJeWw
uQKG48EUIZf0maoK4zwH8//fmdrwJWD2EGRUTevTLgQS/DB3TwOeb1cejRF2NSaufSU58BK7VG5Q
koW9j4Yy/28HUkI/RgEXUnut9MqCeCE+QmofkjSKn/gI18/0pSOf7O1HNd1G4h8xnlxAG/ud4YKe
OikRmKGGSAV1w3kJOXSQ+I5f7GW9eEowfQwopA9hFV+/Yw1wlUx9EGWMYPgjPstkBWqhkpyKziEC
Gw8kkVL5OomUUq00ay0y90ndtkVspPRBvNyBRY1K+UYfI+BrkB8IqDfbHWF0yLj+sPgupUVdWMvv
RD1iLX+++xvPUVihQGS0asyg9wLEoANPMenwwIdyOqOOns9QHS8zls3cEo7K8n1CG4dAuqE70tEA
qQha9YMz6swQEOWyJ+aLYrrRUX17erzh9uqpP2Vrsg91Ou1bES6VMG011dhb2+qCje7GuHURlOHW
9/hvYjMvhj50abkNnCVmrqtRNkPUTFeFbGE4dr5SVj1CVuEm9ngKHVCchUKQGbQpQn4gY+hU+cO1
mtzFjZOMWereiGlGar+uXfuApaqMdsPP6uw2OpzJ7FSFejNeoJvBqwRfQv45gTAloVvADqrKrj7Y
KZNGCbZcIDcVj7bBXOZ7dfN57sfJr9u4/KDsjMTZUwL0ei8NUV9u39jFSLXaI5O31neJmXo+DiKx
rI0EBSmTueBhT5bHrEycw9Pzo32xxNF1EJkikH2eM8qR2YpzqnAhuNiubOfRmDz2vnsaDRfPdzt2
DU+aFz7yM/VbxxuaRojKXI++bfS7n4soo5XcXv5y+bsEM5lDFccCVs9HBCmb87aFvGWZsb2dD225
PKRiQN/O0Vh9aFfrHeposggufnxYN58qk/TgNWiMUMT66/Ck1E+Am4Pdqabae3/6r2CBevtR3Y2Z
IMuAjpgZg4iHFLPecPhIQ4Az1lPeCYfvnohprUauwHJGGNQYK68e11Pa1cWP5ZIH+fyJqE+Q9AK3
woqykv5iIrBh/RObdpRHpe8qGxjMWvooxhU0O3DgXtDhjlixuemBULJvlsqSG31OKp648JyzcAUR
Q5+a309YC0fun5telGflpbsdZLFmgG7Pi+IvUW/+wt0pDNczelLLecWBw6cz4I4OW3b+s/u4AT1F
SxT0gVOapvD5X5jtUxP3Eldz24e/we/TeSGm2UOQJ8GeXoHLjOzliGHFsqtD+OmuP/5WZQnlocbW
gntkhSuipS7nUBHkLZQd2Z6yVABVYkCMl19rnh9gJJpbR0m9rHhpYBWyUBg58WSDZwWuImgOhzxY
Auxx/rk2Pctr9N6EKOv9WH98X5vwgCwC1KLGtikx6Oe0s7bzGhDO6aFxU9I5hclIz58tR+XuVr+L
JyHvM+2UMNlQtJJiCm47l2YGIUgjMWf7RbmwWxkJp6anGTR/8RGMWKgJ1tYFHP6IV5rQJlWmZwOX
iCbfTsKHfsXgKLIFz6aUUnm9g5Rz7G7878Nw55eD+ah17TgTmM+sIWZqHLZ1xrl2+T1tM9bxa9dK
BHXkDVBiJA7vev1lETai9FT7vrLHjcnEgAISqAv1b4ABM8zLovlvT4oPzzidjrQJZ8NgtQYuWDmk
XQvT7UQQQgS9QqurjwPoFSqJwBAOFudCF0XKXwUxHsjbsViNUOv8+dnMwkfuMpndHqvevywD8GSs
eAuvz4iiPUEuS0tfKkLRNe9ahOM/HiZ1v0YgiUlk+nhlC451lWNLvNsmdC9inJVTZ8HKak0E+Jt+
yx9kAOnBye4W5y9t99YhKAGe+mg9C8w6UIe9FeepiRYSY2vba9eVGVdQwbuAoan2Vu5cUEUOEqxj
qYgxb0c3BWDvEN4+cX5FQcWO0P0nzZ9kLSqLrEN8Jfp8yqp4aOIMCsdV9/OSMFVBrNUeVB16l0hn
mPwM5YSIe88/XmgAa4mLHKjM/LgXOplbzXUsqlEDKdMbUU27NtX6Ptm7rUIrCj8jvsfqELVgtuRd
4glNYPA5zksi1QEm6wAUK/Ep3jQwEw1pO84Tz4ac6bilz1BJ2gLXpeVJB1UKfvpwMxM3jG4pa0Xr
6VC3iiicDOkXKobg9DdZAsfl6iE4Bl4TOk/BZJK9B6RsV+zNOi/kOpg6UJayr9KMaleumpTDQgAA
XB/5WqcO4U70p+hCTXh3ppsyo5fkAFgTd6AKQdzzPhg9ehL/uG3dM+TnjJmF1lEAHjC7HkzopJl+
T11xvUDIro78ozCjbDFWJebXG6R51VVRz8DFYRewiOXgH0qTmcIG8i46tIHkX3Rixj4bVYm3tjoM
cum60BWZRmM+5Ra0CnDVe0E+0hLiydix3xVlMvgfeBhJqdyXiGGNnhcmoSzzO0XIFKXDDVvW0dBK
Z+gp+3erO2U5b6SXTUbPY4xwPiL1MRlW+uiPpS2c6ezAlIjyo3FJlXi0Uej1Ij1RWBLFmAp9BvGC
HtXMt4zYpoxzuWz2gFP3xtXjUddzlMxES3+/nC0O18phFQA0HnyfzByoSMY7K9azdym7HPr7A/9T
u5bM1f0IeXAdAGnMEkc3iCAdz5C0Sj96xHfIXmTfra+nv/tL9Qm0XMwli36YkhSbwUOIkP/ti9Fg
ERBj5viODVaRikD/hi5qMeORBPGAxgnOZ8St+DQbhC5UrPPhoMNGDZZjIlF+YpgIRYIJ1oy7v5qb
U1Z15FgLxYLUIXrYp5ARTJsgK3Z0ITOMoBELL+PNKMdeQL+9P3Nhdy58ydBwneqqigsmGDzKZ+2P
b0E4Timwx88ZOHTeOatyGwE42hS+Fscdk5O4h+oE3b13TwFxH8TmUIxTMdDp5H+NdW1PbeT0RHCX
LoANuPL9VIsD+Cp/FvchdFSetDxj7pw62IH2TuHnlPMxOY8stXf3pnjkc/C5ihkp2HrPqLVqZ51Y
fif95NHHmJARmQetaqEUiG2E2H3saWE+WHI5xmAlQnZeliGHfE3kTRKORdD67/7Q2Z/LW/DFhqVy
6n68hPR/W8SJOIs1m1iyqPyDCj6wT8D25gZwjqH8g9T5i1S1nGILaHJz4ZHUmdLtcb2YUxv9w3fc
hXLujsJsqEL0mtP4t20rK74hM8RzxROkyt3WjNcvfHveAi9sLDQNspHzputdCaCMpVs4bmR+zVpY
DGUhWeoR0v6sEPO2rGMHXhUumT4biwoDLjYqXUUY18JHMZKq+arE3t9AhOvs+5epA+vUSS0b0tv0
dTe57cXuZjJiGkCwZysn9hTIoxAcvAWRAXuG3bKHDKOK/iJaale0IFIJZfKVzY+foAJHslxNBxUF
g12mHSHNjdRvqja72icHABGTMPDH13JkeAE2U9Q3cQV7n0hq4B2SC4T9sXcRRGWI0QJLj9RgfUoV
t9KDF3/FakHu7srfrlUHNaojWaxKp0mqPBstPTxADazg3b4QM3+H41AogKszixIHGn+iqg8QoX7p
JqBspvNQ4wvGNzTtrQO7JvxWPxC4XOqWSEEzBsVVZviCxHfT54vipsDytNdWIluCNMndQ2pHpkHK
P874l50EKWqK0Wlfmm1JB5SITVPmeQ/muO4i5RQMk5xjJyYjVV1GciSnrYwJPthw6b0VHy2k9AIN
HACSarZC37+oJhDw7Vt5hF/Z7afPN83haLxUDSpZ0Xg5YcaFM7Uk1tA/T8ouqY5jrk2Pcy+cLsh/
SWlH00GxYPKDt2M3TcPNQJaDmskvynjVcKIvXds0P8EhGJn8hUBPteJ0qTm1dm9n/k5ntld7IPnA
N1Ii+kF1O4FwqcBhhvp/r35LOdIDusGSUKomX0WZubPT75Oqmx5wXM/+cuBaQSyLMw2NoHVoKg/r
7y1hoRCfuUrpJBHdfkZZ27FeiSaOlR3bkYykgepukA47sdMooG5bgkvxpmtcvaQzgmqPz2IWcnOO
mHzRY4YbDQo14W1YlQhs57Am975djpwcSVdh1JHDc4vegV7naLCb3L8gifPA3xj2iVSpTCpBnKHY
/xrFxev48GJmm9AAUg9GPascKhoWyOecbQQxwYtSnGP/BrfTWzzKLpD2BDbjGrR+z2kCAkUNrTna
d5O5Shdl7ZJ08GT58Ntm5npYMRo6IpazACok9kMMdo8YBxAqdTQlt65oZv0K7YD4zS1UTuuOTnZ/
kk23It57sHCoz2h4xQWQSAVnUS6BPewAcjzVMyC7PyvGmg1wlp1lgTx+J8psUEpO85vscz6uaOxF
/DJoAiO0uIXe+AMr8pW0gQRtWBjY6PvecoVuBAsNlW2iXgwwxnZc3+ODu44vKwZ6HfTchK2PQpjD
DVTroSeSYFshzyLvza36hXP9S2r5XoLZf5p7z0XexTXvp2MJu6aIGoXH22GPrRJyuRyRm/qRNUa5
+sjZiMSv0BxO98lRofAXA/JgsYMwD7go1jdoPr2uVsSgR7ti2gzmcB7FRgrJGW2j0DPd0+qq+ebH
dLXk5Xjf41Tdb2q7CjAzOMIbEuB9K/kxcXIbtfBwjWBRmf78Hzd54WfoIAQkn0Iqd1lVgWZxNWjr
Q1vwzHH3VWeZOkprRIFMwAho+6NRTsDNcmy1Q4tKwd5Flz04g0wj8fNV6OVSZB8uw2mMtcEw/9u3
O5POYXgOqSymzBF0o4i+Nv3EKCC1AKfrBV5GCuVnSomkC/qeEG8duFi6QyBBidlA3zW8XJzFBz5R
y/eiqbf2fsPgwN1OpQvk2Q0Ya6aCnbo4jm7ts5zwLQxmfenQoZtEI2iHsu6xEBjhmQ3okV5O/8Re
6/XBf/KQOT9xeymp8zPe1po0VHMU9VRr8hMrgTYeA4jPkYnm0NY/P13k2n0xmI8yxoELmEuSy0FV
dbYhH0ZZ3QcX/UJ6Yf8UQw+8bhCMzrrGn4yZAvidhwiISnRKr8X0pIN8lEq/wOJKdN775Foq+Qz/
47DCinYmPOGEiS7m8wVs9QYnBqPdLKQfpeSO0871bXI1GXEhoJn/v7s1hNFEepzOqse43Sm+VY6Q
FZbwLSY4LCqn+umB5HI07vFR8lDrImUpFQ2aOhOb7gAbHGAfEtkRqTuECIs3t6sWMB+G9z7PORJ+
9UAOV6Wuzdn7u1RQnlGXv8zWxpK9C/WcVVNG6BxOayoW8IOwqxKtwgS2BZgDprUl8T8e3YBraLRN
5bxGOHXeIxIS27LhShk9oU+YKcKE//iI+DNQIaXmx6BhcTnBEXp/ZY9LJfLxCd8652VwwhyfClw8
i7Jy35+KYww4F+FifcBDR4M/0mibOm4LA2e1UzqSqUauxEylneLIsnSLCx2wTUyelt5ZDYY4YCyw
8+v0PXzfcFsQ09NvGR4FRT3bSVPELVxSH0fByilHEIIR8SQ9hv4BX6QijdZKv/5J2skrNUsTno6+
9rBYI9ivVl905rf0jHS6AerpdMLA/JNiHSKk2TiOw5Xeb4zrXfOrjHQvwDuUJDJcSfEWX2LM+UEr
8aI+yktmfYDOrhtdxZUUDEBKcXwGcN0KYla3kqC/MOxYKj2jIhrqizvK2dJWgzkUOoQBPo0QoeAk
bULCnsDhN1cbBuE1fKufdYiDKgPWP0YcFU35ANdEylmeBhOTaa/DZXmCAdEmCnyWc9RW/a9A2VN9
owcTG5SEDloguJI4rJtvfNtN7pbTdMAG6SPyEwraj6qmNwGXxU57KnXF1pf72fL+zgcak2w+b+8c
yNRjCcQET7aa6/TtecSjQeDBF3drOprctdMfozKLrk7jBQ5N/e4fgKgP5CBr6zRNyBc5q61RZsEJ
B/X2Eb0mtADK7ziRI92QuapmXQNSdlimZQrdEHDiVAPzEeDpNrqiV58yugBKDUEsKmSewavBK3mY
mJlwZkkKObbq53LiLo92VfuGL3TeqSPPsWzjIfZ8rNU2r5u0S8xl2vwCvyFe0YQg9pXsK62Z4T6e
loA6RHFXGBVIee0YdRqPerf32Ue+ipHay5HfUclb1lqaLbk7SKN9RMNzf8gIE0CnLJ50dMhMcWKw
56pYiQIIhRQGCO9RHI/WLFbBJ2JT+r/NxXQJLxbvbNFyn1/n2Oa2kGQ0fbzmuUlX/vh3QLblWGof
umWSGYRFg267MOZSwfOaXuv64ikG+iREYprXB0hEeSRX9jradtvd4ClCn31VXc7elC21acl9/9h6
3g4iY0DRSfN3nTv4tKRR63MfEcc2tSRNB7aEEbWm78utPBU+uE8juDilEldHqvT5uz+5x85JFPD+
rnNwTwZtgice4dlMVBZ4EB3fdRyppCr5BAiANS7XtwJAKJrovETZcucqRic+ZdoL6+65tGjGbCcP
pCN3M6ihAHwOeal64a1VAhiuDc1JWZ3oQmrDVnsWAbj1IbwFBhwm/3CxhjXtVmrBa+y/bRuRnRpt
JAQ++RLiGL1OOqY3PKTSLn/o+FISJeAPcV7ZC7UZLITvZLoKXcMUOsEBMnYWyzTNAnmzJHPC9bl1
b533YvTGR8xQ64oVCwplYBVwk71xswcXYg7yQQQuSEOt8kD52c9enZR8+S4eTBfBYDs/jTtf0r2V
A9dn8tyiZjIlaiych3FIAd2X5FnZ08yXLgnyo/fEXPEU5csoZCzuNI512czUoPfVJNWjicgCwo8h
47oa4Xn6pVS+p9qjqRNl724Z7MZnL/a5JPl9rDteKlkHuBfUBFDz+iRdmR7mcVdT1XZmldDTH3Pn
O+dgn09qoE00wp4AwcA7lLLKWB3/A/2pvKmkiLv1fQscJ0tCPtq6lgPFfYidAzFIcjeor1fuLjAz
GYSwK8A8CSYpzmvKy2OQZHTV8RGr0k7CPiZnRADW8w8E1Mx+t6R0vrX9SjPSfjlXglJW6oIO9pIy
4kWy4tPSRxlRD1Tg2MqJKFvt++VOjXWcRnsUv8OK3ievskp58vG5E4EgqVJGuDfJHtZn58bqyLKr
xFYuG4l2fNyNd180ZgCGNlIz11520SemDoI/xOQyAl1NPXgGbaJyDg6AiEW6h4Be1IqNB3Xxl1kY
/YCdPe6xV2hDYdcXrvfRtVZkNFwGMidW+SGWqHmwVEjfzrVPT0WnnGbkU+j2rcBU/KNfVG1G9oUO
w1CRJUlUsCbvfh4ixsJfNL/FEQff1oe6Eipv4asLjKwGpK/qwNQdMPNHtlAFa4keeHMPDNk4rY9X
SagG86ROMRUx3XCnCxRiIzAQqROTNQ+xAT/ukO3rjyXYC3/AcM6DLqwnofav2As6DlNVQu4tf49I
KjBGa+nedkcFdCzSK51+bKikjsQd4FOKrAJ9ani+cov/A5J0dqDJOW31p8lgCh7gf58r2GFLRILa
jj0TBjj9D60GmtxiXe4FDErq6rmJgcMsFoS/kxs7w8j0ugP7MXv67RtFsVAYLAIYKO4ndN2t4gNj
m3D8o/x3rq4DYV8OhHsHLT01lzKDbr8BNL9K5hYFDezJ/S44ijvO6sB4Zg0dUQuED7FBLucyjsmH
Ayhco763oTXe8vIv/Suol7kMkSwDGrclu6b/KWboIoZvxu0GC1cYyY4aLp1DxOkvAIPNIpXLBrmZ
L1w89eT4x2e32hT7lJssteieWdf4BLP+RTzLZCTZSH/5ZRPqNCj4LIPU+W2m0XtAh/P3aCa0fqM4
zKDMY/cRuyJwyNJcYj70HU5yAdew4WUMtDDYPTvcmkdXeRgr/8kSCSLhAfIru4FfWUmqng8smFNS
G04wJTEsZNTFGWKcl+Pb6rg81jPZgD3kdMd4r5f919UuI7biDewiI2y7rf00Ffmb+mled4/v/moG
frzH8At8y+BiNt6PjKYa/fyEhepGjhMtFdFGWWx0i2gyycWOasi7CVZmcVnLHnGJyolwjORKolDe
diKnb/kpDde/RrQaJE/8D/gElLWsR5+xZlDMleICV4gOxTF44TJCYnEsuSEP6kr19daIW+ebBKEg
IizFlJFDJvr4MmcWYdcjVT8ptGkWfCmKhx0VZIz4i4NPlY0cqIuGhVYR7NI6qBd6iMUe4sNxis4U
v+9tNnIGjt2yiUuwqRg3VYsWSrGtA2Tm4pg0oto75kpxU8JFfePg+3z64r7PFLmHNye4ojTib9EB
M3iXooQs8Qdv9O0J+u55DQqzooMx16ruxeXrajtY70u9+af+/eI0RnXwHHu+pmclW220BZrhku37
0pKMFyJ0yLiDJE/ofIL6unDTuAbyw2tjZWkeRVhguV4fBfO6v+RUtDABOu3LV1spFujbd8z2vId/
K9sgK22FZmMLn3f74Vv35eFWf/S5fBhyHiUOSpHmvtZr7KY2gSujX6DX6W8lWZ9uXs42UlOWHIBZ
SfUoEqeFkQUuNBT2BzgPeKFbU3SUAla8OlAysSXf42F1iskpuoVm3GKoK+wvz6vbih2iAGUF9SSC
EvQo1g11LJQdAi1BXctAcO0JB+dmo8W9/nqPcqnxsPBlNXamif5YXXU+ZF36HtwXGyQ+fToTVTxX
47RjZZ/nhAfphNx9Sequs6MdP3192iyGqdDfMziJT9ERm1/xdBIwRgS+VDCiYI6p4NlRh2WHvcTS
jQ00ETG1arvWC5kY4kNy13t5RAlq2yRN5CIYTcawg2z2TUI6xH2mDrhaCuAElBrEmg+dIVwpujiK
uO0ZzfLOxmY0W/cAttxkcFvCzvLsAz8SkZ3UbyiCHi6OfH5ANrW/3YVE7OkGBHLwI1rLTDCJ3/5C
pXcFnSb2eQdUVOArLaPZDM9+jCHyhpDSrr6DyUqY/ugSZRmKePkIpf8Q+qlwOPZ90mz5PuJkXFMn
qh4FxG6NyH2QIM2gAgqP5A3tEkbOdoBqhJx16G8U3+wedyOqpa8xTrz+VntBTBUOJLxJGP3htfYb
5Bx0bR+IT357Rx5Cgh2xboEKPKZpMnKk69q/8h6TWdBuD0Eo//9izZHuU0sUAkv2bpSU1zx2RWbf
vyYDJ85O+WxZgf/On97Ua0e0sMdy9wBOL3oPZHkucK7eMeR/008qlNavGTsQQbnYfhJE3sYLHqdS
KgTa0vKe8hjLqb5krBONCyEva1OC+Temg0/9n5OOPkFbcp9QaPNom8eFEEGKbS7/X1PS7aRvjo/C
XFue7cZ3ii11lPWw+ybQF2ig48ogizpJmaKznWaeuKYsssEGlrmF0u91dQvK2y7IGz1/DMtmMYK2
2J2756mDO3wnyWWQcOKQcy6TbLjhLKSJq8hlQFH3heI+KPdNU2A0mjJ5C1lhTi3EP7C6rKgXySgu
EL5hSiWrP91ZrCCA+05yQVipvdLK1weXoia1Iz9hN6eKSFXK4n01PpbCWcB4lnIIScYQwg1tMs1B
xJQZV9g84Apv997T19WNg1V9v2CyoZ4Yalz5hb48xFat6kG4f5qEMFfOcDxvd6CUEc48rB0cS1i6
HNG2RyRtolZmoqjHnFNAuNLm2MdsXaLyhzq3FlULerSMCgjmV4kNh0BYQDk5X0OYbGCPX8evnRnJ
bC/GQWXvt9A7KPpvh8e+ng1cZu8o3+GCHTuYBd7d/9yGhu1TFgJvC+8OPiaTQkn+RsZlqUbftvky
5XYui8VZAK2asY/Viw/0lh+7eMFDTnyhW7JRgkMmgHyq8joLkXzRA24QsbM0haIybadbW5qduSd1
tJiw+dPaf7XdDMktXdWbs+jn4dCaMrS68ChwtgBTL2wG7nalePH8vuWYqUvg1xPof7IVNygIWN0Q
1//X9AEh0mG/UbqS+nhvbESgaCYu1S1NxFea9DcErWfALwA0SD181VnFNetpmJCD2W3Ha1NVP8nN
hR38s8ufEe4h1i0nM9igBJSKPG5LReoKEVD+bA4febB8qi4cBq/Wx4naO3rlWebnMv51Dua54j/u
JHVv7qRb29Yf3r/ts955T30uJPXBAKf/1qqmACS8D4VeR3BDZEM3onDD9FL71weiuuNXyiV6Mrk6
4NTtFcO+JkVF4vQBXOJdWIsNPwb9OaaNv8piAw7RGwZoxmiftQhcGqy0G49S7Le+T8h43s6mk31I
76adQO1d6O+q4VxjBp9MMnpEL2YJ+Oi+78jSo65Pt4L5KhUcDgVXa9ilceB3+S20ip4OQ+kfMDmP
FRrFVfintJ3Vy3sOPzFyncm7IUoOP81ov5fSWuRlpCoZob4A9xPupL4gKr7+ghHMMduFRUWObjWn
YwWSzD6iEAoIqetux4ZZUt+hAA3s+q/SZURZ7PDc1Xukn2MWv3iutIe+NsEWYGNi+dP6X4lWLJXV
MFmUTznWd9tZKDsCVQu5hOT7S/8W6B2GfwVvAK1CaR+7Qy/+ETJSBWLxZ8BhsfTnOPQqFXPINacr
kSmuQUWh+KlVh/HCAwQvjFSf8sS7An7KSHyaKj13CPcHrKbOF8Hgd0WvfRpBuKxCRcyDIFf7PR/Q
SOJygmQMOWgfvcCd8N+YhziaUkkr1ACpyoIroknOgMy2d8ct8MoqqW62UVZXCGrea11p4l9ckzo2
mJ+Ecq8yKmsuquouhVEahm2oc/aRFoyR07LrmLwORyQvD+xRwMeD7c0z7KxVxrgY4fHrJFewxpY+
0043udi4SoT1dQjfXsX1JoRl8HszlEHWxJdi1+Bp4VvEZ5AC//t9hrxw+KP6aW3hsx6nhhCVv7A3
dXHeVKOWs/B24kfh1eEG0rix+0G4lZ9Zgh+mhOtPwmEXfCRgSI55+uMG0UeJZzVHuR7XKVmjqd4r
ne3cR3+5cIX4czzx9hwUsyUHn1bUSb5u3sq038buA14xctxH/54DiMQzCygP6P9UXETNmSN1W3Mw
SBqYPrdKIU7Cpv3h23Bcfg7RBlPxq/DmAvK1CsotOKaoXfwNAaalpmkH6PknyWZGrhKJkvDV8st0
xF0sg+zmpRMTA7Lljqa6C+5tMqNpXdrvByyXatsfG+gCYmMyQAPaidQjXFlFoKI6dy6yLOkbBZmD
3ACjqxxyiv91DLCuAYr6NktYBlP+9jiQuRZyGYMAeCBuFvsrk03+RxQImDBuXKnbRYDDPi/1dCuF
OijQZWxk8LaF1dn9zWxHvQvyMiipfKK4mz6ImKRk+hec6ueASV9cGmWunqLi5D5j+3RzwB/PzSMF
WQ0ZzBoARDvsgJYoTPm9YCrQw6PdMKyM26D5weDICHBNuonewAExRo7+fO0QEzIQmcYQQL1LmFBu
yguk/hmyhxun87J99d4T94CHuODvfOApzwix5lQiA4oiY2o4e9vLo4YRVR20e4kuNWyw6s6DeQHa
uouiV3d8jJfFYCq7k5+Y6wuYbHqefXNUz7y5cDE4CXTrem2cEefTSUD2kIf3Zliix5IkqbmLOxmr
0VVG8avLGlx9kHpK1casJAdPMWvlxqcBBSADKA8qunvglsYoruLKbNwQGTh8aNFq3TQYnOS/bn4X
GIkUfkC8WCYvQiG2lrAFTlRRtIHQGC6J9nQO/S8i38Hnr6TlPLP/BT12GBrS4fghUHB4AliDsz7N
ZWMQzznqenY3Oy+th/TF7rLn1Y52sNyGtnAP9XgFxS9LoNLknDX8WD2Vk7r52q7d2sQe/bJe5QKY
i3I+LbUkwXka69gfnKTEDVBtvFxA4HHCzIwAsQZ45O6ofmGK1WUXqRxud5WTLovPBRdcHJudSTda
xiEW53+2bCzWTGWwx66Z220kwu5jTTy6i6n1xd8A4S/f6XA6uvrZNI9u7a8fQrWJ+cPWCMyZdeSv
YCl2uDjgEG3txgdfQRxrzZYrxzgPFtGbhCJKSWjX91ugPt+h6boW8Suc90KZZkO/4y0NRlo9EfVx
u/2+K/6+atUBfx7/36YjWHG26V43r6WhDiuHmI3MspDVbccx8A8/ejU3cIFGhI/HTPPYrMjS1+bO
zMxk3S6b0lYrybafipuYDYITcRrs8BR046xTbPnuuo5IxeEE4YgdPqXjg+23CbofebZcSv31zD6c
IbXOTmwW+Mv9LWSVbr13NoFdqd6TSiBDVWn+h5IvHs8BFfHiW086dVJZOdy+h+uV/YEl5IQWdajD
qy2j19BilD7xAdqI8Kc22GB4Cp6m5PObRju9pQo5M/RCx71YOzE0D2RqgkB4GuNl4uUYYey0wBij
IXpqiYygN08Pg1Yb3R0mVl7FqqBSzwUrzIx4hcFjjlEv3fPb1xRTJy4JBmXKPkiG9nBkYM/oW1qy
La5Yfx4nzu5BpurH+322ewygVf4KGwz76jhwE5buTxOEFWvfY0fITfcORewq/pQoXkYrfn8CW6ge
dDaUHWEcVK1QIcoIUKEKbenTZifc5L1iomUkmWOY9+TD/womhyz630EJaf0k3r0vqGKT++rin+xD
vgi1GwOkWbat5zFp9EkOY5NR3VtUPnTHfikPiMKwpaS+EK5UGib9NRDWk5mL2Prc9IpnZ45Dklpo
AwtC5uYpULCuATfknqGIBsvNvKfZ19rgdFMsrYblsv6H4a4rz+kM4hoJpaojcj53PGK8cBRVGArl
AXwNToevMj+Y/7LBFNczOtychaS1VhO+h4XFD/STNMaP2CqI2j+tLgaPSRpvLTY8aS+FupQS5OAo
VaejHgjlypHnEYw1+Mlda0DmgJCdYeBsruJy/s8Mo210tELVBUpNEusEuVNbyI6MyPEjnu6odOt/
1rTbBXy77jHOTLsrgMcZqkCe4qDJVkRKTLupZab1Q+0bApFhARyLQjY1r3BuEQ0Soop4hhxUC9ws
3MTCYzzSH+CNTGwDT11mbDR5SxT0KDIr2t1blap7BFD0TWXUwlrp8Y+H7oyuUR1qYeXLx/tZ/wH8
xLRfzJ6vrezNfasSv9KwokRAPSrKlAJKXPhwbvHNYR287cXkpp4FYJuONBuvm+33ZPfGs/rb61O7
QSAAxiSt7Sser08qD3I1Kpzvjp3sDT37FO1NRNLJjmzK0zliSXRjbgBjef81Xu2+IrLXy18YTiup
RFCMPXOkHfzmz53Mp7sUVxrkp1KgvXROX+d7DLrlbBU6dIojSlvRdOnirmZby8MUXJlmo0iNLU/b
zrJa9HThKVhzQQAgLhHHhUc3KAnZsqkTrGkvccBerKaTJuJXMt3wZSvrd5V2QEojzS1Bb4fjVExy
+t+CcaHE7FG1QVTcmTFhMEA1q+RXVDNpSbPah8TIFQoDzPE375GRlRXPoQpLEbJqwnwVS8Gf6TWS
EmBrhwCZPb+g1XZdeqg/PQddUcx0iAmNfk8t08LXdsab9B6jGSnZ9JqsLw1aFii1yvCnxXABfA8B
NNKiNzqLG6oPe0ZCJsX/fC/h1zcvF3d66Q4zrv/pYuaq2Kd1oGsyCxz0ZWiQuIdfYjRA1sDrntYJ
WR9ZBlaxxu0oPq1qTqyE4Z58IKinYLOVVJ5K1yIf7RZXlPJHzEa5qPmSQ3Iu2pdG3bmeDJnYD+wa
SH20tuA98mRY1uVqSwsYKkeGyUp+YHfc3+b+POXtB+WFaXavYftuupSaautdPWaO+rw24quz3k9k
QM0OEy5WsZZpRlNjos7BytmsPuaASSpFcjBBMt482BGyKrqKGZk5WfrAxNIiMvikbLIU1pR2Mz/u
2jsaFcfb7Zn1PAfgHLuFzktwMVhbaIfIM4Cox9ck8SgO6pgkxYjGu1WWtQV8aCjnIm28rSv0ABD+
uHHTUUB1oyxK15c1FlxlXeCY6HVs40Hd64A8rMrujKFil0T7jX1D8gbKvEf/SdIXxKSQLiurG0fq
fbCkqvHQGvZ3W2VbEbLcw0FpXaV2t2Hx1gOLiHvWc7LMK2IJL84Bjr4pKMiYCmsUJnNjTV42ZlJh
7IjWtEc5SyvjuNi190/ynSN2+HYYFnAMkSTUICCYCaUd8dvMQ7FdDkjl338PdYsy9H64ylrFpL+6
BjrBZWpc9XT7MM4C/lbqNU6UxLV/kd23FXiCHmU8aSBGiZBkn3diBm4YBdrT1qEMo2QgYebQgiZn
H/gx5kLVmptZTgCHRBsIEu+p3uXhDl3FTsTnlLZFs36VZw9s4Dce5fikZC/1hfy9i+quGCTvLAQ0
4Igx4TQxdErJpknMhhIRE1oVcnPPftvBuDKQ41sMGjnbJyYWLOvn+g88mEUfeUITWHvDIUsqIdJA
13HdIeN9/xCFNKRyAeGmdySEcI/gpPrHrkjsL+tOUgDd7DPPB5eNESTZAHGxnEPVnrU9kMEJ1Pme
3R9Zau3fWSUL0dGC5UqN3bdTy/cDzaphcrXM6q6H/mqF6kGy8p9WWGbqxPHU61dC+aqsEvyo2p6B
dF58MZcaCXhYgRbCd/DsdmGZmmCrgc/LEWkXx5yi79tJn2qvC3hGMnnhiIZd7dZxsW1mRJopbwnU
qJqN4AwBP5fAjN+Jc/zk+l0Dqt36giRu1IT4NEgRtxaqWX3/BLFm8xMp3iuhyl/XMKCoD5+Gsk4L
uScgeibmyOa02tdBD0Z1IsLtZu9KiS5e+BTv04am60nsDz2g3aet9OBZ/lxk7h3E8srMbFpG9uKF
kk15HoE5FNYhRFDKmoLMCRKImJE4uC6pBpdGL2i/fL4mS6qpnvsNm2ZWl+Q8jgK18BEYnZRZMFWw
vb7VE21x0VepocTVhcRbFHZU7sqC8j+epZwdJesXxmrS/m3yvO3Vz6scdow7ME9m13MFdRLaCxtH
4P8vXTu96A6JgD09oZovXdEesWVxX+7/rNEBBihEwe0ziaqrY56Z8C66nL3/Ry9r0DWBz5OlSb0k
X0/PXj277LEpzuQq19iU7TDISUuciKCCbvpf9UDSUgYrnDKwmPV/na9SxpTUIbTYHYZqoQjj/1dD
cnx5PJn1axUTQllv8HBQQp5OyFGtH/9+fEsFCpuNnD4j3tF6Vc1NSdGwkXmCuH2FJESL0yPSVrNr
6ClCjP8h2TigwCMdmMRvIV6NJEfodTv0NVHZ+eFgYep4t32xw4ZBRX3JUQpl5JYn38DN+VD0g6ul
UMgeCSRkdv7xu+cslMDNLr/VgyRxuNAhG2Y5EVeyLgBwQFz41XEWFPQYoBPkpXYjqOSwMcpS39aa
PRSM/DxNRb/TkYCVKDJL674ykXwCubpmLVK64mY9Zw3Qhqi3Jhwm04jML0IHcX/+ccDSMwi2v/Jw
3GAzUOu/+v7vqOnXh6FY5njt4rbynbGHg681GCdhLOeeEZJWmdI4rK8HO8B2z5/0QY1O0JojQ0Ra
MmaT6euo9PX/ViDtKKvMWjnX37uDMjSRUDGKs/Jc25Wn+PeUYtwNL1VQq4YB9C50ryExCmC6smIh
J6XIbhJLz0arpYtljh41SF9QPo/3Waj+qT5Py47nET1RJDrMwdp2w+AeNznLUutu1w8DdAY44U0q
1fdbnzeZ0QfXfW2w1grgAVKtsUdXenXIf9fn1ZoraDjeFzuKgxlzahx8QKWvERO0uOgscvJ+Jolv
lDJCdRVfDiHJrynIKF1K6bhZNsNas8vtLwKIpNf8eW6HqCu7liI8FSDL0cuSXpHHkpXTG4m17NjO
psNfsCaLWS1rF95W8Bol0fKX5j5O2u2MkzznpcusTvXbP72TCxLg/5IZCgwX5ujZKKUt9wj2abib
9b3RmyKR9GGJR75FSvKJPsWTsvB6OKXNun3sXeJtbAwHzI6r+S1NprWQ6CBCYPIP0u6uUIB7qjGo
efz7/sIr4qN8EbxMz4T8NBaik4QUSVQsDqsKQgC8zQZfm4H9qfLpMCoAJe3siQEpqdypHMWcaHo0
be7F5sqnmvbfJORJYmIDfK/W7qECUTUCWve4L4vDtZcrvz3L8gHEEHlxO/YC4iY+gvl/nTINqv9U
avvdv32sREUMIf2GJNk7kyrilMSD+1+L3vpMrHcXf/f+fzRxK/U3GpjhM7WGd1n0gkJCJSkv7PE2
p7uFZ/wHaUWsTeCV2F+WLD1emkAI7wLeFqoEF3YKC8Rl6+0UWECkY2gKgL6REMYLB/1t7oB7RBlM
JUK2r3Z4Wt2KQ8eJHe14cs4B8P/+Eb5LukVAn8Ff4e06I1phhkqlTi7nQcjf4pGQctmEWaNCSMqb
NVOhQNWVUmfjFiLnPnv0L6a+MqSX4JPGN4t6kbp3zMU2d08fKe0qpnKfxIIhg2tV/ol7CxViI+V2
Yhtro0BV9lG1U9AWGxPaMbxLwZs8V4JkDNd8I1qucQhDXLUN3lesH3YYm2kmaOhOYatOapGKg2Ch
ZEB6L29d25ZxFdzQU5Qr9QkXUCJ5+6PSvb1yZ/4wDahN6huC/HHF15TtzRgBc0CHdpaBcukZ4vvD
VakPGQySwNqPVq1y7qiH6ZVYAXzIpVTqhmkvonj/fZ35M1ZAK9JrYs+1zpcLK2WoArKYeF7vzg/9
5b591a7Cm7HHTzAbAZuT5WZDwTGEn3b1fv2U9nBYNWyKTVgLR8q6VPtt8lTijyDtc721ylpKjGch
e70VEAbrUMi5ZjaBZYhgEdBZMtpr+xzmHgseyIegVFebyBqkEyytLrP7NJ5g7X2iZA74SCKWweSl
xocQh2slI86cSw16OEPcsbUOHxGceTyISbHcHc80ON9WSkneiMIwMYRWzq9hICOSsUdH/jpvTTli
1xHYivDGULA6lLtpuTY0Pa1pSd64fT7gZ7OuITi+6e310qBRmKijpDxiNE0f1JL/h4UVprDQqbEB
c+t6b9AHFPkV8JoPLNUdyFcI2C+jkTFbuoCvMeajaBRU4XQdbzupE8qMYo+49aeZZgzKky4P9ZQW
rWOBppKIYe2mpvIPjdc31D+onrmdQ5KqdGKJJSBGw/PLFSTgKv9QXLr+tPGnyg+mcmEkGavQqGmN
abfhv/Ny7jXeSC0GTS19XEYlzzN8wTIGEzxxyFtNLNf6BN/7tvqCFWYf6F81P1gHjykMFZAvHRB7
UliwJfi7wt9EmFluKiDOLULcGBj842bBkY576mfCQziCVRnUDAd+ZbWR5d9rIANEHs/BlFjkwKIE
/9kSRbAbfHV4vPzHdGY+sFplYnC0HxIPcpBwP8Fj8iJifHufL4ZpdQKCDgvd9WLh2mRymR2g6oCA
7m5m6scfuKlExdap4rAxHfPZc6Ii5YMwu7xATO9FDiaIIs7KjxYs7vapQRzQ71j8JLMEyZWMOqZ1
rsZNVNO/J76pw3S+8XsQP+wXyDZERPbItzTY9ZrQR0iexqHWlWx0tYSj+dKAKWhMFQNbD5txv5pC
cB5b/fmBzFxdKOBACXgee3SMLBeWY1WBdLmcZdtpoU/3hw/5ZrZcBxOANqXDRFwD7tU2DCQL+QTP
2Fc8r2y3vg+aD5RR3fVv7wK5pW/WIrDr4g8Vc+B0PlJ+YApeBKGYVErYjh8KlHKzz4wkpkQWPICJ
OAitNeGbcW3gxOd4fYawSroLCz9lWHaE+Wv84OipJuNeaPwc4E1bbSFsecQVgWrjjmnUD61CSrsx
pm24M4/QOe4Z4MMnYbwSuKBdCXA+xvTWkjEsybyVS7lsCboBsknAkF3YGZhjkOplARxkRsbfX1vI
Ro/UMVGbnmtH1WzYM6LEaMqQ/zLEg/7QzWStaT+UrHRNcFgQ7LzeeDbIRcGxgqH9ucFKjLXuJ7o8
ke30i77ISPotgys6ld+aMBwrfZ5n3VVt9c4ZKZ6FgCBthPm2jXAyetBWMKYf531+nYcF0wsgWj0L
5URQRSBQShQktj/i++ptdhXxXvMQynfXKBTr/Qu+DNjWzoE7FX89pun41rYBFqvS9v93XSNJfk9K
ApW6aINyrMVA7ujUSTGpXmtdUVWYJCTamVGO2xJny548IT2kcFLHjr6AmyGdqzQvzpydhD56joGj
Kfnd8R6PWTEdUwtFM+v3zgWfuEYVyExctnAaF84BCKyanOeKVgRxMRdE9B7ZQY5q6mTkpOSoVGAi
BgNhczr7oOUL4Kuu5mJO1tgNLaDnxxQxLVgn5T3XTAZsCYRbPLxIOlG1ZZLOK825VrhZ00CvF1q2
j6k1ag7F/31xTGZayy7pn6gmz1VeVFe5pLOS2FojdW71111icELYF1y6VSxJ77J1RfGmKPaZi3J+
1pAlBLBRis+KO6zYKKH/aNd1vzRIMZNPjKOEszp0KJzEsqq0knX/OPtNpLxkmBCQs67fyh3oSMpG
Z09iYKQmWpbopAZh3wnW0WX7VeLFPHL3uK2NThHvKX5vhbfD+O0leQI1/UGZEdCoe2kyNdaorPNN
U4dIg7GoNa0rGzvcAMqMGrABdRBW7irgqARTepBDIQYTiS6gMcn8LgWHn1Zg5VOftoumpnXYVPL3
B3vO5tjHlLWCXXtC1uyGkcSaeOJwV2otIfxqInI4Bom5YVXIklyWKQPqMy+DXMtBkudh5aC51S4V
YiRsWqcrmoDSpulUrLl0pUdn0qvrfsJY0VbfYF0MEEYIebQEcjrk3SsOJPax3fnnTtWkPcD/3O38
WffJXGm7V/DUarK8K6VyGYy/54zv6fx1/EFmEk3CuGS0eHC4JcWxEP3c+qMSZpvcXnz5231d25uM
xGMI5ZBzZQ2T15hiV8ZyqcPX0gcqX5T24+6LYyxsfaMMjui3KXq1QKpPj/gfNPanMSoYMn+g/uHL
e6P6hLaPawd+tWnHguZttM/VVZi34KeQyiAcCFA/8t4Me+K29GEUBlbY/hpG9HAytLFqicVovyhb
mJqocCKyF6zNsOS2VqsdEnDtPI5RZ+YmzcYLU0dxSebvv+yWkTl80Z9DEyAuAKfmSh2O2TZ04xOd
JJveMzbLJJ5xgwGdKrEWjzlONxit4pa9I1K577QOxoLRE3f+0dElK/cj7QkA4vMX1ugE8YJP9Ems
KVN83fJUQr4yguYMVV1yW5sGSe2lP8Jz42DraEaoRnbwTpGJpXSqrW3sRNjIDNcXGfn6/vQ/w71e
1vjaNP3VJ5CQZyzzPXDtXRM6c2pJpHNUYwBnGbDBcXX8Tf3kU5SA8s8P6E37pkIT2WHA58IG0SKb
QggiDiDEcV1ZX0GRZISGO8qNYxRRYXwdA0pYxK4gbJ3Ky8BDkcwCcfYvNkddgQT++rfy4bJm+h8l
ifO8FohG6B4zJBG+htaJvNeE+d51kIqLLQ6QjWfYaiZ3KQV0l5GfW+pN392EnF09fR7KTIhszfeK
JH5fFKaUooz1xyiCM+ysDYpGXGjvOgJuCogwkdMtrZgyxUBHNqCx/lY9XO0J7rKmsxMLbpkuYGUv
/Us7rU5mwjK5eZDFnIJmVPoEpzQMgFg6EgVreJfvMU03URftYbKzIXZCb3tQwvyKsuskXo8320ez
UNRp6FNSFGK6eJBa6hTKtDa3kUSVevFZpYuTofR6iBnOgy9JcQlo1Rnvpu8JAwU+7xJVBEtdVARe
VdCJQ67asoC320loo6HQwjg7Ayt0jxlmK0BN/6FA5Ui5oWsZn4HLnUu5R6ExNRZwPUVquRE9itTN
RcMwphUozyj6czxu2aZx6sUJh42ZdXHhwtqKXbCLY0Lt+aWlzLTc8lHgg84/KPH92cNi7E+vtd/1
lcZLczrKUmLAEfSQuK+/srO30AlHZqpYd634aoVJhi56XeSPc92kHcQwtA5e2VvEQ/6iYTIHW+g/
pqu5fk1k5yy5EBK7nTEguT38vdrbdiwFaSW7QyI1l4iskzeSqZZQ769/Mtjx4iw8E1ol9ywLgtUq
OVGqVOJZ1YR9GLaAqarm9TWJXc285Z0JtPIc2zOxDagLHLZbr8F4f48CZ0njMiC10iJ0ZlDIeHLG
Ie0br8eKjPfrIy1q8T3PwiWTK8hDREYPSuD4BLVwb8vRKTG8/u9v1iHdgBDLlXCP9ruvhzoNJQqZ
Ie2as/Systj8s+KUuQ7Kr1GbMw0e7IO5kKGL9WugSYxz68TwH0GmtECGhtXFTmUkvg+NMKUsBjr2
iF6IKfh/pZtG0VCq9kHDrd5ty8Z2DGHdI4z/nsjGe7kP67FnyMqqzvPNjEIdeC2FGpAcF/mJKVpY
YKr1WgJOCcxjTAHhK3EHh2b7Pb6RJzquF/8CO3XlE6MXEoMnJXPwQcHe34vGNOSqe7m+Rg7TJXr9
0tMFmyF6rpvJHeehCqdHzfo7F5btjiUalmNwTQ40SVRZDxLvreHYoZqzojH97tKcdbNdLPXoLOP5
L51pcVNF2wKo0f3VMJL5OZOhCF7sEJU1XfIBy2AqBmJGSNZcWO1AWE482HXlm96gRqLuP1Vr3iw9
Yv4wI0CAFB/s2+Q4fxSSIJ1pCvM8KioB6wVKegefY3uy7AiyYMLY05nv0Q3zvptdRF97KHARkhe+
mgRid3QQiroG0u6ewmah9JiHSfFlOpetV9y8cZmu9322joyH5BoZTp6+99vCbklQBeg3viYVSMV8
YwM8hAfYRSSgvkIuXZUIYmtzuV2AjUYOq7T/ca62wUrES29UOAfM3BYosFSv2I+YGxmdhEHGmWqs
xQ5l4kFXjgrPDJaIvfi7XZLlqvMIF0wmumEGt6im6ebJOisnjja8J8SVqDTL70gCgQukCaUkgx2v
3ajI4QIPMUTzElYltfREb3q7gdbHJcnwpwHPkTevuKDlzJ5cj+vMUdPUxoJUicRolYTlsmE9fZBt
lRX+2CRKePinpiEiRtsL86YtbvtfRVSCY+PhIKqvgEOTU7HXe+0a2ybeEj8yfB8lIJCF4RuneVmO
TuiN2vQaZqk/1hVMQYAsrv8SguyFj1RWD1cHjvgcU1xCQ30e9SOdaAllT7p027ICGeeQYHByz73T
g7aFD8tZjdsO7Na53p/lIJaOx9t1grOc7F4NynEiJOpsftp4nQFyr9N6Kwi67x7YXCpNeR2K5Nqw
GUCypoLUacYuRPxPTNKZZm6bU2+dGrIlBdat8kwXB8Nnm4LTyEWta5uuDgPYS7/8pjOuPWISuGlu
6feYbbdFADVoO9Ct+nuY0b3ORdSp4AKSthLtxlrwwaGp8/ADOnsK6/785Ii+k1doJk/Iaephe9HH
YKWfpE+1CAZllLdR+hcEayYUqZ54NazcFSm1NOkPAopciASFySCK9nUf8ebrXwKz335kud70HhI/
rFrBmF/+xhoeEhqZo/UMd0yAqqDj/lrk/1JMXLPc9NKK5DXk+yNNdo1AYTEVLhFtHRrLAyynE+30
FuvHQAdLBaEaadHIXwvM/HE1RuHgrmYugL6CBp8SLi+wAdlp4HJLRygixgR0ZjOYOcMLUrcYN3HE
AcpWHz0j9lZL/8A8AOSlDhVYSFELwJzY+cWiuxoryAVw0UvdDzxzi9Y870FB8LSb4mE5S1te1jrM
xHcoDBuOjySAt+MSyicWNMncIZLt5oIJ6vDH9ZNfwjHx1NURoNgwd7L6ouR/7u0nEwbnR3GsCS9O
OM0p3fFSgp8Rtr+A/xv7Xlc54w/gpcRvEJIhHSRIX6lDDktjabB1ydJaMVgeTT/pMSYrIhn4O+uL
b6+NuuJXnD8YK+PqdILyFrdR1xX21E+rqGjKPYJ+Xj47dHtZWKyLUnLpbtfIN/36O1/xp3zIMpVb
6BdpkWJwPB2z7I0DPRZuY36USqh66yzP5dTisWuqP4K+sg91TuvQL7V4wg6BB66P8BSGABhWoHjA
pO1I5OOaiXnhWw6djGEj4np+ZzxPQup4IvAbbHf3sGk61ks9iEXoy3zb3X7hs6yplXSYqgDs3xrv
anHO2BzHeKMEw+8uCcus/TtGbPgrqUPfmVdTE/8Z6wP+DblKPjvOkquHlDite/JizytgfC3sIUkX
e//R68y0rKk0nAKeI0wA46aUaosBbL6+97QU9svSHoywzu14G4SB03Dawik5+SMXxPVpR+Kbhg55
uYsFsNdnF+Flv4+zzJ8tm2uhcOjdrWtTh1VuhRZCv+24S95Vk8E0OZMs16skxrotnEjtlAlOLfce
765iTDt2ZNR7uyY9DbjdaI6XYuPIoipH+mCJ/GsvtN7+Xx16Qx9KnDY7Bob9VFl1qW0ydr3+XHxe
oFM0zLCEVXftg0u2DbmmQ5nZt+ZJE5tbV/1f4EpvYijxcCmvhz9DIaFTCOgYEmsNlMGcjtpAq/Go
BNuu6/RWRwTyWnzNilVjf/cMIZtNfPSMcJgNZ9GDUv4/5VFk5bgrpGf0AO1OcqBvPRm/ishu+yZb
qk8rOeOxwWjJbNwIUYW45qpitB9YpLwydEFnLjWZwvOAMFNftQxHlf8Ua+/ETV8bXU0MOSyEbcMk
CPra2tyS3vNka2TnPnm9yqi3u8JrY4dzLPGocN433vzQ+lI4dfubZMPoaRh08LuhWl4WmYRb1VP2
7SmBbwk0eTxd140/P7UX+6nKhqB9T8OfZlnslr4/GVYR2ZgMSgJI1EF+z8cbG7DjRVTCTzoCXXwJ
w2r9gDUT7QIEcfzqvJjFy4v20TO+sE3FmdoA8q7pF/ayeGp/LWXSqy2quFW/aXkg6rC1vOgSy6PG
unpeysDrMeSbm/9Gqhzl+xaOYTiD2XjrB3OizFgqTeWtANMaXQrrYsXhT5Tiq6LZ/Y5Pgx66x3Nw
ZfoXjeGcZ0Kl1O0eQUHHtA69fwD1E3dV4bIxJmT3Ad59Y/rmLABb9Rb5JlW1T/g2JrNsW6EQDtDo
ycVOeWWJeZPIbYuNKJ4GCkY5gpUhbHHlOOo0FOUQFy318w9hqop9n0lIM/XX/7xrPBxeauVEmwLa
Xso7TQLH0eeOFmHHKsTrEAL8xQU3bZ/1n8gk/19NXqvab4Onr+jioKrak1fN8q9n/v8OWdqJuJDU
i2SW/s9qXJNuyHmxsfsFKcj8QYQY13fgMJ/37wZYvb7w7ZIm5gpmYBvWl72VKxFsnLta6Ye5qWyV
Gd7yJFiJK0tSYnab28HS7h8uLkehtdCA4pXSJiXF0e9xGEAzGfZWrsbWJmwfATpBDdKQ+L8c4xWp
BqymDqsKPeECOV2d4q1wLKNBdEa+gXiRPlKf3akBDadSDWjGAtCWKeZijSeLBgj4TACLxDy/6nko
FKQ2S3kJGBKvWvhMh3A0TWH8XtnbqKwAPlcScfSMY2O4pGSQwcCfOx2NbCLuoJKujRy9JVIEg7DD
Tc1jnDBcW2C2ZaPUamzxD83ViMZOwLiuVb/T8Zjpb0nyJzCiw9PEF0qh6KxzXZG+w7IQGVdvtfMu
VHnK3Uo9+zB1GiUUuZ//pSu4Pm4LNegvBfgYs0ljT3brdl+ADTCxW7Xvkx0RY0pLH+lHwHdKFMwD
OQjk2ZgrRDfD/BtLniO7MSE1r2tgfIrQFvDNyIqeyJr1NdmOJBlPHLJafLxNAauOVSpUjgGSLDSc
PHD6JSAVBqPAMQ9C9re3WYSfQmayHUXvKOTqMqrH3GJICGbd67QyL4Y+qpA1B4xDV01KJ3+v0ScC
BjZqSAc0mvVXWtq0oClQvRT91e35arT4VWGq4Wt9qKVtsbWmeYL1RA5dkTJ2ppJex3/7x6csrfBW
GNNSxxYCCVH/eBJk+FUQcKDGjtWxkIAt5Uq+M9uVOhlOBa/hAGYss/CjhkR6ky46DYItlW2YJqKG
vq9HlBF5u+0z0X0czbH47YmzjhPSFub4Lq5lz298q90ZEy+vcLzLYyHKLcSF3889z5CDTrJp+ej3
MXZEP+qFs3bAIj7/0KFYGOLyJqRNDdTSHB9dQf+nQBQbXX6jWSoNqjUPkXMDhcHy8SnrIV7Pywmc
xbJ7rXxjptxzo3bYj0c+Yr1BAzM1L9GRFMFjVOfAv2QxUPoihQDUZOWB3TaSbjzwZ0xLOEdqrM7c
2r1bAvdJ02k4eOoxxInedcEMy9PEGAmBXeST0SXrjHBOoSXPqNVgpqwMaVJGzOQRb2A+j9wZNGgg
+W/Mza8Fh59bG8lxCdx6l7To3NCf1hg4gU9kuk37iUbs+s9KqTTjBnJu7z+stjJQqfnDByogKX8z
8MAa4vmatryroXjLXNHm3Kz6u0YBtMGDeVSCImWFy3l0ezn5k5f6k707H8Az9+PqIFYNucquDXhK
oQmjpr+6nmXOfimd9g2nS8dKdvMZiD4yC9XIdsm68QcjoZLtq7nlEWI/59pkXkCULtF0i8pJQXkD
Xu7FbvSRI/yUf9w5dcqQpzxOcd3Pzo0UmJrd0pf1iY3OgOe+zODWa9n8hAAPD4D8cnhDAeoASSIo
adf//V48sz2Kv8QLZYMFX2cV+iQBWAB08YCkA0nHkkHSHkkyJF2zxObjg2Uosb5u0BAzgWXajFpX
1eSakLSa7I5d6+umyxBO/+WibB4Zqbe6qWebMgD+mtfz0MppPANxGypMa+KP/pWKup7KA9gcbvT3
Kq/pChJQqSoSEdygSGg7WmVfB9nZyiFjnTvLi3rrTP+YeN5RHO65PehynAaQTW+WzAzLsc6H4lRT
XH8cc5lezygCa/R1epi0yuPB6/nhUMqm2xYXBw5xXMTwsM35RDFUawaA/HS/CbVOCiEJdhS9Fvmg
OXbSnGU3RfeHpyKM8ZHFR0jPK1FadzqsH7Xhue6SzLZcW96v5c2wkvuGwdHJn7BUx5v9+gDz5JJ5
hoF+B8+U4WqI0qGaBLzNyAo8yBG2OSrjsxjcT6e9l8h7X/yD23NFv+rCoattqPRWGnVbLEy95Vm9
hliQvWorvSGf4myU9k5UNTYHOj/CAajZQBeaUME6FQGEBo9i6PT3c1ZxYzicuj6Zs1kXCiYsNoKd
HHJpLIPaRIC8A+Tl8YQ329PTkU6WZRklGJxkaRM4xggI4E9Rh3CEto09LCYfsR3P5tB5cvhGHX0S
G9wjBVlYh7pjMhsumyXCoeYVYiuOO5Cd6rOYCHmAUnH2leE7id9fslsKHnS7snFRz6U3w3Rv8Pru
Cl6zhlGqVKT6UcILRXIGiA5YGoFwYs8suLrds7nYEP9yD5VJlpcW7fRZo/ZvHqfcmUWQRQVSB/C5
FMFcfk52dsBKV59xTT+Ryn23OC23JuhirANpYRPwwXzxLrTc5C6Q8dqjEDvqdi1GUWNmcppwDa70
C9OkJfTy49L0MJ6WuDAjfvji+BNdTnlM6KB7zUsYbz+2XjEAhvaXr5x101HrN+vIdJpGFhpADOqf
7frZp/UYBwpt3KKbTPtkYT/zY3YwsqEa9oZJp9/Z+D7WV3myoPAowGdW2dyASbx6OVzr7zr3bLvP
m4LT4qRc72U2i8uH1QtDcowStbz6iUMh1JJemWfP0vWvAI1Jic/EdNb2t4OmS/dLdkccPHP9bxMB
vYA2Fwifj2cAyM9jZSo1VZskaQtbfNFg2XSG+1uikwy8/q4baDaBybPTmIQBSMYDT+45xqDAqEKI
dBz628+gwN0CpqYRiJ45qYwn1LtLYUn3PRidqOTUjaUSXcXsL6uBx5Q2Q43sjgXx4rnccod3LuEA
Rpr2PATO0w1I9oTn/i49pnzGPt+0rUXI952qBWlPn2ZiuZagGVyU7pVT8NbQyHPtJ+lMhfPcGQTs
lkU01XXAzwFDqdiDeDO6v/pHbm/0wUx221zIjUXaITLwjEHooTq139kl3W3lpsiQE5ZtHVVVe8EK
TLSk3WkqucFNbeucI574kXLLhKxfxV+85XyApeDYTO5i1r04+Js9aB1kTVedTBXF0QMLiM/4xQNb
UVTQmpEhDAbbD3Z0Y/kiSjN4yIabEYIxvfPeY/c0cyhoudwK9I5KnNzpf8pvKbDRShK6rvqBKYi8
wNZZFMn3upIRbDtuGl0fZun4nEisG0MpJ1FcGy6l/y9Lt5hcNsg4PumfcVVQSuuUhoVwPQ1ZIYzH
HjvZzUZlvbRyOXK2mX55nDNFODj+bG5W/SGjVA5CYGoA2uRsxh2ERHkHbUMrP1qjEFhL3ePgga9L
tepwJoJRzlWhdndij4Bp9LoGv9Jh0LQorN/KGg5JiO0Vbad9rYiSFIk6TFyfUxJr08Kdf3H2uxFF
YgvIAJqcnYXh9I6WtQiwx8js9ah2yBR+5qCJTWzA+5d4jVWf0b5UpdRGccoMcgcls0le32+SDyH0
9u3bVu2SN/1MV090ifODn4G1AZYctLlW0UySBWVBBCvirKYOjCIqJbLSjz1J83JT7fbcKPrQFHjN
Z8xoItnaWVQOSU+4LRQx1R+McdOebeZIEL+fErmPQaDZNcCcTTbh6dK+zlJoIPnfZJgna/6hEgKm
07L/yHstilO50Yb/xX72DdWPC0RcGSvQhE1GQSGfrmgAvT3hy5jMe6W+W7TzGQt/rUCQrqVfjAPF
32l052KlnSlyo8eGvMUOooLnniUu2aV4larVbA1s27C3h64gCh2qwVz0bU5L2U/qvPP0s82Kndae
Xje0NR08pDXJRkZZToMucvumZVy+EK5Iz/X4ce5dFlguite3rsFxdKnW00mrSoAFVDWOQUuO4ha+
32/EonQcUpQ6f1/IdJ+SdAYcpTO/z40QYykiyEOgDdyoV+bs9PYI+RlQKQFDGOlGChSmyqkNcAn8
FPi+dwROhBxWgBbM+PP17y1dVw0A1TarSOqYMDmZ4d8iGcj5275r8Y65mKftUNAfqHFPu7qniE5f
p0F2WLEQRmIa1pJ54aYVpjcAHnfeSNlT9MI2vxJB/1fY3bekW3j+SWIpQngXIwDZlR2HngjguryK
V50I4EZ9YzxMojBCH7VwxAEChG9sxoiRxJ1dlpHcOJ4+QpAEWy9e4E7SI50cftmKNWQ6KNoaOx4x
f3Q9FvZ5KF6Z/Kkef8gMP2BF7I3oDzdx7JhcIaBIcEzA0yDFMwpp7n8o33fG4KxgLW3gJjeNmiOM
0rkZlPYvO+/Ay4Ov+UXaprrEwfUvIj8RS/kahoJRmbe2W8B/cy2WA8Y50VUB3Vd/IXxYYy3sB4Ti
dkgZEU0JGj+cI5bqUP6URBtK4sACzXjPVGgXi//rGTwPckvUjiDMIDAbuIkJ0bBj2EaMSUkt6R6q
SBtmCAy6iJfHsD/Ve4+KL4QdSnp2NFIcdocWqAkXuLrCt1744Zdc0aduOlpMLSFGF8SdWGapUcgW
XJwAf7YCrSgXdkQdYqvoKN9wEdmjLf6hveNWCyyfMs5SvoxgCroc0VekRcHUmjkZ7hCBwN3qsX3p
OuIeog7Y4iqGu/VRHTyrurlWCbDjnocrh4YVNp1dQk7pE/b4YmmFpIVJqz+TXqaD/MTqM2aal7Wa
nmnihJGs0YqGQnF9dnYt5yaiK8mjMgC9fHtsuljOq23G3l3ATANajdXlDYCSjmWBvERa3CbJCtgQ
ITdifjYbQYvo4eyOg4xdcfq8SHSQuXDGkIbBo2bubipOLwu/sbt3PbspvBeXYU+pkHJxUwqVFH8E
bmEJZ/4z8sLAxQzYlp00WweYxGF+G8pup2RUhlPgjg3PzJiBmem4kMOtYClv1I2VZ41vTMfLP+Qb
KPnL22ofWBIHEOidLylLef7EcvFPjkH7BBCOmZebObpY4hl04WZudtHYyFOzy/jQiXn6Nk0ksdrE
Tg3pODFH4Cx6HvajsbKl/Fn8rl+1x8KjQTSed+sbGuT/OxoUI6J+bmhc1BnOAnRvnjgEv60LYAID
xJpEo0rzWqH9soGqv79u2yfQtgj+Eveu24H11sd3SjUdJtGJKm3gygeY6QCfPAqULvIk4o0NaVfP
TxCN7pHjGpybQG65zJn3oTburBF1IF9iheJeZm/oRlJ/mEO1NOXOyHclZ9s7lmOv3qQLMk/LeRcF
KK+UwvcFt+TkVdWwLrOXexdUVOjhTNsbuO3x9v9ZPzFDmGnQFxtP09O5nXhselsdWXH0EFaLQJB/
EkzUrDFyG/RkAQaumu4wSTUIDYx2aVWqVpkfv60KDw0CryaOfk/0nE3ast89k+OPY0Uo6ZIaMM+I
PfDrPwiCRoAO5kt0+qdS+VS0O8YO0BK18oBR/AycA4eMZ0pc40oppTyy1sumHRyJrycqZRcyOl3e
1Hu4JXJG/Io7RTmi+IjMM20m4/SkfSzuV4KXCM5kPPInH66cN0iSVvriW5AgOyWAINmjDUERrT5z
VOB9Zmi9j8w5Vyg3J2nSmRNv5TA2sbm8ou1gEZB8LtQEJQY95a0FmmIR1jI29RcaRhdl9BJQigJh
LsrycMKMK9hqp4GzOTC5EqbXDU97wj+myylsGBrZOaNrCtVu+wd4Jgf0ObMBLBv+B43pMK0WPCvp
Orw/IWcIK2lqZVerm9Tvs13HbMm4PN3qCj7KYhtXE/1R1kIRYSg/E3Xioi53QQSwrFnw0K805auJ
l5A4yArhyQFtU9NYkdNys0AjBVR/VsZqpe0sYI+yQ+jnPXoTt1Ln574B6A2VUsHAm74XcFMlVg6D
dRr7GhY7iavxuGF+LCerHsbPgVbO1BSB/wjrk3WhWXcRXsD0nSAHm45TGvYqvAwy2ONzl5/ayJj8
O6B0C2PN8pIYR0/VJuCvcN9/cHSqFkvzBLouV8aLgatrLLGV1zFStcEv6I4hAnngLN/8tdHPnCJ8
H9l3JtD8CAl+77BnAbUddvrsGRwY82bWEq+T1MFDdToS6LkkqGT4maCNl2NiOG5/HcTsiPH1dMer
dI4k5ES5IHVlUQ1PxL+bpJKlQifI4UhNUAR5YT9vmQgjnk20rPwCjEPmqFToP0WGAsxLg4F3P3iO
GleJ/qsaiU0Exx5YqB5so8wpJoKWVgsssA/ejmjulzseSB62M2BPg52Kh1mmooGvnQyGOem7UEqW
4tskW164p8DbVJs5vilQJqZxE4/0rX7QkVFagx9UUFnCb02F+ToCaDWhvAZOQ1eOdKdMNgmB6iLC
++VZWfXyeYFOr7Llt83hzrpsD255x917QSbCaY60oCBy4DVndjfowvEYUSVx3AAteNWkqDNKXRFk
XS/qrdRW+E7ryRhk67JU8JoHpK/kqPTjPG9P0cStVBN1f+/x23uxQQL0oi1PkWeJzMAqd1fHlDxc
7MMeLkBXP4BwfznSHi9DAfpd+QfG063nrRUY36IB2eXpPTJ+BhPClHEU+TWSjCsTSLF2zNX1IGBG
ymBXvitJeKoU8FxP+00uJrkZUvkYDsmliZfbZGnm5JKTnRZb3JJ/33Pe1Bck+gAuld7VutA/7j0Z
napj4X60DnkyD1DTSQpE99UX7LUAhZksV7xYrEV4vfflWiInGNP8vXcJ5Yhg9WgoiMShpWUuHnEX
7xKkGExyTx5jBX67gVWelTvGdEyq46UlLXtv169T5SQJd2OW5Uz2kH0KRoqqWdsAlTKQafxqPDar
KA19tW258L96QFkdqAM5DaxCQKtGowCki38L1mPGK9bpIuuwJtJVpuoDBlTS2/TrahFn3qgr/tAb
y8GvJmFaHXadeczcdNeB1JoT4zvt/jEXwYGoqAsDhOlxmtp4GoEel5erdgEU6KV4FhgBWkvoMMYZ
/J27v2HSRvZM+xY5SmWq9tjFsi8q2R6JPreRL4X4QVNial5MH4F+LEswNolCS7W62IB5Nuuj/4h3
h0HT6wOcn+BkqUVs19RO8DZ94MpQkMi/6kaCK/A08LukEYOsYCEC/RZoLIvMBfRIW7tZ7HdutwJM
xUygsbAggSxIBnRDznWonN0QC91NVBbvpW43HIa/RhRdkatZS8+WLkoUg63/pdN6NFh9oapRfOAb
24pvot+1AtLZUf2/H1olO+KxP3wcJKpJlMsmdbGpRrt3DEC3c88pbUoeDTnoWoCbJ6PM03/is8XG
hoKLIpurSo9Bvk+YuqqCOoXHuknaNvOnU0tJ/E4l74UUEOQ5LZ67w21jwWf3De+ovzMnkd82vlCI
Mz9Fyr2ggoDZmU2UJ6IYhMeSFi2icb7XBQmr21mNv4u8F4vq91/J89DDHUKeLWiUkUtlxHiDVCjW
qDiSwFuTsEG1f4G6Ih7TjeiGZKyXgeS2BT7tbvTSjpToqfydjyTehuqy41gA7tHOJrlb9CGVOPKa
Z42hnEY5DdnclI6NAI8xQz8ZsZhToz2nqPZ5gvBQJcN9gOAl0l9rnYcWm6luuexFY4BJ0ea7jBSb
O3pdVDMrfW8uTyV/QFYjMqV2urgJJkJta6q89XAeyqOAqTIJo3YWikchtofnBU6REiICDs8qZEsA
tgZLIWiwrLFo/auYFk0w/siJVdq+tRvabHmUPI7aGi03Q7Z9uFKYwMsk2BlWmSvsh4RLkcmsuc/y
FvqdwmRP6YUK+4jLOH0TPsR2GThSPpSEbba8AMupO5YmYzyVfhIm6hkN8JVl0eGIEimhtd+d8dEq
XPyURr6WROkh0qVkAVdQ/HhysjIPxiqDhdWh+tjIylY41VrIM4ebeUDu6uzeFsdE4HbGtOwiQk/x
wSJQ7PRl2Xz33zFsnFh/mVqNP5LFzuNCu5KRHK3o5NZdxGmeCIQImrAmyxosEaM1x1Ge9WjOgBAH
HACbs4xvbVS0t12itVDxFa3O5bY0DY7aioOHXlOust8pBFEkUw0uwNSQTBPKjITfCLZqhHrmau+U
grDm5SteYLGuuQJd6Q4r65Ui+4nGnnxJ9F0O8TNIGW2PcSkUdnjF+0SsvjeOjo9/QXGm+AQH3YTj
tyyWXiwwuY4DetCU+LWT/4kX/OPjIeMRFz1gz8/YLFhind08LATVByMZDEiRjiCz7h0sOJpiC20F
DhZYxIB02mzKvlVpKszqa0b/k4lacltKnU3bzwfSVY1jVdfcuIsBGpyYNIYqXzbid++1lB5sVNXE
gUitgLyh+KTa6G7H81zuQ59KVpzB0bZv+aL5m9QLcdfd/5fFyFWxYuq+K+KqC7O9gEw3T2vvAuIa
lExYc/mWC7NuixvYBU6+G5eU5BLZv8U7sG6yJ0oK99dFbednZdeLuZ0sPDSvJo/lUYuHhIsab1K+
3j5j1VsVhwEAGqoG+zG/HpHaMPfRzLLuhaCMjASHb9iFU8xQxxePLbGCiMD+f2+yYmhKouuIAdQW
zfXWoSd9U7I6rHv2dZhZ8ERSo9Gh6P/4V6xME8SMQ/YHZCmbge40YGs0Nw46Tz9GLiJpRCfgxG29
2dRdA0JDUiVPWKYFnRCqbbAWQNijl92ocyZUmX/yH6OS9SFRqIiNr/YYUTbdIjhqkzsIEypvzYuL
77EZ/EIKM8csot5Pl7Di54S0MtOlmwFUaepMT/XINfi8nxz6If2gV8tF9xJwHsJEmNptBGqbu6xN
ttPuUfyb5C0tWjtqlnLV207QpfHI37Rru49y27KYLZHvp1KteFN0D2RT5JzFVyka5jcDCqU30+dr
CYXSFS+KtRMAAA8kYXHa92Pimd1MqFheDL7nDqXFyo5IIuzFWhXypbCR6I+qceRMr+6ZV2KaGtL3
4PzITRA1hrpU3zSWmjS7++aSFHGwKgDH0a8YV8ldtHtHSjkB0cc3G7WsLwl0ZGDqgxVfDSe5xQ0y
lEUVmYyMQqwQdnXfUo+sJQjzxz4yMBLgCiVCiLARfvV+SQwc8eZCBftSWDMhOQWEdEfnwBbk09mX
aB5p2gMoDxx9m/9J8p0n6Dz8IU2oYKCJJTRAZAovvz0sF+MDyxKyXBJaUMBtLUr9A5Y7+aNk6DVU
lEBrfJC+Otd+tCux2RCCTdOUrBvgTX6wxhtH8/mYxCVRRHCRzn6Gmbbd36b5N1wfblCeHaopudHG
Y+I8IkmQTjWKU/jMbwbCHhHVrPP747uFzUSbBfLppORraT9TMFwkihqMROBLoxa3IwRpUhAa0e1q
RambDTZvEnigBsOFbFng3dkMG4zGnjetPuLfIH6jbVS9vuZOSd7AKU7B+WHH07qWiVfl88X2RnG+
io/xDeWdQKngAPZbgExs/wkE2/zhPEshkd3gUkyoknrLqUHKrhecssokFEQyJhZ0ZMqLWJD56kAg
GxBYGsR/LtWWbmBuUf4/5nYrvYVLnor0NSqyfjDe5Zfr4tXr0LYaCsqM4xzP9k7e3cu+4YgzF/w6
OlAQcAxfGIzbl2ZHOO+zdCcCgit/xJG9D6XacrdE9AgGacPtsOedK4/ikbKINbpaN2Y5dtyRDEwV
UmZrIBc4RUlo4y+hHNWOQDQ8fPKA4dvSLNpSpVd4r1P85gPMq/C14f6ti4ifaIWhgtV16ifnPIbE
r2I+NFhSN7V9MxGb2u3vzoFxHUljG/38bhsiz4VnjUAe4ezd5JP7pHWJw+XKKulf1QpXJovFOvgL
Ps9VHDjBGxwn9SLAc/qDnCdyHnA34n69wT9FFWb5XsNiheD+1CWZOESNXLRKW2FbWns8uXNU0YqU
TJVZ1DyuDfUN5LMHOPrpyXqR1MdheBvSiCoTGCjvEqlBrvHkyeid4Izezo1gGwOsKwAKAfHdLWT6
cdkygbZwcTUGCw/YWLStelReGQuHbWMmqWmhnm3ujh0lcEnfwYSmcht2QQVJk5ClcQSe/aHdcDLJ
amTG56jPKuvHP505yS92U1IkR71rf98abNBK249rhRHv/lo+ZdeovYa0dYzfBwUix32Vn+UPp7wt
Spk1f4ykrKIbv4okGnPEdIXibeVkXzj4b+Md4uuydEKJOW+BvopYc0ybPeBptxCwKzzKmGKsqDdN
WTQfaiPmbW/h/nplhupBf8BO2DhjM7QC2c4ZfL4LVVCnjoOk6m+yOaJodIECYi3o+hlndhssc9Nr
EyXyfzXXoZt0GAQ3DFBauGY91ZzV9+eZnYwvjUpW3vGYpG69CiboYpvjUPTC12M+RRR6vKpICmvV
qzp9WSLhipNATsql9YmCwoIB/nc2kw2skBNkVV4FNTNnalQngx6B8PWJpn2nrOVUD6Y8aQXI2pEj
zMVEYCXzpHmIDvEDFlYJVcUCntWgqHmimxGiRWawjKRUl2iAXRoWp5/Saka3zWV6Kbvu6W6xnYXu
MIXvYK6hgAUTMUqF98JOe8CG9vQxZjlP1NaZ6wFA7b98CA46xf4iuYBpVfL3VS7AG1KXPPY9/BSg
/Nk9cedHBLMWazzEE/+RN1qZa0HKoZ/4JN1AAhuIzzYt7wP5uzH8w+K0HGpbtsZNzKoPQYSKhW2X
5/SgwZSyC4wynSitzlJYtd8cQn/pJzsGBY4/OX7JXYsoj1M/zcI2ovikh7WOz0ILIVI8c3anhv1k
ykQrIJyGnSOuE6y6K/LrmWCbqV+5Au2oSZhz+DAWB9ogq59icj2ON+Oo/KrsiOj+PhPM9EwQOT3s
YIqvsXl8PPIeRV6EkhSPdJ2XNYNqA9FFM5rvdSNRiqyaQGZm0YxJBxV7wmnVxOr6jD4M+RA9lDuk
qRU6jTX1BHfUKiG8Mi3NoWo/bHGG2TdKgf5atJbvM+p5klpY/ktifKwWjLE8WYWcay9mxipECeRl
whVnlgRIslS6FtktdN5M3S+NgOxE3ydN/R3+nyUYe0Z0HfNxfTj3d86EfkniQ3KCZW8cX3shDo11
LUL9Q/9iVitBehrIgNpqldDYj56Ul3lKKFcCNJ1OfxffNLXpSb4vRMnJmt1iX1C7eMvFKJlux41P
X5t86W5p/15zGtlHIdQle66s+nvU8jOmnSvLwpGMDDD0ZW8yUiwKXrxjlAgPC2rEGLhZIKQet6V7
2PxgdTiEML5IrH0glYUhJKDaAwkZ6XKcmoPQ9t0CAykOfCTAtoUNIqg7cHxFUD3K9mk5GK6BF1+p
mIiAEmDRxlNwfe83ujf5MVl3WhF8hP66xoizp/BU5g3n7/YDGzzxoDNDfnkW34pwZCYsbc4jgr2z
SaqxgHJ/7h2mYYh5iSwWbNrO8mkRTrNat6VTNTcIpdb9PQqol57tX4Zcb0ji+Uu4A188InWwxv1L
/Nr3gqII9Cn4ZMrMINOES9j8u0VKkGp9vEwo6cSdDvsZKy8pG+oNsunej6ejc4sRxYVdUk+wDVW0
ugJr+B0F/bxowKx/4lLmzc8mafngAIK2gD4cDPYNMzmXbmSwEtD8/wU/He07zRtdoeEaE4NqIgkJ
9EDqIW5VxGMPhcrpXYhmlVRuZp1XXvqsJwpIXSXdTtdm22fGKyyhzKpCOo/J6praP56YsDwN038p
JZDhwmwVIjmkckPrXHNRXRSlB1Q3c+ukTz5NoRj+JHWNqD8UjNDJW7IAGCcI7tyApDB2fWtkngiw
avT1mDM6Dx2sNTwjfbQtQd17E+I+QzVHMe16fCZmfwPGrS57P9WVzhXfmqcvZWDqKogfPg9DR6k2
15gJclqPPo3ibW4Um58kd3Gweeb2bcyIUWRzpE5CQ9NHo684Rhmf2MB2A1QfWemeZ7gHZq/I/xbE
jhKLOHPW93i0638n3ooBwbyx8G+2TBnkvYLyuHmXjGZswX0rBVn49GmlTp9H9lJFO0BHJZTyYejQ
UWbBqVUWBU+sb/FI3PPYSXjdlEL9hKuLsROozgve/jVKaMMVaGS+5nzRLSYBIdzDS8s3WxDuq5Em
5Ofs5mB7iHIBNXRyNWE8rEsSwB9p/GgSZ0B6oZxFWRUoci8aG2l0P99pA9T18r9AyU0RzJ/hlckb
94rZM2VSvis7k8Nbcqv3oCC1Q84zx/b5KGwuBqrs4zizgBymui8hHo+P5TN2erVgFp1x//u4DIPA
Eqv6EcgQzolwR4htbC96HfnJf0FFpJrVaOBkYY6nQcW/wuVlE1ljuRviZQcMK7nUZ8wl8mKh+2Zj
V9BPuh1b3UtijsGQswThUyl2jsvHk18n9FR4JF3UgxauBFh+aKl17wz1mcpcp5g9BosPJzkEBB8B
7YBLWu/HXPchGLNrlemHIQZiXlF84g+9RgnSiiTA9Y8l3JybDiXtUVrvZieug1afpYsyoljFxOIT
TpVDkaCz+RojIdyQjI3o2G5ZrovT4BO2hExUU4ji5/BhpA/dp+TrvAwxTBDTYOVGUBLGEWlNBU8s
5ks4iNXxG+a5g2ZzdsSkukSV23HCdul/T4SGkN631VsU16HaRX+hQohrkdvyNgSIWsVsdioOULi3
qqW+nyp2qyPXO/7PNwd3IKI3l8ZtcAeedM03WpuXKWrVDRA3lbdNqVfSxbLgf41qY9c5UNhTkhDA
qRhIythfwLOhrrV+w8/h8BsJsCF8MSAXgMycTwOg3+SoxgApFHUpDaEWSakUjj43xy0QaRRkJRIB
XlorALZWaLlK7ALyj3V/Z7azmsvlhTeygMY3FuwF58XZUzhMOc6M4uJH4rpqrmKcTzc8QTVpv934
uoszLO7pMNX5gCnI8XyYbgu7Y/nNJcND+YOWBoPKnGPjRYRVPsVQh8xMFBgVg8oR7BF4kswS26az
J7+X2IKtRWV34Q2AtNl+CVKPL6/+2zZ9a+6GfVL+x9vap0VmljhO3YdyD3NMwtwA1m//O9bwJZKK
k69AO5ToT3oLdgUL087IE2ZZwzJEJvy1NdRfIT+0SdObEUmGx3M6Jk5FmcDT+z2rNbDi79U4TM0L
L4lF5qJyIKcaPi7TyC+RO87OPBBosMzEGDj/Zb6FZdwWyFq7wwxrIyy1j5ydePYJM+4x72OAKUin
l9PUS4Vs3ODfZntvX/nPiPgdxFNhJc/5zgF6L4JZyuUNjNlW9z+QPLVHYROHVqqWGseG8DCaPgqI
+AZlysHL+Il/0uVAHwCVah4Z4vHMCha5lgQt7NRr6gruI8ZQAsMwAk8T03GP850ltbuCtCo8WGsi
u9wpNzPlj4RgBnB1ekEc/BA6Vv7k6d723upy/JgYNL+kVRNw87HMkNnnOR2w63yjdPCgJ/Rrf4pz
8aJV0ledOSxbSX0Hg1B6iUkUBiRA83mM42uiMZAmMh0x8aSmMwzXenVOTDmBe/v4MJVZ4colfcie
3ihkAxTTf28VTubGGhqKTGObwzkC2Q/8+B0RQ4bBH6s3GeOpcFkxf9EczF41siOR2dhrYFDYuk0f
QHW3oBggjMZF84MYbp05mHGgYZ0TYArBpjr8nZ/q6RQKgyPWAM+mDX1TFw5nJWPA0+Jx5ZTuUH1M
NnFwpKWoHF7xl/59pZR/HMBUKjBvLbyEjDdmpj+u6VVzLOZTQRZ/LeOsdZcJOz8f3wM6vGmq/dG/
4FQ4zgoVVZwwyqZ4/DYqa1yQ+0GV+4+T1wt2SvaWWvY1hXDOichq5vDwiGf++FdM5h5Dq+/aXUTE
/n14C8EE2MMv5ZUSxWLXZz6zwZC9sfQxyDHXFrFchzwXI/j823eQt06UTFq4Muy63gJFenQrSO6T
u6jZf7SA8eb5UBtTilLsO0v9Wtxk81Z6EY861xsm/5JJm1y4xIK0Taf6D5LhkeRpDa5sojtDdZr7
2E5fVC21ZAr5repX0pS42PjBEraiiRD8y/VzPVfHnXUDv41CPhpRS/7YWAcKZjm/RmIinR8z30/e
jqcHJR5yS3R/Je2/mHDoRa9w3XBEfu+K6d+cQdtYfphaRXZfG3eLceuXHLfrD+digeP9BjUXa6rP
NkcjDAJlAo+kdKArLAceGIGL17gzNZA8bHJjNPXCR7HqW8sfULewmTsqPgbBwHTPpxVbxGXVuAqe
KFm/LePk0v71+v6iwwYdeAqOG66WbVNs2oHk/OmS1gYImpq/bt/CKjS+1Pk7CBYL1RhNC7c1OShv
oLHRwmVUoO/JgXtHv88n8ujr3NgfWbeq4HDx1j1LF/j0PeotG7cLeHk7VhcnjoOdE3Xx07ILnq4m
PinUxXarkiX0fBZ/JzztDcS6lr9vWiEU08BfjgX69QUS9eHpJ8v59LlMVi69DHlw7uYE0BceTG/A
cXlu1VpwKlmwSFYkp6ysrFXwz3Sj9y9M1xRtZWQ//y6lbbXrAUnWzvxnjaLII2jUjIp5Yh70GW4Y
pZorXuD/t51lGVd4V4B4XKdpH5cCEIVKPoeLzV200/9KmDyePNxuMGZZ2AeVCv66qp5AyO/wBOj5
cOC3yyKXvv0yAAXvTsKvmRCzSKcXIbN9lKamoY82zT3GI2axuKK2SLq/DShtu3mc2INWgKGtatCm
agxK2mnw308v12shocuiML3XSXObYsPZvH9qwvE7+j+QdIBsOvMbFYy9UD9jmlJiKoltnXtxplSs
4OOvoufgCdYcGkTsta5biz+e7Wp5gUqtPX9I/voq7Es4pz5RYla0NY/BUxnfYnsP9VWjsAf0BhPm
r3aYBQ1OYjWkOBZnLMA0ufunuz19OiTwt2VpChpfn9+QVjCXoEXJA7KVwlli04srVMOPnKNJNGkV
kgGXl2mJj/zciGf4+U0zMDMOfFeOqptS0dUMPQhgJzQGkGzfVJhQw53cf4aeJet46SrhCXzxQ8GZ
JzSKxJ+Dhu6c251Xf68nPlr6ibdPTcJbUSpxLlphOkZM9aHtAshJIkdJHl1vkGBwrzSGELmJd+/M
a6ZqFPymvx8vT0U+l0Gxde24sKnJ56PxKOVamtIbVzFO2lgyt0YqkBMA967WcSOo/XTUlVvy88hW
xlL39e7A3/9YLOlxN3y3uvoUUB5UYEOAxZHjCiGSRPeLFEKHr9AL+olXgYf2WwFS26gOa7XYQ/Wx
91/U0J8W71cw7R2G7SkOUO0JQisFR6Ms06XBLliHhe1mCqe9PlCJU0WISAtJPkVyb2t2Hc1Zid6E
OZ7jUppkSoXVk1sfzmJ9q18j8uf4eHFMoDjV3C6UjKwz+l1oJFh2JaR3hHe8Zbx8XUqN6fM+e2tl
o4e4L9wS8iE7xM+ifiykQpfF00U5aClvjE5/2dGyA/mCNAszOZGmtH76RltTUF2IG7I4HCEWhuvQ
p+9BVJ/RNNy9aY6ZNCw7hz104U4lZJq4KFuPPZ7NbfdEmcCDBiu7cXt2h21Zhgbe3djwT+dbHSu+
lVlZDOq2gqMv6HwHkqt6hlXv7++RPDtJi9EKIvqPh1KwT5O8BV/JV8mCRzDPKYr584vfLloF2HTO
CQ7fZkhU4RN0Dst13W4SFrOaR4U8CGDfb4GOnxYcFInv8giKLe3HUXJIUoP9HXDNr6ekkM2K+ia1
FAe+oVzOYl+Nr3cRRDiSiFbLtBPgh9UdokT6COH0Pk2++S3zz3MUBMQHweZ9kepEgidO5txA9m0c
EDTD9mKbNEKApd5+FkeBNFLYe0tc5tOWcznmoGwbKAQHOoX8neZcbOkW8rMDXLtmDpJ2a3yanKeU
kZOjO5WF4sR65K+dZ+rbMMbXBQzIfETKqYaSITMThh0V7y7Gg3UBuTstVhVg2WvOJeVwfryw6APF
V/Ss+jTbFPD+Nd2RBHDy1k8NlJgFkMjREHT2uXOGZozWa3JU/P8KQIzBUyUBxmKWmkal5NR1+FRY
fHKNqlIUff4231YLYgVII2gZ0f75L5LDePzc88VndDxH1wtAIxiVSXUVqc0y+JhodxMsPE4dzrLb
n3lUvE5RHtt5ewRQezQToVhhgKUY8ym4euRJSW0gA4S1SGT8H4jfk7voQemAvPkXW0yphyI7VuT6
i+IZ9NE8bqo+9TMHyAEkfPB98l6G/k2zR5SEQOJ8ugEcHOQdnugMbHFfu8ns/8xV4+YQSO0qZNTD
hFYA36fgZcrPGuDMdcDc4ReLeuwEaOZfh20CerCT8ZiUA3nLNvMLk/twbr3DW4zvIOoA8G+lZ2YE
fk3hjalgI23RMCXNAxKEggsDcYykIEhcLNEVMZ49/dfAPpoEhzeJI8GjL3IDGK0qH4BDI68aXk+y
NSpFhsUv5gtvZbCvdp72+znSKaFoLOLA2EJ8GwJs6D4SszCtC0V8semMLQH79/Evf3HE0OhW6B1E
ZsArDqQxTvG2i7+AAeG/rOmZ47qaj8uvLOVqSxqVAPEHtpR1oAVewCvpmzPPIzSFXkWT1oQR1pyG
GrVqA2lV5fJGr+CzhWsFMKeV8X0Dm+nnCLT6xnYoBZLWM8SpTxBFxD4SASE2EminEVFGZccG3YxD
PHBjiw21JakR5gd/cvJ/zoMwkpni8O3oMuakTntXxalFI2Y1G9dGW3j2+NWi8giPoTHcq9rXUGdi
Nhe2ZkiwW+QV+QQlBSFH/Hk63YJvhVjURZvsbckfH6EMJ+sGF4EMXijIQlc/8mc6KuDAgaLQmFza
t0mYl2mTl0LY4bwQwhFfTNzKaZjSzLV8nBf/Dt34DveiWCumrdQ9nBIHn/M9SVtYc6fPykZ4ff/n
mHK8L8/yZUNX46RmJQRf6CnQ0pSnfO7fyqFCuNLXPGp4ViOx5cOB54wATpDqpiEbA8g7Kfgu+zG1
/aevNOq7XLRWOqU2D8aBv9+t6AlVuf+w0ln+y2w5BYUe3CSFLgIglyQW/FZfTPWe+G/jC58U8hYR
5p5IqokK72jBebndFZ7AaQHjGoUzefC+KBGQaGZHBtoJRtHyx1KA++/Yahm4xQDqqSU3Cxz2MNhb
VeF+5t71wtKzkbv1XKvlDYYst+lNHxXlWSrfEbMNk4iMljxyEB3vpfsgCNW8furVqsvruc+C45pz
6lLaW7ASro0tn5FQzDfmI9RHAa/9H9d4b8jiNrZFBGy1++K91NJystKkoxdY3+9mnxNccdq5chwn
1arT95Yok1RpDhBzxg0QJspBhSw43Svs3qRJ0KfByEDz0yYyOXF8A4SKRhOdYTHbishVkOaQNexb
Ie+5ly16KRoycpgPnOZEX029A0OtoB5CtpTLqkOcI6MaYrWuIMlCsjJ/QmLFSOLgPMGGJ+vxPVMk
+FhXbwP4cdIRloJiQMIUC4HzZHzlWwjOQBt6knMH32pIIxYHqxcPvisdg6Poi7oIgHQU6DVWbP2a
a2I9Zv/GWuih9mICOMNAEnRIbT5b/+ZK4bFbFngt0qFz16Xfw6YC0lkFfrVWS4ovMBSYyz3kxbT7
60CBsbodf9IyeDkjpvH9i4UGJqFNRN3fuH7itiD2ou4UUc31DpbBrfzh1ZefNpVqISp2eeFhgNtK
5VaaRpFu9/fPbrwBI9jpy0v3WMvT2TagUgOF6GRj7ib8OGMe6OdJzz2ryZWX1F7z6zIAJi2AhAXV
f6pXBqlP/D8pjv3DH9+V7tdJtJw6GCDe+Ov0vourdImGHy+BkHLPiCp5fOrrks1wrcXNbeGPUmPi
o8BLJ1e49mOXKGIC+NAW+dxPdPrOE6mlxOuk8hXqb3zB9vVRWF7qNfxCQu9zGrsaR7rpfEpr5LLl
zetx2Pj7tcb311hKUl4q9K1+WxhSiqfxEdwBCjY/i2S6e6TgYHhxKuF9BAdn5kmalt4UKo0GgvII
0vq+JbDlQcn4z6o3W+liCgSV5hJG7RSxD4VwJ0wHd8AkN5/5L+Eh5BBtpUHiFqY9EC/YvUCGTCwi
fhYIPie4eXWFP0BtyZuB2/2umN94Sx1efXp5nDa/AN7MUzByZCUmT1Esw2Y5c1ZFryfh91Ly3Fv9
lNO4r/iW2xFFWiv4gZfaLA1pWO62P3rgIUmBsqMMOC178fgsgGMe2u1ZtUDkD2xFPy4LdIoqvnlv
u6iekCsddvAjxGAudjoO9hTzvrnSNIDE+OOVWz1kvr6TCTRSw/u2RZVu+mzdDu1sYJkAXv3TUpfT
Z+1nEJclXV2PhH5BKRNdV26QEtEHTZ0xR+pcPFTIs8qWOa/iDThHHu1ltWES2PzddTqyNEVVnzCb
I87mYSYxYSI2hPW/+QDwK1Aadbu72r1LhF1g6kT5z348VLvAXFmJZ7vYWnxEE6R8BmPmHI+/Wzgv
iBm8sQlhlGMB5CdtnGF+K+aJaQhvLwmiwi0Gg/Y4xPXMVVpGoRPBN7v86VySh7iNw+CM7/WnFEf9
Y3CGn3dNCm9YwV0ozuBkfLL1pymS/8NmA6CzSb6E1vwm0V15C0Cgj3SjE7UEbuFT79dX6kkNXAzg
QSU3GH5QTqHynr02uzfAM2tkcg2HQUXSGADtBGBNLV1pRR9XdtHVc8v+qBuvdCAnQL/Ek2PtkM1Y
ipDPh6aN8eDMbXI98RAQMQjbjutd972BTYFdSa4J1wNB5Eevn7DHLd58ySF31VoT8z8zzhpwitPa
uWeSXNB0BxR+3Z9gHUnkHyLmCrDmq4UPfiY7EbUAwlAigbKv6h6LR7DpphVwEqU/J0obaBwVJ4f9
uu9o1utycrHebEZUflg47AqaoHRPIx7gfFPckn5s6deM+c+rgCc5QcHwrj5FfU6W6azjvvPP/VV7
Pn2CvbS5xYM8+jFST2+mChzFdJG4XLJNG1E/dHReDdQalBT6tjVxUdUV5/P4VeWR+TS6jsh69peQ
ZI5tUTlVLzUPhCvNnyEBu/KItq6ZVWGtKJsrjBqBPPM43yNZ6spJGc0kUL4yXXcvTeSHaB6+zkf3
ICKoOeR6p3QdSOuV5c9AVAUkm+j+G/ZJXl5u4NzWCVZVAvEeoyBeq6rBgquMmAAdpJwB0DJiFguj
MZljFADnV+W5x7vJTb6sZNkb4IgBCGl+0pQLlg6snsZ8QF2iCWgQr9spCHXO/u+11Sp0g9Tar0Gs
9Hk+1jMoZFRnddtuqpmxEh86++fc/Ckkv2B2mqwqpZJ+mW6RA8fsIZFgo3C6ju9Sgjrso2T8Yb/y
nSVxCQwjV9NiqL+kZSdFh3KhqnOqqou6ZBrrV+feKf1dtIW5vWrwGIH6DNluQG1CS+Vu9aSv3p+e
PygNGR9lTmmZXODPWzuP2mWTmWS83Tif7dFTXP8hxLruV9XHJjrvFDNl6cixVblms7jxQp1ISD0/
vqeM25iLU3IWKZoJmWXNTOOHBP7YeUmNQiHW2hbOgFFGxPbz6/tCyWE0TV7f8rFxvX51gyCOn8nA
Whlk8rzZTFnC4Ktj5NgVjlHRNmn4Tcl9jAjcXNIdIo+J0E0MuB8n2yn4tVbxGcw0RFDMG1bgtxr4
+zcWvuEl7yjs6u7e2XngMOJ1BDV5PB0N95Xdoyql/MdRRvicMM2eavR+CF9qaRvqoc2guXcLpCyg
obkI2L91DEPo6lcI0unxvg4uQvCfHGzuqEEfh+diNizTRUpZRGlGcJzxwXd79mitF6wXS5ilnX3y
Kx7E92c3q6TpXCT31CFPJZberNweVWoJNE19lIo7i5HevW/8nppZf6bKiW3CSijXJ3mqQY4BJCML
Mnw3zkaOd2kj+Jdkd/fyGhQp8y8P6t/v5tGJ5hecbF1mmLxJXP8R+aI5e3qWIHygD/1dlUeGHSeS
FZw+dC4J1j2SQwMsn6/SHfZZdgqAIGcLFCaRxFDuiMU0HxR/4YBlg7okrxS4R+sgMMEgjrCOYKKw
r9Lixt6LhGZfVxIg2g2Q11CYVIqXq35Eb3Arvexq4nqNHILwtCEJ0nLh1cbZa/u6lj+yFuE4sGYA
Jt1ZHA1MSweR3XMl6ajYAyQOM1cJXyUsInLPQ2ZwctWSoeriTDBnOuecb7ArSX2Xv3CS8QjGH2om
9NJBwnGjEYUeNByUBkqd/pP0XEu9L1kOriZaoYuV6NvL36HRHyYZvq0lGtzrZ7vH1LdbQD8JgCMM
Fk1l6xvfrXDyu03Hy0fm/egdPt6to6SQHHt00q9HpfeiAtFUTYnWnbm6SeP0mZeyEC0qoq0IcTfV
6SKLFpUJ+sOkLtVYamGyHFvEgmINjIUkR4XGd70TWbGDCz3/OlSthklYZIiOo/lS1DMzNSaart8i
yFyBSD6TeBeJ42c/mP57winlYIO/QyFkmFhkFxwGr8J3OrJGJL+FVuwukl0FLObqBummUZzkrv4t
3xU7tiTSwUxB8EnS6KSveKXsUPwgYJd+CVWaJhET1kOha1xOY0FLWR3GQJ8bCepB3nH8TtoO8g4a
cV8AN2BSgv4bhAXUcIGQZbcCJFFKno7L6aLwuGwjPzbVfhZH2XH4y/4odtzT44vIQhrAgwhwaNVM
cLBhDad05p9umtjySgQYLULTxcy9tdKqvrW7gWHE5iLbjeWs4yZyBlfT0d5ulwX0sAcyE8k+Wa2c
ibjLzI3Si9++FbpktAWMJ9+QUHA490aeFZEvBLn/JyO8dWlu6NYw3eQDwSqxyHKFVUrkEucqqto/
8FCqWLwr30RDM7O1N8svztwuBbBgiw3f9oOnWkaAxL7w6l6vvj0Nxn7cRM//9aSveR17/9gzGLJm
uHObls3gGa/lxp6giBe7xVnG8gqq9i03GAzT37sQ3ogchM5F+XTdQjG4H6PC8iO/NT8D24QeTxwh
AqlQASImmA9cmZIZhjBxLXsSuaZEUVVtCVfmKiHgoQ9XbKDa5fQh+lt5yNXSr8Quyqo9JjEB9rkS
sccuKOux501UsXx8x1k5Ly5rXKfT2v1F5/M8p2jQqserltVISxWDcRYSwbvGUPuDcv+M9X2Y5+J1
JMVO/40XZdZ+eIYGumYyECplPsfmm6jbZyz6ZW/d3QjVHFCifNTcrxkVTQS3MIE2B92cAmpI31hx
VizDCXjkHllr/TSqd5RM27kWuMd5nrvbFM0iLeH/yevLguPGSvK/PWHO13+IW1Ut4jeRWUj0fCDM
wQYYq44yl96rnzpnIkEeTG3c8pVPDLZjOKPPPIMQuyVWtVMlSl5vhiYCY4ubmE2kSBxFChWj+ej5
FZoBvxMSBVF9JOjwMgifVpLMmzRB+JCvo9Ba1D/rkDxeiTKuk+0tc780OusEzefVtHW+/KJB5Ooy
QSyoFz64+whmKlJiSzdrCGahoHocbJ4ybyrH/O9oO8dPjKTCR5P6wBUdIQ4CACFizVM7XvzX/AUo
V5CLFLyj10lQSgJ7k/UmHi2oXIfAY3nJoLNvP7G/IfMm5b60PGZBegvn9wYFRDeYToUpCROe+fen
wkW2eWwGRPwGXWRqupDcLWNHKD+kAOPv2pgsbEVHnHS2IA0KOhLpsnt7tA+DrFTrAO+IhYx0HV8S
wjJiWPDaV3IbAHzi8cKDaOEPTU/aeZsMX+92Ef1VIeC1IV9Gv6CSkUsqmO72SdSzgsCjb3abauwr
xNdwzjGSU/Lwo/sdQHbuf9IHhLwOvTEdbfd6+FzY+TNHgNfj8HyW39/8pKDFsENK5bFLmtYXglHw
FMCVBhM2/PIXi3f0EJ3gQSOR3GLo0q7RUIG/xShwKWmOemrg0Esg0Y1WIM+MD6GW/sejLGbFo5Pa
PXDOmzS9/EGQujT2QWj6n0PPvqS/PG/83KKUKFaFlGkRY+/CT0bno2uCcQfi1Pk1oqYLfMQNR2uS
0JaAtN27cKLFCn227+OzPSTqyUE/l3/SSJKmK61CR8uOFGwgJ8DWjIfZbogbctpVSmXMtp4qjFbR
In6TNVl2EAAwd5ZmL86+1oBbKxCV9ZHWCoCooGFt5Lyl5LblbUdvW2JdS4U46545jfGvvg5qroiD
6DY2/CCl9Tlf/qKjrJJw9EzfAXSi3FufY6Hea2WFIWAfvQDJFnbc3V7vHM3apQ7EnUii2fD/s5Qo
JkKVZBgjI9gKfstoXxrKzSuz8lKiC2Gj9j/wWYCpoItlc1EzDgG/n7wIbw/Jy66sNWYMfFF6yhZn
Ie//Fw7DodK2N5VoouQ31wAwnpmjfoqlHO48RQM3QO7GQH68bI2OHpEkSQehcmf8GnXXSlLXTLaC
uWXQzVRX/DU4f3kNrl6/D58HK4fsdgCZVVZ1k6FdG5nkMIxed2Cu/nTjxfbF2FAfVhsUA3XdR/0W
T6O8Vh0UpNyPwX9IOoMmMntrwrV//QT42+pvDwiIlI97OxT0R3EvPIQ0xkMmadadg6iBTz5nkUhA
Bx0SImI4F45Eda/ui9tylHZ3/vtLWEwgba/IajDmZlNSxtzAy+RkcgDQkA4+h6lPprszX6rdx6OI
LhzmIk8+nIqOhGIg5fwihglo3ebsTxuHbjfQ97/nJbAmWsF/1que+zU26UpumxAwpEmS+B8dW+M9
JH5a3UC5ZXYaDUgYVNON43alcc7hQUwPGPdcSzpPZ6vWek7RpBaX6F2mZ38Ts7QACzuRf9D5eXn1
cYPSDQCxmfzwSJ8TdwV+LIG7E2ZFUTA68seUYPdgm5bWZ6+EIzBhQ9185Xv5Atxt2zRhOQgTEEkp
TSPUvTRxL+j3oEp6V/NVGmD8rVbz0j/FloI/Ew610Gx7TUSNWmu0Cx2LDlKqj/bFaFWFCVRY5aDO
YS9SKbHwX4D8qiraKGJHF8wYa/gqHJahyr/DRVzKschRAD+sfKFKu4uDOi4Bn1rFxtsxFzqoOptp
97vFxRGfWPjZnrfYSrIylCDuNxCyTc0LxLKTZls9Hjl5In1RM4RIpql9HYkrcR1MTMVHT36McGz8
y3gtJpuiJ4GQrQzPsarox4gaCvyRtEAUfORalI0ScYgI+UZgRJcUwZZMsfYFEjHGHuEu2RhYto+K
PYW7vS5k/df6mTrELabgqq7bpswrOq0o+zcJcRrR7tgJRNjCiS4r9Twaocmj0XBEyRawNR987UWS
Xr+2pCqp6gfUGL7Ns6zdJxOV8jsj8zI/x0Rq0iImBBwmnNZx0KWE+pYAcxgYu6U4qNPAqY0ndV1d
BXqWmfo/udP1S7gnFnY+SG9a5C12p0LFwKpLEFEs7uqFXLFREKjbDJFFmRDvZOGr9JVCO9rR5pZE
xu63cdnLK0KOBhoToIWPqP18noPz5OFn5a+XZTEdL9ruEmheq7PDNi5N6cbGOw7ZgR1yDInHRdg/
M4EJrkWy9RCW7LmLFhR4jS1ZqYchyvEjADDOxUGw5mcFxNknzu3cAlUbyGYIQ/SneihJ+AL4rK60
doYiqR1Kt/eax0siII3P5FHwY10HGHHkip53yQuEUZ9u/lf6eBkq3QUCSj+7JL5U3olsra8xr4zy
dLPtr1NvVpO4mzNMVtgl/ZKckXIu1tNc3BfJ+Iu5iv5PW9OeOtLGI5PK1Wubw/1I8gHMvnafXjoZ
KUFMwUD2ZNPzWIvAVdnPva+ItZ//JHT2KqVJay1OZLhuYFRpfhM1/Y91mOP3k91NqUbYEFG516tJ
r3GSlKnUjOhUNBhzbF2Q6PRytYXXzogjiqQKFxpLhu3ErNKh4Y78FK0V3btFSJyRxxENL+uIES7q
59u+b3yveqD1H9jFLXjd0htfRIGcUVIZo2kxtqdR0At9jJoNSLczy9D7zuYIZwVq00Dekc7a1Kk2
SDhiQ6jaVHaREJG0oC0Z5Foi2CJtgzZp92Vn7EE5JU14N7G955BrMmu3ShN3VeksfZ/KW528u8PI
nxEoie8/euckubAIN/ebhBXS5Rlr1d2y9sWnf31eOtOLG4HPJrfXOmV72+jfo9i7W6pEATPi3RD3
kdIwNueAmphq640ZgGoF+kZl3v3tiuEtwE2Xy4jMD5qkEEtRxm2RGH6ZF3Rvo3R9on8u4jATy06E
20s6LEU4ypMFeMTGlrPLoL7Pa9fW/q9nUMNqJQBRua8kcsKbv4rYz8hFuYDB5z6luifDYsy8VuJ/
W2Qw1IfvHAwpXi4c/WbaCe443RJZqRwSviPlaDHK4IVRd1vFBZVODH5ff2VCLL+Q9TQzcORTgYNI
9sUz89wJuqdrimI4CPbvE37MWy92NzP/Z/imkNM3FXJaUmcJrXRZE37IWniaIKSjG6VRFmpYsuuV
XbpNR+DsEiUqjzoGo6AVjehUu2XKxl8XMw4JxUTKkS+6emGus3UjkbOCZRO4QCRJNEPhBRU9wCo4
Bj4Fi059xqlVtq/RBcTgaWJlb1VnHVI7FCPR2kyWUlZVfRjsfGwHoMMtHDQHxEzHny7k+2j6EsfM
p9d4yj7jb27b/NI4uZMkpKVH11L8s/PXaa2hkdULuc55Lf3u7+AAY2LAloFw65Ihw8ma//kwG98T
HfEXaRxDgTsWivIM9+wpG5w5mjwV3FDM5A/de2KL9Z7JFLCJhlzgWhQ74K3CHFqbIX4BVFJ+Sh77
7U3RM1yNvwXpTecYc6JWhiZBnyz1e5tIhGq79w315v3OmH+pXRpxuTRQiZAkZxnWxUX5rqd8B1pu
mAnn8Hx5xqU1J5HdpUjYhfEV1Rmaatd0aSXnyqUm3jM3L1RUdObHMBB5gpxxpdzCrkcARvgUf1QS
PvwehxkDNK7zrJiLsZyYmnm/tUc6kP2fthZrH/iFAqBMpEjuk5AAUI5ZA95am8T+SUqeThukxhBE
Dv66bWXnIUKNOw0NHfl4SUajXPFQX/74BBhXQoI9wc6wlCaDK/0V027dKYBj1UNRgeW+jiz8K2h7
xGUhOob9ppja+sATDzsgMhZ5O+zSimFVUHc3vwlXKD9IVcdFY1k1xYLGfOtyakb5HC/lVzsRYP0A
577S7CYh7g4y09uIEGVAa+mK7See/Hq+b+r8hkZSDwaYl/benOyiRllpPVOHYLFMXy8kUWix4xZF
WeiceFW8egMetXtnapycLTSTS27SCTGBKkcqkUJYCCY5sUwcSAlLTnbL5VegqwuKemoJvzeNvend
UG9VmSEOkm+ZIn7q+iCnY24T1R7bPpJ5CSmra0zMA4izuPJj3BgvZ0CY4mZDqWGJiDEqBfIF37Rq
L5vhTVJwh+JN3hFI4JQhL+NJDiqfhVvQuLDmLw0UHC4oe0meMvs2TtHv74HJH1oVoOavTiOXTp/m
VbGFL+jA1BYza9sqL94iKB66lSi9PrD/axUp6ZRu3wNra3eDkNI+6w3RZQbI/3U+6GYTDJ8jOFq6
7CF2l6Ex2PSmlKWMP+BURhk2v5mBgCfRqRJtrIJLc8QeVkeY7FTauJrs7zLpzQgZFA5RCoE/m+Al
YOwlU90+iLIJ0LoCAa6qMniDNVXqkFHgMOnNZXnBiaHdP7/AYBbxGNQyp6yaEjLTbKpBhBvtE++H
Bf1PlyyDcDaY3uTy4i1euV61+PatD/9ub7eYVLKw9PGixyq7/HdVZ6bAeX1bR+ICF5/SgYntYT0Q
9yq9JNGx3/d+ENnYcKBUprouQ2WEx2+YxlyRS4e54qYb/v065XrCcHxo6rihwO425/8n2a1ZPjYa
xdy+uxtN4iekTEteVww4LGc3J5dmALxf/+j/8w3cWG8fYuBRjft4flkRT3x9Kca/y/wEzdvM/Na9
Ue/H8YhBTqiMLphNzbpL+GsJxhu9+CVRzEkXcCC5GelIIO5gGGmCRqJF02QHVb7OnySchInhqv0E
2T9Clu7jPCc2c++gBFpuPMwhPv9uWksazk9zzk+eNuQ7ABhQsG35XRqNINhCFH3GEbnE8NJiFWwN
nV3AD4G/fEa6vdW2vBPGvBawR04SuMI/lH3XL6FwvN46kFxaReAfpez21dQV218sdTVGMganURvj
9pyiNPK3pRxTSKKWwqvMNiTXPwlosaqoAglMUDBUt6MxcuBUUn3/HxJnPbz424oipVBEbPDjeT/a
dMLcjRriRMJeYic64Od/IKgEI83CbYpkP5+Vspbhvy2gUSBdCSgdZarlQS4XAQbnqFK6w9wEVL8S
216NeXXqaAQIpz1zYcegacr1Xf5rL5Titj3Bp/YX+YCrKmgWyOaw40VEWnnsNsQEH4y1JdxG/cAz
zHz3qP24sExpZnVzNKr5WtU3tq2J9Fqp83yaK61mvVplRCtFvT6W4m+l0aER9/FUMgcMk3l5KoEZ
PidbODqUzMmvleo8QJQcIfos2O219QhvuKQFZ2XIfZvGPQ0zXLri1bKE3HwKniDQ8q/D6AyL+5mi
QJ7yrLC/bBGBriqVhIuB3/sdfdQBFtqV3m/Eda3/J7FqHYuzUWjDE6oLtdGvfHKxJOUZQ5GYCUd/
/o33qv3KpZGh7ioF6CZyOwSPe0b1D4iCb7B7bg+g9ZmdwgyOHcgzfS9IMsGtaxJqed8gXAEnLVfG
hzx6MJW9CkuKsoYnMv0fPtcOzz6G0eT8U8aE2l/6/HomSuPB4i11xUeTV8pAKKl65iFz0qQgN3b6
BGklb3HPz0eHbf/SvCMCXS5GoWZAkKsg2ggLUjjKJVo3uICKriVfnCC0o8S4uumFvtE8lpLBtL7P
rv5d7vdEDnNOQb13R0zkeWhbaeB5aE7hm5JTVte9UEIvwq3IoHzreGO3Bzc2UMu9vbgAM62wouCN
oJMp7kLYeRKBBfYMeBwXB616tFJvCWMqxWssHCd+gyjsR6eiNuijFQo3FMerF7TxHMf4uAoYgkyc
t1Fo3kGsVpNWe77Er4g3kuVCUQZE2jAVBwjeHLZc2SBArRL5ZaYrmSY/j7yRxYqZYFsXlK8anApA
7o784lJb7+sdWbIThpP14DPQqDwQ08Z42dMWX66zdRdCATDf2Tg9s14wvJhWeTjMJhlaqWQ4pcl/
dKUQ+KJSIOs3Jh5jlLvmhrs+98rylXwoXBZifMmc5aF9R5zmetyENyaB6Hyf+4294AAFSbRIsJQ3
KmwNhfQ132OOHm9iCTQaMz1iUPjYy2VKFfgoQYe/oOlombzvnIHGdQWIsBy1Zc91h0Pptq0EDekE
YV0f77WvgizAfga9iHK2Dp8bndD7seibEsvmpVBkcZDlkcCF6soAJwiFK1rJNZ9/h9HKWuOgrT71
pQJNpLpIMBRPBdcpLMLxyURd52mae4C0VPSWLQWqkHi93mRjJ8nZM2SMaDbu268OaUKoIPmkO5ZD
+QuEBJtFXt5rPEW0GeEwvzpWzZ4ZVMDjDNGUwZg3plGvUkDVQXtdilotRCnLArC8stWYxVK7e59L
KmXzxIOvdxkcDqENZk7xa6WF4X1Mnp6k6JVRZcMaFy0mgJBL2TdIXO69bT7K3BDC/5xsY4PzmU5t
AaItnBXtl/hfTGEpf08bvfhiBh8nmAR5rMPONG+el4HAr9SDXfeTq850wkTOvsY22YoMypNKHJSc
AfOWyHEnTztipso19nOHTbbAwa3g0uPECFLiP2RubFvXJy8TYeOI8eZfJ/uPvZBisN08KTb5xZuP
OnakgvoVXgwrPUyghzT5kGUkA45Rxo4b0JI+klSxWohnRUHv1qqXakQk00F5wfNdJTHA5xVN1z7f
aUjwcyhtRNi/SDn4BGzUeILwRKTntf3omHNa2c1wEnL1PfTX5r7OBpAqiQWmg6w2FiZ9TSr6Efpm
NvysrcouBsFxnsguF9ceO0kcMsR1AQMnw4VeqrJM9augqYHlajOTew6ySjwCS07ZxczBqxajKe8U
2wS4qoNBz/ml44/cLJX3SXLLco0w9zKkRtBB64475qWX1XjSr3sdcdcZZsml9NWzEAtTOLRE5uAg
LyQtkGmZEE/0cHKCzwLa0W6+PgeTdsssiKfYw9+5aNOS7PZQGpGZn/octN/5qrXkFhYBb+hCgkGy
FbXHAWU5JufC6fZp/S5j1tO5BEILSJAoSnFPB7uocVFlmwvyyH6z/gPzD0gXN4Zs/R6h+rMaLTz8
UtoKZyhFcanH1+ilc36pZIlOQrvTa64A+yJxA1CcFCm8jBl6zWjMCI3s3aycgFTaOkrulqw4Z7PP
zMgUpYNDg1d+mIkzpbRFn5NhuXYlzAQN0eP5Q+3Jn6ldvK9OcEK0uCUFltqJWbwkIxjgdJxCf5wI
13z5VE+TH0XIGgRqeQHBOpxWNK4KytesBkvnwm23EfFzR1HDtK7xjP5b6aQNXa6q2IpEYhdmPBAJ
DTGMDzU2IUJXyDHOemy1xbdIgTMzLy4PWWdtLRXEjUtHGA0oGAkBCumLe3yGJlIdie5Pb5iXdP0D
/hXKhTdNHLwJZfJ3YGeqK+lscjdaxm2AjCxsvD5ba/+xnfjvWrcunO3DolLit7mx4yTjurtw92cE
sEND9UV8Fx+wYV5kTNFEI/DeoLu0PoQ9IqxLCqJkSiyPFwaVEF26Vko3Hs43CLEp9NzVyS//Xgsx
pXAsqZ7KbvbxtZ4XV+zAUbQqAKvZrLB4cZX6sdt7xmcXLqo5WgpnrhzpK7zadL7sD6BcLa9mEVzj
4D06fWjtnzyqL3O39MeOL15l+OuywbYesC+EC3UDWj6T52ZGte/Mrqr5V1pH7jSeVCyRC8bhKr/r
IuRjMZoadTFizDZ9q3xKopr9nBaxb42+lwbUPG3EVgsY9rKW0y2KwYKrA1eziu5r4lei6vtfg26E
1bH/+F/l5ckBzSkGbaOJosgrh9hfTFoVEhBQULdVnyvBP7HBQFQBuijjtT9E9Nz4FVUHfq+gM7DV
MM9UJXVcWNacvIEY4FcqHFyuGxv1LvLPN8lPUDwudUkSRZs3KsJQJZYCzHm+laE1QPyZ7io6dwXk
LExZUpBizM0DoH1qc1xSG3xLwb27J6RjWicX3VlgAFTdNBsGOe1TV3wFYs3lZYJ1x0N98IArK9Fp
ER0E7iJ7JZPUhwRsctKILLEbw4ECLX0VCDQQeBdOsd74iV3dOERz2D4ij/7XpIUQsv1R8Z8XSkX4
kctI3t+kQOKKcT37bSMCLnZ6PO/czHaPI4eOhgnP4t8hH+2fSvBuaJm3NS8PI+Wk3AcxqlFVefdc
dhl+l9yTragKE2YiW9uxO3VhMDtqwNb326eMbW2YhJZTKi1WXqLaZsoGUr6EEKO0ydAL9OhP7+zO
sV1KGs0giz+/8fqpGBjX5lL3sr88rUSNp0bzlRGsWfuDXQrkHddcITb4lhPceyWiC37IvC9pESxi
3pNYRyPqDkUMSJW1j1r3VfIHuNBTjtF+SKjRQCjRCHZ1u1MHBj7zBZGSDq8DDgAUFt9z4ZgYbf6e
IUduBhHDmGwNut6/RfNsKVB54e479fC/xogU4PLHPuAaT1Yfu3gNo1lSD5rtABtaeZieUdZY7kw+
0rFx69TVBAjGy/WmMpek5IrzZB2f00cs6S41XnbkXbAV7oRmNDrCnAQkzSRbPMdaWecZvtrzwKzF
aNplp+5rDGVxLqJjqCyNTYgINfgq477gxpsH4I5/1hLpr0PIzpCKvKDmQbUnUDx0dRlyXZ3UDOy6
utlbPoNvLr2tm9Wpgz4Q1l5AA0JubA/jr1t/I/tg/TfdZFW5T2jRyy2F1GG2hx6NQY89jTOPPQjI
mbSS+x2QYBz/C/wvxJPWimeZgoKFzsw65VDZlnfY68ZIksPMvvSZlNwWgqRoXf6t0Y1iE6c2AAjt
2oE6u2uzDTaUxmmuCKOWyjfmHeKud9YcjWCOcl7DxiYVSKQjjop/9P3EUREs7yiV9E9O1KFx0VnC
JWEVnPElZM7dJdtNB/EQFt6UyvLWcXIr+x4LjZFojh1GMWTD0Z0NbL6cAK/tDeogsbt8b3fif7UA
t/AKXVHeCyfaZ498vpVrg/YpFtUeCKyv3QX9qjL6Wj9tOCDUr6Hg88sV4HByTSmvm8M2JyLkyj5c
gqFCye20for4MCaPUb8WnmpKwWLaRXs1nr/u4GAQ7GDnODOsICba/aG9Eq97+ClXdHXqViIXOVHn
O2EW7B16RQsbGxxbFr/AvuHk7iIDluePuGui0MA+5hBf4B7RTSpf3PIIfMr0iGn90Ifpj7DwkbIU
uW/5lLB2oneOwWCj3NuB3V0kYO3HsKcDUAlU3lscRSzcZ+SFb3jTvHBkuDzFRszd27vbNrYO+4fH
GuI0KTr00CVI495HCy8JJ/u+MLL0jPc+D1uTAeuqu31syA2wTy/oCtsEPp4MKCcwnQo9/vjz2eD5
N3g5j8ii5mkWRTGkkRGxjYpxdJTm64TcqDPm70Af+Dgj2lNg+FG+ICv96DS5xIQI75LLBIFWeyFz
f8rZTT1lNRLdf3O9U6I31k1FaGXCjoZ2qZzhJy7a+FPGaLpavYnX2LaKmaj6E3TYjWNWJaD9Nux+
5wK0RdsoT4BcIPFOFLSULZYc8kkLo9aie4lyze55yCuPTESEKp6xvvZ3MOjo5hIIXgLUQh1aq4Gh
63XXJHyWSrAlMCY7ugvHrvKXA52oNT9dMIgpMe/o4pCKd6njmrGUvChxHwCaEwb8wm2gup8ptoIt
dYu4eS4xzAphoLbUiT5vmeeilVOJu6bkY7wAIqDgLPg3QsV/FO4JxXnhOxFT4o/WWO9jGz4IoIDq
TM35DJ1yfVeoFgKCTiHVvmKQXoGxXxSAjlZw01h71kOh9Tm5bG8xkSN4iqKjr9BWQqYg/7w5S/Cc
nWqY7eVb69IdzmsfMRnaANUX1dKGx47bXzFCUVOVmViWHK4tgfBnAZzS0MHYkqvRtKT938LV9ur5
JSuSBq1m6ritOXdi7MRJ2U3Lg/Q0TBhnj7GHxzvYL/QcO8u3UHkF8s5CRLIrA17K+hf4gD+WEzZw
J36dy52aLPVIlZ7G2kPoTyDA8+sswsgMiRwtra+6P8sJs3AdcStHDEd6V6rr+KJnSJdIA7McQquz
o49i6HLeGSWE3Gvv44kPM26UlaggT7VUEpEob9UKSRNGfbmqOG1a+1XoC84wG4qEOvvnR+0zBg/W
0DIR03dUE1kTpIbLoJFAlbqiQk2NrRYLJ1Mva5LWo8rCZX2sxS/FII+q5NHt/ZoDxPR9dWLPdgMN
jXYiiX6wwI9uDx/+dDVN2sQtFKRz3HyPFmGd98AEjfMcEbp6tHsNSi9GaGt0dFDfTpQUzLbv8YM8
VbwhKms//ajweKeZjrJsh/uuL/v+5cF93BoaJ54PcrZD7jVCzAmn/bzE74A30bLY/F9NUko5Nudq
92/3bzOsfhluItDxWmyktr+vuxzrykmog8gPOz3Q989NOCSpQT2ZIUJ5NkAacRy6DdNtU+ZfBssf
6gkyIG2eQ1KDaUbX7jN+zeuzvwhAZKbNu5kV0fbL88x2eascfoPGC5jZmNQrPgnOMdATDlzIPBLa
b/MIdupCCb2JSLALioAO/LH+PTeUV2ZSdOAxH6WAd+vpGRzANLZ8C7yx6TDQPVrCk2w49PWLH8r3
xy8b7FJrloAhf1ofmZOVDvJrGzgIQzrfrFLYXfCmYwMQGGaQ00bdbBEbdqjRlFufLn9KTSFqJNzU
wQGd6iOI9Hm5fmYs3J1ESsPXCoftgaLuQHM++gl93k9qryV+ChAZT2qRrQESUt1D5DwI1MiUQ6T/
q4KWBRVhuSRGuCiVYwMWjsT5k3eK+R11a7IotQFN2EeB2JBIIYmuqZy+Jr5LVDVCaw45fUqeU+Oe
G3NRbqHkS426AX9Z73vEOvHdn2ISHl1pwahYYWp5yZ5wigWXGCK9ZekWVs47nyC0z7dHQjyc8L2c
lMxqb1yeStthU+BR+yHUckVBINaO9k5IHBlTo4uPURltZujV7e+HfVs4IBAZCAIka1T7jd7a11ky
ofkO1QFSvtaZrTOxBgYhg4N0BXYaFFGLWunI2qOMK1EduMV2o/k1NLkmdciMm/PW0JkfxgyvzKHz
G348wdl+x/APTwGXxIZs6oGO2WlQUQ6ciALgdgM7BVBxzm7sX51sG5dfHRkcGjlW/iWv7PUFFLmx
D1oqphZ0xlrEjuMa6AIz9Gg5ekF56PFkQhwcYP0ajw1bZFUmEZ6lU/Dqh7UoYbey1PDj19F4rdD6
gHoqwmtFbiLgiK42dycAtcA+jGQZb4Cv4QmY1w61TEFW2DTqM7F9XkVcfkV6u29J/yC1UzGa11tF
OAH0WesAgE8KdBrCNUaibexKPvLAbNi8Az/sZjkFfAc83PwT/509ur+x5N3rqX3WNvm6LwB+u77q
UmViuwLWIqT8ExpvwnkCqDLIDqZPbjqEiYPfd7/ygSVsLd/s5LF0/mrytxEeZp4mIRWxTV8FRT1V
H1ld0FO/g+7znQimZB7zoJbgb/wc0mMKXPr3mVtOzvx1u+EuGPctqawhaLLqpxbMD/PwtZDZRzCB
+7fjh9nyLJH+kMjk/aiRxAztyBYagrIXbxSYnLgJkifhtq8XrzHnD4oG1/0mZ8aNTpMrDglqNJCK
j5JE4tMD48VAnrkVt8V7CiS8vWlZPhMUEURh/R/UuSIJcOn2twbwoct3jpy1m63sYyrQNzT5fveI
AEe3o8jyxMNsykIE8J9vo6PXY1pR0DhWKr9ZQvYpxPGcPJVS55jeYilCYq3V49WVdDrei30FVN2P
r/wrP2hVKFocJbDSjszLeBKEMdxJDDJwC/KkYa2VWhdIfc1K7B1Xwo+ouwaaUTgj02J+U958Snl6
4wrVHwHp540MpPUbo3ZO/bB2YReZZEa86rG7GDh5s8ytwoo1SjeCLvoZfDLVnPj3nTbnt4XAYNnE
PvwzErzc7ijrO50zLRyOZaZ8hIqBIjVt8C5nWP7d+clKICvfiC+DHJuVWgt3H0RkAuDyymAurHWo
oQ/GYsSBi1BMvfLGlepWidXytuGw3PdCCLk3RW2Uw8vBQu5E13Z+UFbLeq65UfkocyKibxQAy1Ip
7L4mETyrkWGnngrCX04YGsLIOVTu02Y5ZZkQaK3B7oX5tLuiPc+Wc+WsszT1+gMA7AoAgFEashwc
1ylYu98JFXNOdYdZnyrCquDGwQi4MzmKjzuV+jsWzEhITL2Yg6jyWvD7k/sxS1JjjMqMl8O9B5Se
nDi50LmdYLRR38WDNVnfTYafkePp9lx+O5PVC31h9G9Kd2tLN+bralLUacx4nj87dPUF80vseDmL
iPhZIlrVXSO/UVJtqeTFU1icVpl7b59onhyk9SXg0EKS5GHIEU3EDwy94YvsDwaNzLw39oLwpvWz
lIu9b8iGuOy462qR6ETn8GnSsgdlSyDFD73cUzFDELwt07iB6ef30InYFc0uWiBOecHNuwszDXgZ
rtKA9zJOaIrZzpzuILRwLwD0zdbuw/fppYhIr9DXYNXTakdOnvsYz9/Z4jw9ZLLlIbmDbjFIrH9i
d+uhxaSE77lZM/j62+PLcjsx9iUhlEkSz42U4oe8fSOoOUaqwUJD5iqFHY8EA43uF/82sZveJGzl
GOj+8byEZdGxwTnOk1aCW30riRQZkhW5PWGFZyMMQwpg4CIXYLCXOS9SFWtCqwBKcr6YydNoWNOm
8vyXwHFJBY6ZWrUqR2OhjjKXN8DZB7S1bGLzzrFfjty3V7bqLoNsWPjfkDtNirft5qzoPuqV7gBf
BTbWA6u3HFMFcFzudbIVxEYzoqnBNsi5rQh8dXs7acekBuCJcUBqbpQGklkBmiVR9EJPivpuZ6wP
0eyrXALUTxB/ZYvCypzXF7cBL6fInAo8bWu3b9pE7aM49pLrEPdmjsrSMn/UuoIrIVu5mQG4DohP
LUYwrJe32HzGOv2NsG6/HDdpq6Pd66QVSr6IiQpaiVA5QCkJJTCjqHc4ciOl90U9Hp0ZQVDFTYCy
FeZ5k9DI02XIIbh28n76ViR8MHMupKDz5/Cwg/1YgUQs00gq77qBbSOaY+s4akXPKvD0oQCfqND9
V5xVLZ9RKSUNd5diluARU8osDE0/54q8AEcNjL1UBwOuoFe0SZQ1VPH42wTF31JSVagu1FefLSc8
dR8CQvx9+POXd3x3D7R2hl7LzqJhLTKK1WWSfIxfxAfC5Lbn7fbzs8YiuTS467RTMVHN/ADzopP/
v0QeyrxeMVUu70nt/ZWq1z4KwGmBJxNljFEf9Z7hGykBO2OoaPA7ZMFB6x6KpuroA8RkijZ1mR2i
FvNxYEKZAnaQ7R7LZclovs7xviq4HrtklgGqayM/YCfWcMxvGy8/M4uWdwExrmsTseHPJ8o3T/V/
Ybs6t96Qysz3MMvcvDgtL5ffWIKzoOnt3pqPmPv8LOokIwFCXkq3axuh0ud5K5w7ArYGiGF8CUon
BAdlMcYm/VphRABQuJ5GHUIwoL0llrVejH/fF9Nqd2EgXvCG27AwXj1t/dvWcsc6LO47K2UAvo8h
Wj6wzaCJXuynsfHuybZSkHsnthq6BuqLhwZXBEuJpBCB/exT+s5ClGiG5DU31UyvhqfnWJ9KhVdQ
ywwBFpERbjqPunRVp/wNYaX1fY5LioSHUeqHIU6EQqBGLUIq6ynqH3UukNLkf8eSNFU9WejyMffI
9vQsJK+50YtxrMIzYgaRrupefxHInkblkm+ExC0jIjzXs3mzFFLqx0J6PMMsa6zmGteNdUZJXMku
SAO/yyuHaB2YgGYeB0KpCUcw22Ut3WFCsr0ZUd7WNiqYjye1owKP14hJt+3AiWb0v5/Qy7v3StXQ
gp08m+nRMS5VlpGKLlljzIWwRIQzkcx2t6BmNbu/Fn7meIrOwMtdvjnFU6OvNlBObH03NXCfvFk7
8rWSYdqLguqo2XLbn040L2tp1FedmkPxDdnwLj+Je8VMoT537ETGBKdD2wl7ajDB9y27fG5SZG/u
uFH6q+lf1vXVrzSx1s/Nin9oI4gq4gZpvFbZRU0UIORBm7k9ibdxsThII4hFU1WAtXB97QnpIUtU
lVmnWSerF9eG79ptvDNJWnrJznraNnHrvFK15bRZE/eV9KH5XW+WvQ2Vap49PN1L1fXhoMJpLbFm
EV6s0u5YNJFZ7mZ209GhnYoT7HjOZQvjrY26OvQ4RRmGzFIABuCNuEQ+gmeRLKiG0CdMKC4rPEJS
5OEKzjLpGgGNb22Qtoq1yihQEC9/4qfe2xwZ/tOXIrD+Eqeoll1VrPDbBorfI9Ia5c7Zz2gMhbDc
Bp/DCAnn4M21P2Tt0U+vHp0zIXeHqMLkO6bHQ4s2HDYrAJOKKWpCy+ritBvXR4xf3tynHJt4y+jp
ov78/0LV3vggcW2fCq77qxfwQ0otlgmxNtkSEVKHjXo9QDDZ1KBapSrbnlvw5rTm3X94+Dmw6jSa
ewzvOVwkNp2+3NzoSygaQVlAE6VaOHO3DYbq0ke+dutGx6QBhpi+ExjdsXoRVikisXNVcH44j7BZ
VeAd5vNnuA7OBCRak1uJxTv9NQrd0jCLz7N4n2Y0DTR0jtzD2UNmf/l/cR096RCNR04CryX0cXhA
CduBip8s/zFlOJMIr0vpUsmU293Ar5a7MCHU6rgosORwldDnjmBxTKyQnY4yyLSEeQz0s/5hCHZy
WoksZXWWEC6Cl7CT13l2ud2/6/8sYS9/1SYLhoeT0hEbR6nyUm1rEazTTXw5ZMeszAOyTjylCEhr
apGsAb5OTRc/zxPeEXy7E+vwB3JkJf7+G6yRo1oz2UQsLqk+7Fvlu0SGM5SXUPdvyUNRo4Hi0u8U
IouWFhGh6Kqa1ExK3zOH/tAydG3LxduXvWNVkJUZRGeXniTponFwluhFbEaCZFHFaYdv0LDQvkYt
b5MGajLqA9uueo3G8h3h9RrH9HExMyXe7mhcYtt+3OCg8nnuh9QOYQMqtaCYOIzliSd6Lht1kY52
oXL3JFVL6ItNsTlprDEhJLBp0KP6C78pnm9rt0fq7TpOV9OLBw/rMH2wGBG/uar2g7NFWYDpJEfm
JxxSL4sW2dV6BO853reAwiN8wMR0SHIri7rtdHVnrnlClQ3KbFS6uqfLPDnoEcw1C5dUm6EzvCUd
k0T7ADbrFewl0gNFzyLWo4cdztSBJRfT5VoYJkF4I3igiyVIv4kDtbTZd2c1IRc62MpqqsYfSkKE
K0ehU8DKunc4FWl8xYYhUfSTHD7q8sYNI1aLjpvNNLZXDND7Sw1tBBnGXEgtdYpExU1k0zy6T5N5
vSexBdD7IDYAJ46T5VBec5sJUvakMzuIc+x2baJtf4MclTdESfw41cRGJnDvum0x+T2JpQcyhRRr
qUWCco/6Mt/8h8JGQ3KKEG97HEVfE7LZw1TFV3MVvCQrXOt8Q4NGPTHXChu4PKfQYWwrakqnxMcM
E6JztrEsXGzDW4Dh0VFZZTYU4eJumeJMxktaQ6lLbAo3aiA66hU9LsqoblJqF5hMHxPDPRbzvdMH
iAsNFzZZGoW5+SReTxg2LiyiCWLzee7LQAtyHAZ+AfO34B39RMT20ZE7+wN0XBwBBVgzei4B73RL
B+b+gmI60Sg2EqKn+CbMyA2k/UwQqO7ysqb7s5kvtl+yNI08jhRjlvGN9nE3747REpNwZv3HSH0j
W1qq7GRQ0SZNOSDNq6OqT30dziAmy+O7268Uf2w+0KaPo50Ir9IH/ZRfygSEBMnxRH8WH6XiLq67
gedZSGGUwBDgO9EaRb9b22zCVIX2br0CecbnV78ycCHP4qeclS6JeCvJV+6QBktbMAgehISYBWcS
w3ZeuQsOiHpPifSHqklwrL3N+i7NMJp7bN6QUQ0n/2coZEm4Jsfgpre0UbBFbbnaATC4iY0zKa53
hLfJcF61JvHQQzAzKgt+iVyQz7eGX35G5s49KB9Qvw0esc9R47/mahA38FxCusgNxDxHk1ziG0xa
tNPg6K34aVWiPEqRFk2av0WaxEWblqP0RahSFi5AEJXMUedp+ZO0H550r2DjQnhOWfFesjodmOw3
abp9BX0eyRX8uxVomviSV0iy2aYkqvNLKMtNGNAyOXxAuOzv+szO8yf5b3S3zhDmS/g4jx1FA9a8
0dZuJXHsKt6Pi3nvjVoKKTDJn6O9izgMuhs81YE0Pj4Hv0DRLUdxhkREjbsMLcTrSMwPO98tNUY0
QeyD2KdbKLyvdF9FzWdR3/VveOrkcvkdyJlkyq7bsj0Fj9uQN87bsk9AWyhdJXUnAjo2TxFC+1FK
exW4Fq3LbIXlVs/f2wcBXa0wFofqa8dKX+v5vU29k66vH+/k7FMjdOWaisGgNkeCL6r9jrwIXTrZ
8ULHkN0kvU3Ld9m3bVOdk5R9tj0XmGnwGiy/dkQ3cF5gyM/qJFNaZv31QYQQNxJLMUulpRcDDE9Z
yHuLlC3ki3mYOXw3XV8SnS7CydronsTsdiBQjAz0daa0+gACv2RhRMDQ1HLM2pQWRJEPbGnXgpm4
KcfErN6rZqOG464/haVH/clDeyR06PBbENQXPQZOVuYPANvPV3eLvbuaz9mvO+UgNT6wZR/jbgQR
72UrSDKQELGbhFOSPGAEXs5cBp5zfrxJipkk8QWcFBfg3eJmsifQ4dwW5bDGo31oDx7CENwIVY7C
bB6hSmdbgGjB3hyrCnVWhL6lpf57i8R9BCXzhDkJubrP6/LMyqgQSVaVmJQzcAbECCOW1+VQPWRn
XBZaAIrxIlRyW1OzpLt4OLPFuN/RW9W3sLSmKDBKRsJxYQjZhQchKKG8SwiwZOhg0Q8ReyWiSAyy
1x+tCn/Kh/T9H/Bv3X4djCd+i7215A3IXxZGKaUK87RBGLiFID6qgI3Ws8H4YNlYPt7ebyU7Ke4q
F1PtIffkUqTRjYEhMV7Mj59/GeG6692F9C67rDUrReIM1Mtno/v3OqTW1wELuXj2JywdMgVONXnZ
QALgJ7pXW/kiuWfwURUhD6fK5y0hc4IUn34q/pzvx7GE1emBh0MNsmw3tIdULAaTG5+xR+MF5ho0
3/sRtN4kqWOWZ5qkjdyuusxH3trolgwXN4BsLE7qJWNc5bSRUJauHNQsAorToxXi9cI542cOqDDZ
2QpmwcDq4z1sFOXi8/GfNI9GHNsJxgZKBiL53d4L2o/I/bTEsP4Ug45dIsveHVOCNVS+dIvYUp1j
9Rq+AhZoN3oHeHZHkK+RJ07jqhjdpBascWItUClLlhnAousm93CmS7dihV5CoS2JDUZeyXV4VnwW
b3GxCvBLG0aVcKUwHaE/fcxehNlSR3wasI7K4jGzuECCIbB90OY6AsVBOEw3xxvDVmW1bd0pkH0t
gDAFHtKMUxyt7zFrAou+UL5z7hNNYZBtJxEq+qaxYJoFMjIPApwsoBDctB5iFUd18tS2Qup0S0Yr
BAL0OBKDi01NBwW3bYR3KOb4/Hmted1YQJnypbF2U6v+Uvz00Wz8fkGPsnxqfECH50vIgedy03Ns
lvtN6IKl6CtQmIIZNTINJesltTOSp5yaseLkw89hHM2wjIArufWcE7t4le6oZ+6U330P+9cn3OxY
ScRz7a8nY1HgZiT9hrmdcAS1sbn8bIb7q+YuLBstqPuTwCwzon7I9s0By5pNJqX8QDr1ftlf+yY5
37P4/g2MXRN7WKmPJtnqvRvHSA90YIzNDYVRPhyvTSvJLVLdljCDPk1K4Zp5xwLD1rNrnMi2lZKJ
P5Zn7rjqsIOmDkC/yvnbVvk3xnYBUCfN5E6wlwFVA9Abqaahhz95k3gxElhhkCd2xGacQLVFUHMB
vG+S4+di0IAbTvQ9IkooHfm70iy3fBBHTXp4e16s5LsYm+QCVMUSo33A7HwV6c/BAiAkxOwxfqLC
gb6Q8X8pimqzg7OmBGidDc3CnapUN4//IGehbe9WKiwHcIK1g14P/p32cE92FUluBmDOHLWxUR+G
7KBJwY7jmomTNj3SZdMbxOC09X4DgAlALgWnu6RQ7nbdzYdmIyPzR2kWGgOUj7fqq3LVMOAmdtGv
TEIdQOjXOrLB1iAa/Ibm+T0SmcEIh1JAkA3JOmbjNah3QP/KHjeo3MVBTCKB7TUmjUS2X38/RHF3
b4POI9Uic7cduf7Xz9vWHresJO8EGTQotIQi3v4hn21aTtwVIgEs+GdIDLKrUx9HNfrja11qzpcc
hNMt3DIH5o9QhTLxfFG0iB6cSbppw37HAbnBf7ZHpTc/tzLMMrweYuKA48KVAG6SoOVwCS/H3ioD
YyLR4tSwPnBrbqHJ8i3ZoEkeNnJ6dqSI9YagwRzarel1Y3viipMTM6CHbZFFgmqMQZPuYHESYVKx
b8BNInVMQ6wXRWaQUHnLXUbd7j2KPUT0rt/G/J/xRkDDClQS34QvRv/XUEF28Zw4XnNyTr8KQ1pf
SJcahH9olO9m14S8t+38s+GBzJMb3c28MAlAFCdjt+An3mJ1+IT00YnZIdE73sbn2xM0YYvD4V5g
HA2s8CFN/CuaQbNDEYKbqEs9WJVt3gc0A7LOkLnmYPgKHXnaGama2FJdy0E/gGVX9hze4uuac4T6
dVCSPIykwRJ2MZlAfSqj1c8MyRoe7Y8XN/MUa2BT/XCnSMqqp2Z3VpbiVdBk8l58cT2e9Z2Nw2ej
z6454M5gu3GiHxIvq8Hf3LheYICxZ4ZHbBOEC2aBHy7ZkUp0XtBmz/N35upwP+kXg8Iez9mFk70+
6CKWLdvZkbahYzdzIIW1MGzI1USrL6rfsL8ncpk2HwyxrQw+TDtLSIt21mGmmGQQtgN/dfHSAimY
BKsBikDngl+C2yuTjaQvQ4jA5ya9jr7NEesLxGteWcO+lLoCuMQ2bk2rARe1RIyWaY8K1qwf26bl
282mKMY78Vsz24UcsKGoze9r71/01Eg9/G4ELLMwFnu6pqjryxpRCuZeqQVDZQjwqTAUZbx9q1f5
B0onkM57ed+Ov4CGuO9cTu7HyuGvAjNSEafAiXoo2Z+Ppeot4Ewd9RBauSAf6p1Qb0ZDMg73kgtr
ZEO9s9WbMGGx5YYGe4VUte+/VWsm+RoWjcW/jJXFGi2jA+J0ziJN3pJaoXL37Etnf6mLUAT0IP4K
iZTTVsJxtgEpAFeCesqP7jP0lNMAM+8mhdge158qohA3TyDq573WD3Zi82Vu7uWdiWJ14QU8heCH
CdqDi9vztbTyANeSW1MEWuRIp0n2KQRf5KBf/9dAJkDnT6ddFeqQyPwh70x2RZnUkpYfnlMUJkEd
sjprVnZ+TzBh9CFOOq4oPrHMN9zYBxwLCuY1pD2oBcrmUX2dEdsJH4NArjGYLf3HAJ7To/tEoXw3
sky1meSOS+b/Y5MTAUa/wEInjN141Jg/4/q88gd7wNG4GHeW/CN0sEqEhr4fmC53qd5ZuZTlGRBr
4CbJ8KpR2AsuuMmNci2KO6kMmkr4qBQ6KpDYup+ZwJthTb1eufkg/5lQanSlmOeppGwYE0IJ2wIG
qlXGXJ9KwTpTIxyo72LbSg4OFbJlwGdVSm4+YlMgKktE2S7dP1/tE+d5PAblkFvaTFDDsswaa1O4
qbtCIbZlyisDtkvR96EeUmR165QtgNXPArgunOAhUugs5luTtayuoJYEOMBAEiJeWcvCNfc5haGx
4zos4Arr5B60bTWbLR6AdfzVWdJxfKnwWW3GJ8L7lx1HJ3Vf9UMQ12kIVTT4736CgScaExKhuh+e
TjNU5sHTXV7fwy2QfyDMlde/endHIKLcm2IbHDV7WluK6e11fcXmqtair3grz1UrtlaQiFfWhHRP
5bcoJJSDtR4KiGaAsGsfuF+z3uFKXJ439E3TmXzSxRWhHM/fFYVtQTzU7CTgYq+FMvPy3hE+98Ee
DNyQbRCZDZp8XQXPJzjh/vGuLzm3zxmyEU/iaKh3n1KGo0zTqQEVnjo5OUJyoEGDY2rU9SerKun7
kDLvBWW0Kp6cm7K9a0G+vOs7uNXH09aV/DzTK2BNted58M34QLm5xB7GR+08S+eiATfZBiHkHtMj
ofQmjYJnDd+RT9XAEaZ7mnGuMG7Gz8cOpkgdAVXdtDYPJ0R8Jo1UYixU8IiApYQPaw4wk9IagK0F
o90GJuedY0qxouPrrHnKzGLPaas3GqGSdwIYsUjnrvEX2oPiTsdZw1DolYavqay56WXWHhadncVq
GzcWjoklRPPlc3XUT/R7oYP8e17AcJL4Z+f0r+8fApxMsAXGr+S/t833hy4gOOPrZXSiaR7+M6K2
7eLVq8SNuU0EobMAGpRIj9UyrGGBx3HYjQf18FxHW+uhFGljB43cF9naoNge2cpBHxzgQlj+BCFW
JbigfOgYA2Xh/1zInYlsSE9XOtdB6L8d2CRwivLIcfkS+5ZLNbMTekueu38vJzegjRVfBMV1J3n6
yA2PS49XEjGBarOHqgCWApfVCdosESaHhlL0cj48zhSumVWreRwd0PeYHwFx3tCzlHyaFrsiAHyo
AlpeqdS5Ij3WwX7Qvh16H5MtvzF+Qtua/1hanfByBOdzCyi92UYhW1AK/Wk4gf3nwYEWpAZlILqO
501rJTJhQPymXvgZFP7FtJ/ejpxheb0z+ZfZHQUxfmz+IDB6DgeMvgsF304MJ+eNDQN6an5DjP1A
EGjpu25Gmy5e3CRA2OloA3URFp82JfUBIQZzo2HRcNUPGK8/SEruCtK4B9vu6RlhQRjG00QaHbCu
IH/qdqNo2Ijyu3UhCFErXA/y2cKQoomEhUuIglszXx8B9Evhsk5BOwOxpehiP+s7qlI0RwbT3602
VFJSza5841/h4qpVGgkRm7po+oGfhQ6Oz2zYH7BeoEZxMGOlwz+3jVbsxet/L5so6JB9Bcms5R5s
KSmwN0LvXLLjLo8Mh8x2azj7QeNhIJ+mKStC9ysqfVFaBnkbGngvbNZ4zAwPn6i1KSMilLWccpZU
+SEv3wGJGKRNqQWN6u6/2u3rqio+f25D1hQo4Gn1Igj0Z2SzPkSIedrbwb3jjzAv8YlYQSSWtuO/
Pgpj/BrTsvaxq2dbcPwfNDYig2kngvY5JqKTzriCBqVJfFDulkXtX7wWdYyyHlyw3eRBVAYsfmab
esVBiBnYfxPxcB0uNcnpC4c0f9/3nto61KPczi1myVJywtpenPAeQnLfpeA+xSvwfE2C/vjmlik8
x+2axbPTDqYbilJx7jZczBIYKM5oUYOMg2sGAIWzLU6IUxGSBQzDBucWsa6vfUiZe+iNJNaRwGa3
ugW6xxydiBewwMXYrnSNaXObq53J4aCbTbGD2V9DoqEbQx7BNUeGAZKv/u6w7IcWd+wV7JZk4z6w
MSD7vdanL4gjX8VHFLnr49yBhYt14kp4gQC/Z8GYnkm/ziBmPTi96zZkY/ldkA4QTroH2wfiKWWk
Ydt0aCArRexcCWp3vL0Xj0sQWL4+tox/yg8DxMrKkA/BYVa3ROY6MM8zUyHg6+fR+6v5BP1NhNDu
AB2vJx2Rkd4/2zXbU9k8kJRM4RZ8VNAoXjV8fY/ovPvTl1RnxSvPdvg3tW9I/ZOGJcdclF+jV8KV
ElK2RDnrlKrMqrBrOpJnSjacWtaPdyd0SFq0zUxChoBe8V5pKdkkhkSkjb3t2KNsf5QOu5ITflnd
kXJrp6F8UjCsun8mXFs0fsNxRnDXlESE+V98WSXaXPIsdL2GnDO3AfIiwoOL5SPHsbwA7tR1yrDR
viiJzdphiQwuStdmFWDdHJiTROa+Qh4guEC9vOLNBOrTh4ETqExU6MHFKi0eJKKUSYtS8qwtOICR
o9FpN5bQ/Pez+mCp8Jve1nqryE58xKilrcytn4IeUqi9slIlEII0AJ3OZXIpLtFxmd8n/XRzWfQt
+0kYViaIJLQUnwk5FX2WxMyA8R6/sQ0VSdUDWzAk1zPcmLEc88tPr6iGpQeLEN0N7ZlHrivmfnJy
eGBkORyPOeYuB4ZxgFECrGxeDA7UR0L9yc5z3SekDikXzRN/JS/3wXbUiyIYnRWVH2sBM+Cbxxa+
GNtPjPrptOmy33+K+GoaKGl8LSTiDgoiLsC3XqZVWsZ/XBTeis0mK7OSj6jz+EBWye4Cv7oiWze6
20CkeQUDmvpuR0AXygqKXnL57yA/3f+BoX8O5dSCkC0ZeVuL9Fj3Y1aO12/5gETBsAJOLZnR/PGp
qLOtVW9cjdcMufyxBPA87XJmQHsCS0knfm739owtSigPm8mhJibEfUaCBhzfRUzNoRIWOGbknQdS
iitCU//vxuti4PyE+4ipO+u6XF3FIqkE0Sef3icy/hM1GflPmxf5URiwDv1WJLcMzEey3difrmR6
XyKBHyAN8Gho6RTz0L9Unv5gDOGiih7kvwW2qSAaEt2z1TAH4aWMJlRT+TgLduJKRH125L7zbzSR
2SxwwSdYhPEYeo3quLzrSBP8HwqEN0Cmms49Up3t9GbfEc1mLGPIGZNIBFRAKad4viSgDpPs6elh
GgNqex/f58khPw9ojRb6xrPWewpKk2k0LdwLAfm21arNQw4t1cTwCfR1AHc/79ohNiH+JdoUEAH9
2DllAtBvZ8gRYS8R4S/ct4NTBqh4DF4Ni08H8G6gsUF/MQC6fiMTrE0zoeOPqO1PkWTIQcbawc6q
oaj9erz0Y2uvDbirSWqY39cBu2uQrji6pBCeEtdy9lD7nqIQnaxzsP9c8NrgwRkWx2Qp9hkIxbRj
lcwFr+N150AtYfnpYl0ZVtTrL8lrb/s8M2avGdnnluOV5S0fYEG4McyIjSzvYAoOIKhJQ61jmgky
EbnSeO2zFouq3MHx73DC0dygvnYJdStTBUkdbCQVUvIlBgsg8eFqpM03L4XWPhY+1UGmqJN6ObI7
JnJME4Cdymop/bDj9ktJPyQeYSkRI7rmzWEUYnoQoddhHqHaLNyYX772xPg6Vtvs3w6aVfzJFQEA
7q/lnpWVOoe6ZJjyNe/bS5EMJ2tQOya8XFVaSBBUKZpiz2T3R21BqCmaUgpNFUfjUNqCTSs9xEJ6
+PI4gbPqQn/re/59KX6M3xqkX52PjcoPtkUGJ8S5WmZwcGGNxM/nXYvrw+DfETltgYEZnrWIJTlz
5HmN3hUqYqnP9sUrI2MqfIKrB1IT22YrSbEiE3Jn6sDr0VbVhdMM9PfOrfmIYJfBz035M2v961qe
GOEDisFhK2n5bJM4oqnsmG060GVHgqAYiwD3Uuvy8bC0zv7ikcas5Rv0m3BdbTRnYTLMC98kOmm0
wooDq0GO3cMh3/J3AECQDG4Pqh2ucGw7lJiAAdbaGS/JEmf8M5BS2g5y1ZTR+qbW+ajz8QZVOXxY
yrujYmun2EJhHYtnVkxfPHZBXd4ZqktHF6dznGbLRhoJS6yHZoicDuZSlf7FOnmn3Q/kkYXxxEHC
P7iDbVKDMvphdlBE4/ZafT2ygM8Bp+ACv9YuWz72yy/ePKsDmOKs3fhTC7PY2HD/SVngN54JyTjN
z+wsm2M8LAskx5m7YumlNdFiEScFYyda9FLv0UxYkzsPFyL1bTPWqZNvuvld5upFbluNm1g6ePOB
+1VrJQRk+nWKgNMchISNq1wEOjJ+7aiWbwpUZ7rZK7zAopd9eOeEmS8mJvuM15G6wPmqc0tcBCvU
enoItelssaj80VFwXZsRFbFld80w0O22kX7cAGdQRSR4fWdfJjCozOuxlNtmy5wkOhcMd9KTn3tk
EDvCw/95P59jNy2mKpNAAfMWLEdmnJA+ZqtVhFZVgMt9dWxUJD36NJCFGeBDO+LehtTVMGm2TiGm
2T7/tPIyiCBB3vNcuTuf1XAoCrTO6QJ3YtwAKyxLvUpAwHAVag8vqvbjQg7K9cwpTpiqNvpiTiny
izYj6+7AlY06NcvvwOyJCGEs6OeSiIUe3RZI9rUfsc2wzWYI8yx6TfaeLeA5+ulnufABBni29e6J
+XnoAtvAc6tt8eN1MIwoRwXNt559kvmOvlrQJGLP3JCagiDIYpLarP/zmCWp6xA2MWStyiZtaTt3
LRCfZhNk7h6BRCqUrqPuCIM5xRA8IzyTvuEUpYtpRtFsI6/+AjcyhWJhPdBL7Lk9Jyr0XN59Z1LZ
DlQWR3+q+SwyKo6yi6vQKKIUMJu9j9WoYJK4sa1OQo1v0xA6psJDH4djRtScNTTIcx787KvHuULc
r+siMFEXdK4lmFTc+nJ/1Rmcq7xWAuElQ7fBK/bqt3LmY5vE82V2NfLhyyekIFajcpE9DZI7M17H
+MOmVgsr0rgkK82fWPDAb1gHmcCCk1DN/qQVLIexHkOq31IkuKCWmim2E3DQvC4G8dpka544SqON
02YUHIzYk08SjW5ADXiZAM0cpVuC+UZZFs6iSks4xlTCSikUCFAcEwO/czomFGqKOZgoegIQ5Pzp
pXdgt2hRgIheQrNNDx5AdPjO1STxFYnVEAKeI1++vvr5hIFWDU2lZwZWfOeX4Lh0AD1W8VG15WJn
zHRJ+81NutSUkN0l5Eecm4t5EpHwuzZNtezRcr0TzPfimsvd8UmjIBSEz5zhUbV/rYlDlnECdi2C
oR377spnxvsvXCDtDQ9UaATRhlL5YwjSHmi2yzRGLIxsLx7+Jh7KroUuGpD0HHdFLZ9Yxx4a4Als
L6y0+fUvW2wAG/QcQ4dkuhBswPIaNk4rlqp8tkoVqsFuJumx7VAQRCKr7SMKBDgPwhxZY9I283QN
ENS/Gspo2r5bGWoVTa4ObVS6r3WydUoEsLWlTJ0/4QFYjFH/Zv3+9sN4H697pKVjOgwpB72nBiM5
Ymr3mbercXzCiqe3jasBD/A1SL42/jfpJ55WglYR7DvXS5HKAVkFejdGe3FMonmmReEeUCAUelNi
KWh+5f5aOmrMSVfvPtA9DYCLkNnXHpD9bE+M339vGUO44lZ/1IdnN3j1+Hpmbq9UxHI3uHnn0I3f
wcZvAfho4zeGKuUrHwRv8axsRhegIMebePQgB8g3fkosmHepLvIfzZISNCGPdWKxw980L3t14JZ/
4MBj0UWndxXf2zhx2iL164XTp7UCX+u342F8IvqUK5CETBr9miEXCwSCPRaw85yn6rJlXSzTFVEs
t7kKO1tp1pkGa9gG/YirMkSDXf8QqX/c8Nt7eEm+19f+M68WT4Po0VzIUtWEwFFmWXSon7+0C/gL
UKEgExe4rXp9LuOsV4RZZBnH28hLAeGRObrLhzpb2DtZD/J4YnGEgR7k2gFAvmBkSzjgUZNgsUdq
D8VTXrd3hKX7aEP/bxTTXjQ0l7hM3Q0e8yiEFf4Cdk5bJiJDQ7ifvj3onwEL9JOQgeFtV8avUz7j
GEN7q+l4nTROw4Xg1VyQkeN8M10131YUaC1sC0xXyuJH7rEUJdcoiJm93k0tL09ZHEMN9cZ3GvhB
0QoK/6a5840w+PnK+NxAd/5qvjnm9VEAm9DXuyQjv7Mdjklg+0qVnSPo0Yreg+Gr8o4Nv4Rskanc
YQZtJMrdxuGLe/bjiSOEDuKTCBfkPn4iMwaNMP6DY2MEyV6+mMkL0L6qiMuQLGYAIYVFDcfXREbZ
xFvIElgBY0MtfKZo/0+Dv7OXF//wLMXwrdF0VfJZClcUVOOSx/QNJQ1UXzExmGR+WGITb9LIU54Q
WPI/6t2L7yeYznCsFlQyoJL6ExKpTx5PcHInceHdVhd5DLlqoLwAM0S2KwPRw7VVAO5GP/Gnoh8j
AZxYHyy+hbDokGqwdtecuKJZWDJ5xWprz6SRVmywsji4STMQhp+tixTQSfhtj0lCaI2ylY0geHFK
OL1ZpjAIhVxKfZGrv88OWjZeyXAeXMl2wLOIusKFapYO1JYHf3Wb9A06rwYJku1wJSlIXQzUV1P8
NA1MZWa8qGMjN6hIyOCy9YnmrQOC1+0NA0lfdUwwo1vOLt3x9gLqiqaW4Yrx9sQvzz7GnNg88Gow
0VP+KkbK4BIG5p7wUqc6E6eQObqKncfW/hCGNR9CuEOUiLOpMn0JWs8vDzhbdJjOM7ovHO+Q0eag
eLfPN4hCGuFiX/ZUqbdw6OTG9jg887Jj6d6eG5n3utlNAsLIi9Qf91Yf8HcmHoEZJ8WaRKxs8QVA
M2k9JuMV+wMFF79S+u6XHB81rMPNh6avo4N1ZGTOj1f0KZ7M9D4yJ29gjtwxDRXr9dROmG1lqEMS
HvFWBUskaZbH6ctzFTaz72hXpXMin7rgbj8LEAb7tyhZmAKT5v2O870RJr3s+iDU9F/ZVwx1tLEH
xtLJsQYUhNfA6IL7IDSc8cGtLxbr3v0jPfGdprtaqdhfNRPZcR+FQIDT/jGYMxoEVq7A6tElB/NC
DE8TytHL7YV010otSqqJwvRwiY+KfB6qDuoE/VYGoTIBTQOdNY5aAcrtetJm9rl3Tsr79YVFdEtA
W+d2sjvJ48ibYUywC0modemu01e+KozinA8Vm+JV1Vo933kovNTo4l8s5aqCW1d7qWTIj0AJlNWe
uN+5DC5VyWpdLLu0fjA2y1Cb4W9WVf9baZ7eyZfI8zpcXzwlHI+P/Haa6s8PAHu/AqFxsoxm12tw
hr4WSqiUuS35z2eQFNR/w30VbYmmSaMI+/NJVgRLsrMciQKZz97xZYM8RLgq8sddtz70JQoblW3H
tdj/cMbzRu8X48JOlnXQ7kKcQVx05FUCe4LO1EKr6LB8k9pzogiY1VsxDPaiPNnenhWSfYdBM98c
ThYtCGDvJaGSe4RR/kblFaPDrwCZZ74fKhLd5k5AVUS3mFQGzsY7Mti9NFhrZmHYHwaS/lcuTH9s
TAluOSDgF2m2Ub/dQ9eeRfgerQnW3XMlnIrZHjfBeFo9uLa1CET9aTURJYba0OdQCUTOWmrlYqDP
Tp/gORbEWzwFu2GUkqZs+8bwXycjBrGz2qlIWzzWo5rWrL/DBaNQMX6A9W+tW00jwn7JOLb/b+JA
DTKC1uBXCWqxq9nYcxlM0sG66KP67DECpKq++slxOk/wzRdgpYp4H2QxItpOiOwUWPwIQX5FiwWV
r5Z3l8rsrnG9g7zs8jm6uaEqOfUGVyHOXFDxhL26ktDwFnkYODOB9SUrsnzrFFYxX55P1N28A2if
VaGCsprx1G4uuznyLfWMejrbwAedGd6Q9/AnwQVWpKc5UvELK4xHHwXK2rlYksckxpgr2TNEGKxJ
TenZapA72L+iIKa7MynkwXieXQVY8CsdTLStU6SC194jRm/x/OWMMESJIPu+oGm6GIsVvfMgqE2+
y0zpyfxqElZfAFoun5SjAbzo7U3Q/RDQdVpnHteQt4XwZ5awYLKdMpYc1ncJ6ASeHVyTIQ7cCgCN
PL/kYkpTTbxto6dN1/Y/wY3gpy7SkQh1xFQMN3A4dLYo/C34/KNCWWqGnoGox8t6dUABarwkPus0
u9lJceScMBMRmhy6+EagEHLHbCAqUI+ohidMG6+cFRu+5SDfrsNk4NkUzRW2ScVU/qWCFe5ozdr5
QbxF639VyKO2hbODC0+suq0TQz6k5XXYfaM1Yv1n/yBHHLKpIzGYfYVs+HTjhdk1w87EFUA0+Oop
LI6aX05LtT9HCHLEoBxDuCtZ8ncKR5FRR61wd7yhCcSp7Ijohj6GHrVLpIF8xe958BI9gOD4TFK/
0/eU16MCk3voJk/WI57url4ZcojriXCclTVfUGiiHQ/E7jZLg9vzk9aGQo+pwJkmbJzhbjrbZ/jK
3erY7yrpbD5kV9+9IKfYAwJH16SeMCiv97Fyi3MI51R5YTlv0S2+g1p6LlshTw6QHfWpCpSc7drx
ljlOFkAL7K+45k69akFOVEcDmXof+Cdd/DyzRU+69zZoVWk5k+pXZCihMwSKiCPpOQ+SIl8z0wfX
niKN1/7glKrcQAegksTClB6mgTE8xdxl2anAe9DzVMGWkpqUbrMlSm5ha9YF5Tlhj5t2YnJIxt+d
9/RI12NHH1atV57lo/jj2BY30D+1xZVxpNDEmGXoiQNdlSz+ULdeHHbYT7fnvyBvd1/UPw4TzlPp
DUrs+gLMA2NPiwVux5CM6eSXo9NJMbIRiOsNEa4mCE/HWAdhVdG7D4IBPVs31YYRtX9VmYquaJ6A
cE6jEeF6/NDhkH1tZgK6wzIN7TL/2EJoUhJsY4GkUXkJyvqyQQP8XwhO45CsuA4K6C+3LJ0jkend
QYxx9jmfvTTOSFNckeMiXPX0qqgkg7WRJnHfPxnEr7a7MXoNBGBXSXFKYDHtwmZy2Z8qxinYKlOC
mRRDTMabaaPVJmLt9Fqz2M624kfi9YRRVeY7y1SHtCKVq434gpzGcz/CdzFOICNxGjBIIZGiDI94
6sA6AML35dTh74sXd4chHTTV14a9itsGYXMcqLsCguWfMSRYAd4UPwtAA2ejOcYay+w+DDAz1QG1
ZaHcCr4WPx6rStgXWpF7Sxp5Jsd5v5PMo08EWI5g+flWBoNfA8sMpiHMdpsoJGt/VE+Juc9dgg8/
x99jvnuZ2w5ybl4QccWptxrdpK8ewzg40SGVxGybiCdTRgvSO/TvGEbyIovDy8I+REI3PBEvr9bm
1YPLpwb87ceoAs0UhHmrp1HY7HWQN/m97QPF/RcuQPevBibYSLw5vpWGleZ0ZJl0BcMnDyuLRpj7
thbh0tZ+/onGtZHAETZJjaYTgVWVoRWh4OrjYKcgYieBeydjPEkkqplo/x0ydn2mtexIevzgEFax
0FlssJ3VJxPXe4iz2DS3hYjflZEJA4Bn2EzdrmC1/O8F0wG+9c++qZbFRyrAsb0UoQkkHvoRNACo
VhDauAItUHY8xiC1uwAyoxtvb83CfJzNYTqrGlkdtZYkmTd2Xd1+WFraF13x5SVy+sCQLDNaUet8
uLYeAutA5mG7qe/fqlykSuZ9YNcjWBrSXWBuayQCk7frUfajT5OgVuFIKvotOOzTM08HT21ZlNPP
fbqFXy4v7dYUdrPklUNcdyHJ3T2varN+vjp/AN5uwR+3ZUNenjxZ+3cP7/8CuhkwLd2BPxK8ip8t
yikSgYKYEkxs4xnRMi6Fhm8KirBaPRndEsfzBRtkawsnwV6K9CVv5tJkr27Fd9gM+sD+cqhN68CZ
XAgbtuhZT6gqRkhfn8+D6/KX+hKKlDqpo/Mnv3HohMEITZzSE9T0K03z9N6XIXXFAHERvzc/WNs4
ieaM8lEuVIsIW5ikkWz7BbQD5rN5t/fMblmG+6sNtYCB0i2qoU9rkdCxY5+WwmPwo+rM2WTqsAov
WakADyKrDwa3YRtz4+QA6kICyJpMY/jlYzChDt5Ynkp5m+yQKXpCSDLUmCsRJ8MBF+IFftn8oKeU
iEmCGUmLTAW6YcOorIm0A55HlC/dZWjPS4iT7PeiYDvMITRn2onXmWRFxhNEoIn/JVoZCXqzORRr
73m+4dHQux9JOedCc1GsmYLiRYdjzdq3HWM7irs2QNIir+UawijpqkUmGIQUigNze101uG/UTb7T
W0Gi62YQPWaJ8CWZfbQrDlKH1D+Gg+dh7SZV0EqUxYHWo4rPG7wriZmURt+Hd4Yr+mTLA/ZXPkK8
SjalaQ7zEklxlffm7IPrHLTiwxIlJ58n3a9lSRbJUmxd1S9o9GP4rCJixk6L+FfzWeMOc6jymytm
jCa639oD4VPoKRr697OPrTsmxeHMwPDryBPUGS5NlbarjwffPWon9hSYR9gyZBB10/4WeGxtsr+N
eD9mMUwo7/YlOX08k3do6TVA8Tf1PSkijekVc9mUYqkcTizhoTqgjp73dWaqNYlxL4fpAJ+JqAci
46/MZfpntaV2OHBCpkrhhdR6hscwW3HecXv6lL0bJ+7AP22rvhDsAHvkQPZkNhWw2m84cvItOrFY
Y+4IJj6PWVSPmhYDQcyViKhUzmlvIfB2io9uweQbolQV9zMOksor7emlXnA3ebYXRv+j1+4uxvpv
CIHpQD2TH9QNhj7gPLnPicTGjQ67Xm5rxf7l+AvLRqQGIKMguJupQNEjPjsjMqXAjcUj8hiwO3WO
VulQjsxD00OmKkof5PKJxDfIUP25LOd958MDkOv2lI8alLF5oPHQLlNx8l5S1nLfC7p+0oVqwnPi
9zxd3jsg1eAGwEKD8zB0TY6mBcxMcdjqe6J4SGN891rY4mKwPZVKW0JEI1boENY9+RU8NrrMZR7m
A7njgKfNtilujf6ZbVhmSzNEGODwx32n0vl53jdiKrH8wHd62FaxVHbm5Nt+obNexw7U8xjS0OWh
aQDmrqYRakhMLdSq4PZmc6iH8IB3kYhVlXMkWEo0wwPoGkBBKHFtsFY1mkqGg7ZccPs76QQ12bdx
2MSBUunCd+yhscrOtgHtMHHkGHp1U70bwdOGx0tzuyc3ca9+/2VwOSOcMj4HnUTF9aIiX5ONyEG4
Q6FqoW5zwu+ZlR9uFMBymauo1dAVrMrtLfHLdJBOJVduSsPxYCIsv0P7Bjp3HoLTEuFR+yzqz1nx
ejnyZQk/ariWasOIAPO/prcBB/taCwHwrntel9q/2JLbWCx/XF03v0MSFaFs14DUIanPh8zW1A/N
DWOO68ZZaw48hJsFGCFSfiYv8iiyhOLIhpU2IwgHPnBLsaa0DMCi4roKsDY3BTLfVszeV6s+28ds
J7+2e8s7ayUKL54uzT4E9UKpwOSlaOJ/XunOeRQmMX5HOM9U3ehylYSkPNnEE4zRvrHaUkNw0z6L
WQ0MpdzVpgR4YJpk9MvjsfmFo86YXfvP1AlcEWEgbGl9Tlbi7moGaRXRPHlrK9nXsNFXcHtWdSfA
x4TJDK+0RytKP98CtUL8xDV9ccOFxZb9QPNb2ultK8TTfQ2txhiSuBmlgesp+sYxWIfbqo7BKsUG
ufZZ4gk58+ihSmDGiguGc7AOWHG/PkE7F7r8ZaBf9/5aqJ2qzNTsmA8xvl+t8RRafTD0yxZ7Dt1V
SEH9yrdi9cdTWGhXMkxJz+1W7pkYPtO4dNufb1CEIsrbuyP8K2Yc5TIpUaF9lH+tEYyrmxXPd9cR
6oi38bKi3C6JRwQvRNgve2GnLjACp19L11sXXwqON4sT/MD0Uzc7Wj2MYGuV0RcsZ6P3sAuSsN12
3R8iqNZWXZZRGcvchkjMkQ3kbsZxqtdHdRH7Wwz5BO9ywUwF5cTH4FUqJYzp6tY3kfmiUSiULlAp
1mIqYWMj+1Wkq4dZvt5444a6UJQJ/EJXpem7qMQ6hSUxOK+VD0XHpF2m/wsE666sayb9OAz7JVJ6
DvFFiHiFGeLsbq9AOkguU4F0qPIr8dXrrD7i4EDuVpVAgzrUfpn87xI8vClaEYCT1Q+DQfsVlNUM
v98YYA/0hBbcvIfiFwkkHgN2SNMdPw1Qb0A1u2BWkpKvfDQuzQCCOL8+IWHA5cdLEUSPX0PCZqgC
TzK4DYRtk5HbS0nUjwiWg+3A8uVEKA/wiXw7UUevcn1/grOedlSEfhIY06oZXkDrJLpVPVSkGvVX
IDzA+Rdk3Z0At0PYRP+XT1uxJo7uNOwETiLAQPybeIpt777EOC0j6ZfNyK5FRFyv8ekJkD5ZEVpe
2Nt8nc2qAm6skeZZkN4KopR/iFnC9atekeV2bSla2Qmiv+I9QIieCaNm2prsuLAphC29+UArih6z
5YfnotRWlbZaDXRuG48K8/iQhqzLVuOArXDATmGYRX665X4K0Cl8IQXG3oyiwnErAgkVjEhO+3tB
YdqSZ3nwqMaiIGp+lBhsorwtpU+sAkvsrPOVQ7pqM3K36bWcjzU7V3ONp6baY65XIcwrrbV5FFor
m4B3xVGCkQqreJW9O3OcI3J432EUg07J2ciRonl8A/aYar3HSreI8znSczHbXDfCe/fpyJxG2K/5
PAs0+AtUvPEjP3aTe8JGOP8nbC87qOjTrndBSp0OjjFDbYX2u1pSJ5cHgA2w7ohEmRM/B75ml4Yy
RSRUJfUTjiWKdpXLhNy8pmNpwjxlEKZvQR/pwJDkfP6wOKElbBEImnQVLTCTvRPqUkYKcNgbptbj
c71BndN2+s2DHBII/552hrB5I39mFLXLy4ZknysEqmrQQDDzNmfiGoGw1EPryfkYUGQEU3gx31ox
eGdN3ZMVphxYn0kbwjiqFZTecow9+8Ahs16HFiZO95Lur0tRBNnpvqgo3kab5DbCSPKBXYAtUMYJ
WhKMw6GDIUmJOEeN4sJHDUGSgL711pgRqa8fPYXc+RPkSAKutHZt1AM3bUckq8s6LeBhsEJpp54N
/7o2R2zByAQhyXN8REmCYmU6plsx445wVzXZKuVdM9J7/x+058e5AnrBDeZ2unN/wj/txpNoxXVc
Tg0AOcTY31Cl2Zio96R0uyh85wthBy/EMth37s5Jo464CUf8q0Dr2JZ+UH5OMQzPPFeKC4XBFDBv
UZv/dzQB9b/lgsUR2PvftyHNoR76WQjXomxQIB1usi14C2v+moJ1ZW3+zjmkzav89C9eZRJ78OX0
QZdF7TM5enL5Ur2TeBUtPUJAmoU3Gj7pfxJUwSlTLrh685hFOnrEn+1gbIqB10NDX3DabUqEOyxy
yYfWSmlngNK/PKU432NI/SqICZyQouB67piyE04WxD0uSVoh9uDKizPxWfS+KBDHbh/gRwNyLbRj
8LoGBxdnUa4qXod9fwcFBOJxZe58KvUvgZllNwdX7H/xQazEVxq4/TP2y0eXwE7laOgiYU6/V7ox
T3ot2qFdDBWvDEyiQ1e/9yAhxsm5xErJz2FoeBZVGs8RpNd5sq2mBvKX7fYGzLMeQnV1YgoGBEPx
oYAMPCopmrhHAfc4sKoLxDi1cVRc+HSBbCTpgy93q/oLTsYXzVSae938b1Jy1xD5Xe+WO4RKxH56
h4hMAhjL+RstoDt8XZhHJLqv5CExxRTq5HmnrRpTu8cH73CGGUwyUZZHGludbAY+In0z2Fi53iiO
fqIJ+3n/4mqogqxmmrKDuOmZYbdCmwPccQhkUon4lfJ6xry0mmGNZWLp6iFro45fZp6tqxMMmJl3
6DMTI5wvPurNUYsSJmVIyvGz2EHwEcUGKeQwgKvUk9Yn1Zwf4/LQ0FlPgNmxG+1aQdjt87ZurO6l
GEkoJYlQWdBJqm9SyfKjkATfl0Mm1aN91ICvUT0Bpqm8toRNxwgqf5uNbWXb702ll7nlWW90+wDU
TonD5+Zjj9eMPXNj0dEA7cW8lOVOqZQSs/4MFEobNtX/kEB1vCNMzvi1pu+ZL76CPb5yFi3Cugsq
QQtHK3ozasIdLF6HFGRwE+eAz2pFMHd3tyhnwdiQVSp8DF4rrPKcxNSSLKWyu+9yT2kCRRLGYluu
PUOolUHcyyMdky1+AHEA5RpDHTyqcaD3rQ+jqoYSfrlN5dgtJuxqZYEdO0fpbs6qMWumK0ZUP6/G
lPLDKDQ/YkgcpWqWYBiM2hl9vegaw/T34FwzKXPrTZyZpNFpRizNhwCTla0ttEGg2xkjdpzdTgLl
nhx7prmuirJoIbUCDMDQx87PDx99VOe6DOHCTO//WdE7mY9Aso6zMPAgNQg+ui05XlFIAEdrpyuk
RfZmNP/e0odeFEkZcgIDe0GPs1No98gK8p9Oxiu/SXGmSAhEYna4f87QpNwQhD7euRifbf8C9nlM
3rpiW40nJv26L4ywgxEWBq3AtXRm897gE0Wd1Kd8VsaeXoc3ZTQNkz+8LPIZv+NV2ZhhGl7NOCVw
7Qu6yGJ2xn/2JFMZfGIxAcCHn3HOU0uNZgD2yQwxLARgCuujKW3vd8CMPziXMleo2uZqvl9fZapj
K+f17fykV4y0ejfrvxwcmsb4lkH027ls5+ScRAia2fWHMM52t6XJLTTo+mNktPZ1rTfRsfX4XfFJ
VibNQLmMbh2e78NZ6gW2dGEF0Yst9P7kzZFHeBfhH6+0gSFQbO67HsB0cPC+UjUDBgrJ5O56PENL
5QnYFyZ289iLPspq+9ktNFVT/aoyxiy6VVN8Fwz7/JWdecDJ17LK/xj6k/+r8YaAJflmphRWOAbh
9HRkCiL6PrZuzAY+qe6J7dNYL5epbAjwIIB0MSESIZSA3HDEtapZBXUnXWTzmXCH9hfych/nbpkb
Os1PESB8zTcW9ys9ldoaceVRRoGT1ih9T9YwYY+IFmzfX/KRCkman0Q5uTRqZuEn7MZPZyJl6HnO
kn8Odg5mBaul2LsJl+i9VuVEBeqqx7Z9nQDxURDmlmM0V3Qrig04UIoRtNlcAA29TFMjcz8zPFxY
Regz9gnUN2wIooho54Yw1PegU2WpWCGW4j0K9jmjDCZqc/0R/hpfVvYItaAPEGMDosUsSEwKgaZb
BE53rUKqd5wMIDwcgF8VEma6mdyWOBeYhcHM45XEgJdKDmZJXMTTsWcEMm+g78bwD96WWA6rLcNF
2jy2xp9CB2NmLgTRoNMrv0Bet0eOQYxDGLPZlnpfgmbp4+EjLpREerVmzX4FJifx9hanTGLZuErG
63QWRZltoKMEduvJaYXBuMm62OOf2DcLy6RHIOLQyfrv/2SMAku7MGDLbmOBzO9cZVW93h0G03oO
lIhtb5uK3W8BbD77jJL+e5yK1lvj8tkDET6cbQnuvNQVmBclv+u5IOOhhEu4I3ZHnVnztES/UsBe
PtIBUP3VYhqfS1UreAMUeWQUg6DHWB1RKHdLnhz065dBPRTENIPoDrzzrcVlvFYiR3wd2yG5nWzf
/4dhdO26kzkvF+IiwR1pmMIOL81xV0PVOP6kHtCw6rH++pdbT4kbCjsM3tCQciKlriNUC787BQAN
jJkjGUgee49FJKZSuV5+UhrlKrchBepXm7M26VkCXMyDTk+Qzoejdw4/aD7A6k43p3gcjqRq8H6h
5t7ajlrTn2qen7jS5uDAWgkxjqaVjcozebman5f6SKx7DcDrxcs0vMxaeEGRD1F+CqiI+PsRrwxI
FC3mikW9jot2koQ8c8k/ANr9YtOF3leedngdO8XgwRo+v4kdUFhsV+h8ngp+i+KLdrT+fxDt12Zb
e7q670YepFuasjm0rmiZZLL7gMKVk19KxrYyELgP6j99wacEQzsMFF/pcBhF+db/j1AhiTqiX5TQ
4VM4w7AdjapFxnnH0eL3z7N0HSFr4t8hBegyKyIr/Jg2fF+6FyOzdxJSgdEUPDHWYFXWp7eSWi8/
YAMWsW4p125EfHtdkH3/qRhmk/RClMfa16ByWv76TemNJ1Mlx6d80tuTvRce/kegfaueT4WbdjDv
xybC28S7xrobYMl7HzaNyX8LCRtBoTEmEFjAkIt+CMAxNk7YWUiwvmsgQSl5COx9RebUYk/+FYQb
Yb56O2xsZKT8Q0FPu3ROfHZ+hrC7zXjnPbF/B97YUX4gjAjeAI/N8plcUSlm8jyd1sSlRbnvgW2k
wZ70UcFaAKe9EB22Xu5lVr6AfHBTlR8Mg9kO4qmOB9+U1l8Kbrne+PAAaDbea7QLVlR/LvjDG41F
nO03neyfW7j3C82DSqMSwNozCZTTp+Wz7gTNc9qGMX+fa0bsUD9+IgA2S4tSIW+p1U2nFncvwHuM
jUr7eonUsz5pBJI4adJHT5x92UhZcmqzhEEUci6saXHbibJy3v3yIKB0vV3U6bI9MHoFMMx9/3V1
qMMiNGpnZi+4OT5avzf+xx2fQWKoCFgO4fT9Kj+DFu/FydBEPclSqCbj6e27AkTSlD/9FHuZXpal
/utSTAVe2ewj+vQn09P1qFkuJYJrf5Y0zFq6xOcjMElfFrI4tDGWc+nN3gslzCUn9MA5Cv1zyZXC
FQOaTq14wToqtYyuIjO93WqTL5roVh8qCGPVhT+rpQuV5aL68Ec+ffs9ZSWMCf8/YqSCjHbf0/Lf
boKFNztNm/IJRUZK2y75oxDA1NbmsEqOd1/6fylegSAUNHfqdFPEVTAIoy80hECBfC5L7idZy8fx
neMan/IwlsnvfEO2aaQjoaVWUFG4QizNZirxquUkbG0cVyJ48PiRbX1BEOJPckUetcrjDRYIke2R
7Rgy+WsxLSy4xrXe0xYqK7Th3enq/dKnnuOHis9zj8fGQ7cmeM1vkykg6sLlvk0bt+HCFVT5R6Vj
52FzEaatQ7J6YENtByK175E0asf4XCYXSb0yUTtqTrSB5pmoQbgiGSdQD1vve1Y4XfnGvz+1iz2F
sX6p9QdKIBzb4V0AAL9VJS1W58zs1UUPAPTDG8iMdqMVCHYO7XJdjSw4dDW/vgdunVaNGK5VpFoA
zZE/muXut6w856iI9SejjwphpyssqhFoDuHdFdjJBbykhFGlMiXXiLnNAsLB5Bj43d2SvGjO3EsD
pI11ka8SJYEgN7WYLCqyKImvqW8DZy4cOPGk1cvxZK95VEg5jYjh5IGTCMOPRG+brT99Su8q17bi
ff1WPTu5qCZYtuREqJrwNnt/QjRrzFhjw6u033IWS4op3ydGm0Xe98rDgBV+K14ATubNEcdSWIMu
nLrB+BjJ9rqntVAs89p8JYK3/JVGNQrNnL5L3luBtvS8Mefiw1DT7kMa3FIa1rZySWO64nC+G/vw
qFAZWyKa/p/19dlhdUwJOEoSSrsZLNRTyjso7C+Q92W8Uwu/mnrxxNpL7+arLwZ2DoGQaN68wtIk
Yx+/DD0OSaXeGZkhcvxLZ7f7Um15gzLlNtyw0XKtWnkldazWynTwvms4Bb1mK/csGXaBT11XGDBK
HoNifVaFjLhCoEmFWOytCfbb1i9qbpDpliNtim4HscvIz47ubGnx8tUgDLUyGQ/XFgEp3b9GUMUW
oc2+PWwDvyOtOz2AEJ2uzKc5hCaT3ahyhAMtJCShtmAtUhGc4UwM9/yTsMSNssErRM9vh6+HfLGj
5vs7NATLZq7S6dmQBEShX2BykD1H4sEZQos+NTKHnnwoW90zch85YKfFII7mvPuGHNf6PsYAh9bY
gdU00jm/XwzryD4EoC5iJHCoY4MAXxKw4227T3Rzm2HxLuzgMGqUIbqnpUfaCIsZcitkgpKWrhqc
BR6rreZXiqKXIRKfmNS+iQcfLiP/Pi3PKPDUGPjxcFeMm/9qRHimozz7UoNLKuLpNav19tDq0KDz
ZR2WK6cisQ7XeJfH+4/ptL1k9Xv8x3SLwcrGhE0d5yC2P5qRaMO1JTExGj0Tb9dHeaGEUx8Z5QKS
UA3JGfAYKr98kZjuaF7BN2f+aJWXouHzT2DK0wYF7H19tX8YIV3jw9xACZf0V4Q0SRHDK9MilDSw
pkCtL0VPL19ypN+GJuKOwWm9N8StGF9H1bby3qKOLa218yadjb7k0J/W0JWNEAfBwcA9q+Y7XDpE
kZKzailwdxJ7iJGDuDZasNxAdaY8RXZjbv7mMvwxmuCWdgBzx4yPOr6B3xcq2UbXS+8v0MkkJMMR
l+LKNq3bLfxxraKshiGLjKZfagIGRwBhSKoydYcW3pKfMqNJ/u6N7cYZ/8AVxAVBYK2IqMv00RcT
4pjYFvA1tc3l323fyOf7PixBQTSjjq953Vs04cn+E3d33F7lU35qUR7C20/IUcQQvwU5AzeMbPME
Q6MmGN4YzfQ13jaVzAzavtNaA1if5zflTgeUzP3V/ZAm5xHDwL8ubjtMkoYIoKYXWXwyn8chKkjm
5frhvJ5/wM4jQ+EI4/nizOvpXGEUnE2vMUBX2GIyVzmvsGnboVuHGNNK9eFmmUbrc42Tu+c+eyLp
kZuK3FKAw3AYj6ThShy7PBijABwsscglNqhMeh5Ry6WSX/S4tETb9SE1FfBG6cqKjMHhURb/mcC0
uSNgofjq8zcdC6832JyLntgdJq9lFydTHR7it23mWatMD9nwo7uFqKIzRsoXO6ZQa7oym+PbnGry
2teIvKB/A5HgohsMaRnSQx66/hYOncUmGroYPownr3smDsVl3AdyLC/+wQ5zcbLu9lGPkJ1+2+/X
zLMUJuqegnknG2Ox/ipmzY+nXXwIjIlLq5T3h/83eShJ1Rk8CPs4uzDS4iDbn3vtx2tZpT081uBy
17fBle4dOgAG48M//7YICmiMo2yDsuNV4ZX4p+GPkQUcJbx3cWHtwIVQOMOdSbguWm2RRmjAkIua
q00B9HZYMn3RcAIEAj07eRQE/5anSk0c2zvA1s8oilEsz6hIEem/7L2EBqJb840xA+fRY+lNWiPz
0mtaVo+3iGlzFGW5TDWf/fFmJH8ZbxPUwbPe+TImXG0AhKvWryZITe8Y7e3z6g7nsIQ2wOuchWii
Rpl+l9k5J3MDeYqCrbKUrctT6RHjDJD7d6PIw1UqQNvQjkrOO3IS0E7gkxt5PpUwzCdCA1IjquNb
I+W8PgsO4N/QNj1yK6URL3jdnzhivIRY0T9DYnUNUqUjVl+RSK4g/e9e44NkEKs1AIAUbPJyft8k
hS4kqUCol+1BB5wQEQRLteoOsB0mOjinvpU83X1aeWKirSrEYLvZI82t2R1Ow1O5Wzwu8lFPdFY4
4wTsSH8zrTfnKBux+IIHW3WZBBgyuoMtLB6Hb4EPotzpOQBbFebBinnzZHwRsE2tjd69MsvfKJg9
EHGRxkD+iJ7lBA6H5zzEpIArE3PMVzRgY7mWIAZULs6JuEeJ8bntUg07qsaje+8yeaR5bctKxGlP
y0T7mnOoy3ioKj+b3Gg4+qz32kRKyNar7gO+WVMULlLEAwBP+wthsSKJ3+9mi8hd5O7gafwo3L3x
BgFN1wOSxC7VHKlqQqUBTYmCR2r0ll6p53sx8dUR29PAx2vnn+cTn87XNXMNVTm9O1bYUww0scq+
qV3wRSXRUg9ADd/E9wcrh5iRn+IeVvMNQvxJq3YQ/aWsY0z7kTp+TT2AwQ3Bh8OeATa/zUexpaYJ
RkllV6rwLX9vTuBe415CYM/MhJQ6PXzgcH/GtsXN0jyhfk40pUIn/o67K81wB9AEAm0MiQBymCJ/
rmH2Q05n1JxTk2ploT4Bzw+b4Xp3uVwoMtaXICx94vzFZgiqdvnXKnj/ZzLhCpxr0IsyeW5dnt3y
rJmRkZdcaE1bv7zbuDB9BhgQyNpeRs1vmh4msGwJvm7wa1Pqaf6mqO6LpOuz1aiVjN81BJ3B0Urm
Nq4fl67WA7JqBRF2n883M7tDXlLENo/wNT6BByhTwmlFOsxZVn+mIGC7U/y6bq8hSmUT0te16y0s
LMsz6Tx72LdXXThhCtsl/32ZMkEhQs0ENReRUSyEI2Z6wluPAKk4jG3ZznmqgreYFixeOy8/U6Gk
11NpHveC/U2hgehN4aDrdYRByR7QPsKX6nc30SvyfBk8egfARigesEWZ2nNfsKgBCWZ1uWYrZ8gu
XrZoF2E6rQOg5n/fjRPocFPoKFaXHqsw5D51G187CJKKbpQoGoM6U8M3kfrGelnz/VAT/ZXfh3fM
T040iAqL7BQlxQFHGJCRlXElB5Szk9zqansWJhG264/NNEdysBIbpN1lgJ6Q5Nk1uk7sMI2IZW2s
f/lgzZGTla1hvZ96v87gQapDK8d/rtH3hZD7iMJMWmEhF2KcVkMjnuATmZ+qY0s5xGNOz66+nDNB
2+UAVc5ndxcZBuJqtpojJ3ggrlvBVaiHtA8ynsS2z+Frt4AU5rFPS3fEGW6oQf1LizaMKXQ/7ynY
dY5nzQVrpc3VZ8XT93+dmDU9ZZP0EUzo9TiOKNaIGfsgNoqBXE+XN1jaM9cFpodZ41IJxbJK+9wg
yEMYvdvT0SOtcKGrpbSsz+7BObn9IUsO0UWkqXbRK2AuNMeyCHxMXdpKfww4W3qBy+YKxM8tS0fq
2PhNKa2OcCeX0sSV+XDw6HcjPdhbvELgPqtMDs8rN9mS0Fdre12og7kzk9MlOQ7h0nHoaaamR7CW
I678XmnvR+gRYEcaNX3zXqFSC5QrZsEMoMGI7vyUeROqlo9ht84wl3o0+JJICgr/CGMSHOaAW1ZT
LlqZndgY+APyuS+TYm0mnkIIByDyaIpGAzGeXAbePj9djtZvotqDXDRaWAwDRyIfba4LuRmHwE0w
FxfAB/sP2RChgQtCMdhnH8gAUt7z6ZP1nyZzYXvRAcF8CWXIi2fGOTpRzmgrsoCYMx13/NDh/Kcm
+yslfjG3gRxNTwXi3OO6PhC1xroFLIzPOHMvDr0Wi4AT3Js9TAsMyI+OdVA03/WcIY8xyfbZIyFa
k1tmJaYo8XFhe1CI+i8v1kxXRaBinW0rz/KJJndEcBV1aRdNvZFtdXRSbejoqB/dLnEBs5ZdLhdA
7aB2UAJ4ZO/7sTx1k6q6uRBRjydtcLA+b96QuD78VmA+pa7nM7LovmHTXvl2gamTwlB5nVJjxm9l
nRcq6GszxnRTfnwgMSpVfof3YmWtD1nI6cuxw7TqMYMk4Sf2Q86PBYpt1lso6Mz090fzxFJNft0h
f5BGk060LhQraUYQI8fJjV3tcCzjUfqDnz4yKFTp012fqp3EfDbQ5WLwbVd8dm/Kn7/OYWCG2np3
Q8hbbF4Hib4Pryv/YkR5z8f2NPJgec/IjXguaSX4xjAZKQTH4eZagbMF+96dvAy0YWl8PWrKbzbH
UST35684gVRYsmWzJ3FXMssAZqhGyPXaeI26RcMq97UFOtTmp6T6tYlG7udNF9MxQPwhTkc7Z27a
dcbaEj7s1SK+pafaFyNqrGDUj4vs8X9rzPM/vAYVYuGyqesbu23HoQB78KNJJTl5XXDJA1LpexGT
7DfzmqSaoyUiCfKxZR870iyXWpbH4usG46zCIcYRkxaBqdZtdsM/LD0+WB3ajNL1d54E20PNgYoP
YmEZe6Yk66eQaVgi2Tms8DqPMQoxYnZTdEOl4rKLL/nm8b0JMCIJ9mNPWv0XUzZt111ceushmpjh
YcaDOj9mO8ZcSKDoK/49x3Biv0SxDEP0NGgOckMiFqIOhsWrYWU+GlcxDkUTi8UmpMrqFC4U5nBv
oa4xXzK6IAqIG76fXu7up/JwfE0p01KkPrLr/vlRZuvM7FEkgp6bt++NzDmB4CNY/vUSNeCY9snx
LczskOwh1qNGWiPjZbXbhCKOt/z5HFzeaE0Ieo28+Q5eVQnNR6jsERqe26DvLqGlLiBIQotSys03
+fl6Xe0ExtgOfH2SDWGqhMPP/18i9UVHJMrF9u1UTVEtH+LxOQEkY2bAgvbjXuZoh22PuriZ6aV/
l4Jjf6xmR05tX88MvZJ5su6+uAAEIu/DasFrFsmeOJ78E+57P6TB/3N+X4gc/OXbqC21RN7CfmER
B97VaKGyMxCQFP2Eg5pYtKjjZnPRQAcRf5Bj3THZh5K2fbUvkrnSr+SlpTEO+FaNlpXvI5Qc4CnU
EEtE0pdSMIwhKCLEzZztlsjNtgo9kfe7Nqbff6dsSQYazPG2KSWrFYOzeEGprX+ZZQ0YQcF1KNvw
Q8m6rbdqPRbrtrQP63V+KrnAtdU+edWyOYbBGuggfLBwbN6dsaAV56/NOIbDWEpN+6SaMmf9m9HE
GSwg5/J9r9zIUy4UbvRy8Q9uJe4Dak8VeKx7ae6sDApz5pgSon/edvfP3xvATH2BUlk7nN/odhiq
U7FIo0AiRhFku5l3KMMbqCUxVRIyra2/EyaMrl/cyf7uWj5JQBmX5D03sHKMZ1yi0vSBXx1j1iA7
umtZxnhhx71omLbUivhioJvkQ7k+JRAf6ytbgkgS2r5bDLiq02JyFVVLtzUey2OrO7X/tbeqUVwp
Yv3ZQEO/FtzQjqJfC9mPy05MPdaLrKIdBpDx9B+Ru5UTUaVnNQw641WrmXYUCEtOdfTNCid7Is+U
zW8zCJV2SVVOwF0Zr6c5moyPW8SmGIMNQD0Yd3jOoyWR7cyw16y9o2SITa6Er9bGzPwMZw/AVyf/
zWpTMiTkxHkgKZP2LScvjkqELkQfPqrBGYXgD8/B1Y2JvPfRdT+wBNsUxVaXid9njGv8yCnmReds
rPKCOwtRMMG67fbNZvT4Bz18w+NTu5NugSRu5ZPpR5feQR1IJeAB0XNwQ6MUrboQaGy4IsSSYMPc
jsali0so9l5Xvbm2UPkadoJrtxHyYfG+7mffR8cqvrJ68dV+WYLMjULtAFiqfZvRYHiyhN4jlS0d
lzbK1W5wHfQC3PkPa4I9egHyb/cxkA1ld+chCB4UQOn/7pRo6E6AVw6BJroFCcHA9jjjudTeFUZO
rQ1iDI6hjC7almwK2GQfbDheQVHzqOd1BqzsNu6xHxfqZbXfzImhrxAj3SC3Q5AP6Mkq05HJk46t
gpvd0YMvlvYZPT6toNZ9Y/+cxxPyF4RUBIyDWtKwNt9EKoQBW9npWX1vdDFCJOQ3iaXj8q4fdGEK
VGcDOINfWM7X5Ga2O7IkPX6YyHa68FBrKTBxhDGf7Hz33P3uRtn6MOHtMH9LyNK1/qmB7TwgDQux
P1WT1HiYMQ+jD14KE55ic53IjjjYgrxLpy9/QWZpiWpxpsjNeRcpfa9LGprhI5DCAmgKZPuuciR0
h0KRMkDsxfn8P0nNoKRXecKuhKuk7n6WhlDO/yqlko5n5s2cBXYY/Hib/bBSWlwdCcljs/UzGEPC
aRs4ZGKk7t/ulDa800jqZFgiTLqhx5OwEcuRHkay4zYJQXHU4icA0ufyfSmaiLLdWfsr4IwjYSfy
px5O+OmWb4umiw2UhZz/iRPV7z/fzWxUeaRxgJs84UF4x7d1q1h48G/YkwkZdAEzoy7WUamk0sDN
PgC2Lk18rLlKzw9DB6TlmhMRgIaElimEP77CHZjEA63iCE3++JK0Y7IMlBTqGCXGsovzr/yk53ze
lKZTLddomjQRlF546puReZFYl9SeyE/42NWuB3GWzNBxm7LmGDa19ASDAVzGedUgdoBKHeZ9pFh0
O9siHo3qkYm5fj0oo/11CvmNTbgzw8oeSX3TtdZljsj6NOVGU+do1lm6yxjCWmcAFlfd2uNa3KyU
g2VyzyzbACbCm/NhkJ55+RgMSLVZVAILb9HkDWNZPvoeh5JoOl/7DuZBm+Mz8XVBRLY6JmHmoF98
8uQ0T1a6cpIBvlN9EMpOZ4B7uifKHNZZZ+PeIiIKRH3fcGrC4agZta1n9OE/b9mGtN44h0NHRGpK
JexF45ZwwhUPLO4wDVouOxE+P4NG8vZH1Ci/kvvZS/Xs4Un45kxLm1GQ7qx+NLoI3OSvUyZgD0a4
41nxukhz7VYD7DwDMR8KkPlvuQRznzHNXi/M3N8o8DiZEJkgnBm5thg5HLKm1JyQ0+bLZ1+R1i4T
hGjijDjq4Tca/k93n3HE1LiJ/sDeMOfaPmquJWJ1qnaHQ7vxi1+SPJNhGAhrzzpK+heSunLSINfP
9iv2VHNKqjjuT9O2VZRNwoF2D8BqeZGfLENSHcJ6FtA+O6Y7MGGcTnXBsgAbExfsy171nPSWWhvK
4L2+gahHeys+2P+w+pGgI6oa27+nw4sXw8MN0u/q0Ld5mmqkW6e79i4rdJJ5pIfPuMUKKIaItNk8
qk/MB620z1GXOMfG+A+C/M6GYafK4v6GHg55Eq5Tvnpz8fkxeMxeF4/LwTz8wLHKEeC1RSuT+rwC
7xBl3SvyvXufNXY1d6R31MUrn+4OTgYpHUSm52X+3yp4V9emrsITgmBe7pr+WUgOFO8XDArYTw6t
3gF0UyBfhgjcldT00MNh6pFuxb5euXGrcfwKp4/DB+No02qsqXEZ4DnQhhsHxcUAbetEsuqE91xg
wMT9enxmvuWxUA34FEbqhL5MpLNIZjUJVi/CIvyp8QaB4MSKxcaNdmQMJSWE/ZF/4Gz0zjMriGru
Pgs3L17jMoHyqFNvvjMP7tgyUFlW8D95KrySMdCu4gb4EBToumIZlJu69ins4OuZVPKLTjmL2O+4
DkucqICcac0HvZMvLvyYkgjares56ewXjAoX7YXdlZ33c+wRmOcVHw1mqI4DXhzJu6qT8+iZPvfY
lhX0Zh9JpjXo08wXcyiWdwg+uHMplCcb798TOTVA7dqrXUePh9pUf0Ou1uf952feK5Hr2Mv6SCj5
y3OxLFJMYcAy/JdeF5VRYrPCJtMwKhuR8JNp+LpnrPFZ/BPN1IqUpaOjhTxoX9EZRZj0wTI8hgE9
CR1JFTDwLjpBSzfSYoR5jo2sgLh5yLloaZ/0UOhWww0FXYXF+zwU3g7rjZHGj5fTmqNA5qEty5Pp
tsLmUet8HkQPFEtGe36zAXFjXKq/Xs/OeJAVc/FMbuitUxZHutb3MWGxAuKfiD1UUSWR/U/Uw0Mw
FXPq58mTg/EPZ1EbBSYnQf+O3kEYHxvyJXUQq1jc9NttSWxHRhd1DqpuBjbwL3/RM+2xA8sIrs/3
0Yfu4QUl7Z987d49lA6WVanYLO/CIseA70BlF4zgWwYFc6hrfbpZx1N12O0UEe/ql0kL5h1G3ZB2
UMt22IUg2fxdY9QQHuDzbzxW90yyBVnjq3W1Z+NRqGPYlTy1z4SQaFROMbhZxPtbzoE1iNZllZVQ
6LetSYprOihpb9cd6Bm4szP0tq1LvgD2+77m+4fe72O9XrTKqD4+YSah/1+iXpTBLH3iO5OHLbh/
hjug62iUEHxF5YsPOm+XidYAFdnZKHsQ+Dsi8QcSbeEY4XhP2EML17RHHXyQPRxpNwTGZY+991OW
oAXJKcxSxcB45zHlmiuj8GG2Raq2SxLqxCUZXVdsN37NBqZoc6hVXvWNFUVzPmQZJDPeIBW/PQC3
C2bFTUtPnvnquZFJ4VpptaqWF68ACFXem3fbfmiP2Nsd8GSEwFtiPqi9yB0ZT+sDFeHu6ch+ydfU
6Vy/soXonISb5FUfVqJOYDgUkWMBL8XLLWXtJGT+1BfM2Nqq4TlsCNFASUBd+Z15WHUpuQ3Dkasw
d+nAxVDQTo0Tc66B/B/R+erel54vB+a3Vr9uQjbt8x2Vrh43sSYd+74rRYaf0B6oV7te5kGMkK7Z
SlQjy2EvXHEhh5bmSAU/YbBjdWHzsSXtlDLTxzuxN5+qZsUslQOCoat7iED/LaY5bOE8g28YXjZp
GLzS07+5l+4V77VkYo7o2YMSh1JeFrJw2/tGvjyBPR2F0aPoQf5EtcxPzoiQNjbZqv4Oxcvx2zJm
yiMI/29mpF6FlHnfzL4R7qXTuSUn0zDqsIFtHn7AksjFnvv/N8cQnh6n4P8yruaCr+7cptiIraXs
3i4e+HJ0ti7sI5ZaI10mk9sQW/nvZCOR7iibbZ1b/QSEgQz6r9p9kzymd0L9IpXfpDj43KHblqHj
+VAOLnTKVgT/JQ1H8I82+ZvEugWj8k45026xYvVy+IbesCnEw/l3rokMNosHOMc7CQb06bICFfLX
2LUbNiwgT9u9EWBdw/rypXFCizFG4w/QgIvR8Azr42PnH7sSnz2KzDw5DosYHFwrPIwnsh4u0pi3
GYqdADIoGx59UTr+hn3/CFXSarregG1+oEipPVSEJ3+s7U8rkruzjZyqV4NubNTLHu8ZjVawgCe1
l2wr0WIykfgNsNPuWJe/j1wgu2nctc8PgS/Rg2L+U4g9qFtvNl1SXYzYZmxnj4bWjetiNuNNPlL1
Vm31gwAAB7ueiG1snrPwd7wX5ZJH+O13EZqE2sElUk892CANycheJz+u1L0/M0XpnTqj/CCmcmWZ
9dHq+W4/TY71qpdMmcrk8Q8o0zn2eUulqpecX+2aTI5nDKlOdFCHR3oJtRnAAD3PyOjWZIbERzyP
LyPpRixFX/yH5VrEPF10fty3lqeiWa1acAejN6UWDjkY+3UlQmsnPog/EAx0osuUWlRIJAGv9/sX
g9OluM3zMaM5MYXqWPmbb4y/7yJYIA9CEqXRwIDT6JbJaW0eL7EOYjOdcbJ6zUtbIDBHrAElV/+W
YCsHslqZ/eyalpNcsl5aPA3gR3yIZo41Ztb1T1gjWrluEMVBfKabFiJhMmO/g82W/2ljR2bZ4Roo
hQupNyAkqbeRkoE0R6l+NDicAmFf3Sqijccg0dNe3uCNjgK+rOw/8jZsqRMZ6/x3lp+l4qpOTnVA
KxUftdb1TeN8liCDnfFZWHN9/RDyjK3V/2E0a5ChTGGS7LLtA2Lx4j3vBcpWj6+d3IF6OZhiB8Tv
zpM75ouLPLGqqYVUNqsLcuHtbhBIxKeCGMD7DbOv8v0a0C7+XGQ+zTYVETwmX/aPiuT1mwBWBvqF
c9OzT7j5RJdKQr+TJCPYvW3I2bHKLR51sx5I+E+wyQF9/3e4mWpHanGukal1zu/+Q0Cl9CfgngcB
3r5BgFKtUm8z4tjMNhO2l/PzIgU8DYAY7KPrvQmUpMXI5ApSN0WBfHzw+gO3Kc+kJGxi0sJuSAnk
7Gb/trWJBrVslppJtEPXb15v2/nDWN2fz8feB52nnD3k2ux3qXDutkg/bGpTjjFr+AwpObw2ZLTb
SNkA03YIDLUy0FDZQYWkg/USgFFAWqIPl9hFaZBY0lhTg1BUTLkNSfDd7uCpOT6vmtnDPbFTSrb+
LP1xxR352JNfM0GYA2uBRf3yifPWnBgihJo+JBODYB5eEXlVO4PxBXhKTGxRCMJdb5h0UqviQgNw
vlnO7OYL9GgX1AdD2cUuj3O9XItr0rZ2nf17hgCKxbnpLXU+AOa3/i/Qk8rYne3aSDtrj8PP3fe6
4m6T+c6U53tnIa0uhT6mUhdh+0z7T5pYGDkRrH7WcuF/IF78Q/1mIBReo7UOhfQ2NFBdZ6t7RjIb
l6/YojnL9JpGjBj7y1Sz7bj3T7BU2g5d/AQSPnk/5KfafcAS4CdGj2gIxzfZgv/cY8sIfDVoYRRn
zJoQuIch1NT0kWlnanSIhEfnbCLVFmlfeDzHXxQd0utToLV+Rt3JLcFHyGROcAZ86arI2g5OWrxA
8Shm6F4jFS6yTtW2pvgtkyOn8Zhp/WGLidSx/ChUIFm4SNobi2HmOZaLN4d6PSk1ymWBohQ1roKr
wy4s+Iv9cc/BgFwONyP9/x/TksH99Is1VPjJw4Uj+Q3MRNokMY/33UF5R4llK6PblBePf9mdvlww
0rB/989zvFQh9wV3SVP3ntvutOMNRRm1LXqUr5x1jqaH6Gt0NYMKwRY7/j2Rn1WwG19wO9YYg8vW
N20Hh2TRp3BceDJFTXS/bu2zShCWvaSKc3qGEBQeUpNK0DUS5YiCIVOE4r7nvrEpFD92TnsBYvyQ
X3upQpOcpMMoGmQDUHP7L5R7HcOrBf6f2wBEtZiH5k9E0v1DZYMX8HObdFyjeADwLFYPJbC2Zqo1
3/JB2vTUjT9Q25oKpvVhPq2baP6vec1NdN46haJpkyWMtiU4CCvHCS1c88jcF8LMldcW0+aO5gpY
zWTm2ri3A8oaS7GbJKBKtDs/ZhEF+A0r0wFarFgUCGAxR2DrenBrUv+5T9VXgSX6dVbgeA+ZhOyc
bM2xKKl+e7nEGfCEc9YaWzFuJHYPn3SsWUfT6pxnlAjmaWfUzDbwDQsnfjHewDQJU3Cp1A3YMWFN
1G8iNFuCeImWPqX3HbTG0v8aqMIcX77/Rlx+MYRZJ/lKnJd0n+E2sJQIuY7/JTQZPnw429Br4Kw/
eMCdodqTKJ6Hb+jo2LUXilWSZZTEnRMVWU6ZDeapGuM+RLZ/A780q6/EDD1qzpH40IjaEk7Eoiaf
d0RkLpsHbrb9XPI4387LouSoDARSITdXkijExtSlq02Gx3YRClEgdx+o9HwipzuFh4L4uOmQmeYm
uzxCkbaKAWx85LFvejrPwIEQ75wX62qAc+b5Hh40YVype8CEt1UzFuszdfb+EypjllCV2BOUXxBu
qdecpldgdGqclGCO1JiHtWdAFIeW5KI5HGvLfOd3PngLM7qb33ZXjg9HtIM7jJiNNakkaeUZcQHu
VNXkFAfcQ/o17chVCvy3XQR0xWevZlsGSatwT6UISCIV4CJ7wzaiR2Z0fB8TiTpLICzcO1H0AkyE
bPNvIdf5b6mExJ+759HjckjMi7BABaa2GQXk1NMvhrdgPtIt/lQwHvs5eOdgpPsOoo1qHsRliQUK
B0NF1Vlr6M/EUq4Yiji6RXMg8sbpUiB9NeOkd2/CAVRGJtKuAzaUUR76Idcl25M+IsOZyXxBHO2S
273MoApFOqOlGSE9GJd65ZgoPg4pc7fwCrVOFtlWAjgOmmC345ZQFEMV5gSvUP7iz1flYMCdBdnd
8GwkAzd6nGl0/i/rpe1XruKofooxl4n5T2BYv7Ur4b6mgUT3quKJ1Zpw8C+dZbwxl+WNxPSekB36
iTNlJnXhx7Yl8L6vf9p/0GGaAjCJUlj9WMOmEvuUC9LS5wpTjLRZvpVFnNLz++NFKOOS8d2fS+m5
oRetHzKZhbnmAtUT/BQ8uGGr0hqzQxY0InbZblQHvOVRTI76Iq/WBIAiCnOdPVOJbJi4Mvy6TRoo
czVY5pKCrWrMPV/x2HPzPgLRmdsI+2bFf2wwYKkWOsruk2+iLkXi8vAQppAMT7ma9/MlC3bztPkJ
G4OvDplVTuybECTSbYsKQN3zL82j2m3lXDAE68/2/ksnrJxDi7kGdgL9T0k37xrKM143CXR09mV/
SsuR1dLMFR/EuMJHmF9QGs98Oqt5JIblBhTtMO/o9xwPIR+1vaSfShOdGM/5+CWkUYWmZLyLD2zw
U44BKD4y/TMjhczKtlZlWJvZR0nTT2IqthdQzk0XQzbyso+l3Zd+Ld4UMOJjIwK4UrHSEln/E6bu
C6SwWUOdnLk7h95QWScE48FfRM5Y4DtloELA8pIQYgL+clmQ5qQA1Y6N3sDBcuVCHst4vxl5Etky
WkDLNZKMeGVnb6UGfx4TrI3jZGLwpL93D9tsGClUxpJgAkDNINoQFbMeA9w/g/c0CvpEJfnqAaRt
pTO7D395G+YDezsGnYVQ9nGwlcEt0NMUyZQXQq32DTevLmQ5OKquqV/9+vZxSLBAJleoFWs54PC4
dyQyigC8x4SS7P1C6brbT4jISo4HobFUKYqoIdftZobWO9cI6jxhKb/w/R6YrhYIMM+HieEFMCKu
OyUDz7FPzTlyMuAUPw5LFWd3EejGSZfM9ho5FSf5jGvkOutsxw30EJ23sVK+cX6zKl7zb2LUhlRx
LJ87eyhrF5CbPN4fALH0F9JyiN0cFZFKOPNbNYRqZ69P54GU1uPp65yMHRp9D+xPgoqHinxemvJE
PUbUAIFzEsqzvysNxpDqwfHdPDdbamKiWZWm7kLNyZstTSyG3k2VyE9uHPMJaeaJRJMx+RkNWV5n
lmKq9aeOtnNldVfsDUMturBJEMVU84N6I9eTKhP3M6PoanfIHKAEHAb1J15rbFzpgeY2nDdwvcE7
PfXHbcTbn7OQud7KrHwgCSnkmXUY1So39dvLBLPEPFI8YdfGFURZ7dn3HWwru7aIkDPD113xry7E
h1hooqKyxDd/gF8J4lDyOjt041oDvO3LLb4TYTs8A8PPulLJnzJmT6/CO3UYinZEpdxshyKE/STw
RrsdLBRU0E23H/jQSR13+P8ikNkDB6lU+CP1hjukCD1K6POhOwXyVEZMjeBql1CRU4YfDB0ZNY9+
uHcqOrLXaOssX0OhmK3R2FgLujE2OMvOxwYantSLv72hGCsO5kcgLXfCtRfMVl29hk7czVLFg5en
KevrpzC7VjnHLjLp0fU/Ao6j3ol0ZUO+SC5hn2HaKxmyEBcBP+zFP+ZwIGHWtItNItuTU39naRSG
hp7zXjiruw23o+p1s6pRJpfiG47XupzLF0ZKBubGxoKCHveh71GI0xlR4FbRWTZLxFVN8qLdx7yw
bGLPU8yCMDAT+A/LqqOi5JMrkWfbrDEirmAe2XRBxr4UOAx/nPCDR6YF5cuozVbnsNQIg/bGq6ak
Mv4F4Biek+cuuH4eGMwg35CwlAEIR0Jnss4PRgmS97JYtT2fBzUnosz8O/8bQ9+toAfW7TG5Tq3d
HJy4DupqN3yo8KSZJbz8Cb+KWSlxQwzhSApPwa595cnhtOBjF14sb6Z3z0mhIMB0/Ke4VXl1R+rc
985olhifF7dE6gzzTZ37aIIJj9cyLFyztJTz5boVbo0zUmYtpzD9fczjVjTunWy90fBIfTorTjWo
Ar/vAYDg+f1jBHVepOuIvjM+dbogqdXZAB0NcDl4ZOBOzZVEeJJYDz+4oVq1owC7yS1r8tMZ6aBe
3GuVsoDxzaOTeZTWS+iyVJdaEfFTkRqkZRodfgxX3kQvqlbrx/JF9xFSLLp0Mu1WJJA13W/OEI/P
BnV0me4pOs6NlY3UaNatswghkcTTkOV6Y1Izn7KbRnRPTlrSJ0sG96889ou2cJ1PTe0e11tAHs35
PpaM6im+2PHX1po3VeURaeNKCKVK6TjBy08cdEDvG72oX8qzhVh79cB23X2fPQDScXbxu8abDqxt
XyiVFf3YYvlYnEmb3Y2faS4OEGGpWlkc5SLKl8QoSPXnIpHfZBTG9B9BWiO0Gzyi0Ng3Ffa3GUuY
QS8rdRvP3Yi4pz8SQUNaGtQrl9Laz2McVZV5BDaJ3nwz7Gp6kmZo7RWgc5TzltMzMZjDyjNcNG8U
77wafKFytbO6bGb3vsjRmXZyKi90DifPYa2V6DQIuDX9hYzLk+c4db+J1F/ICrdkmrZJlNfcmhVJ
t5+2ilm0z8cJqogb8ZFROxlitCfZpRHBJENTblL06rnSn4G/JCnB/7W9nLAJ7rxja98pXLMe/5oM
nC6gf+pd1/TtQkQ97yPu2vrfs3wdFsLu/Wj5Rh7e0b7Ghlsw6gXuICD0ngXUtKul2C/a1PrmkJex
+PQm+DJ5QKYuJIuRYtI3dLShy7HB9UebwLvMK7/TFKkLCvDkMTuIl0rFz/tlUWRvehewVHREQU6v
e4hNrKAOYm7W8i9S+Gshvod6Dgc9od2iKoTR8WGW0BjclpAVFqsq9CZbpAqeujZxdZfIFo9oG5Y4
K3CnuGRjlf5p/pYTdjyAl6FIZFZB7fiaJHx3N2sRlIuvv/tcZUY1xIehbJZcskw57vIvvMOhksRj
KEUXiqI4rM/fyb2ANSvQs+0acwUettFrUiXTgFA9ixJY32YDeQPtgl13TqoLV44hP4CPtqY2wEKH
SxR4KG4epJPjqfR2pRdvmvtdxFpeAe06MczRkzHuG/Yo7xf26AkJBfY6rVJBVGDYd9sVKO/4IOXv
RyTw8LXf0fVO+nJ++405rcOrqsuPD9Ujl/dJzzpx+Zjj7SErxF9j/wBRMy8TCAxXBnucwThgjFa/
lCG4fCz60HwGcIJy2RXLIPC4peVFvfDJlVAizp0UY4NOsQk3aua0/tiaY6Hshw/Ur3M6cxL8xfXt
5VIzo1s5p1NQI1cgizI/6BiZPHnCoDZXqTaqoMZ2eMxGF3ma/NyV+3IFpASJemrxBIua5MtSblqD
S1luoXjeG3IMFzigvPeVtPiRrW0Gs/M3wLme2FpLToDMIsYZ87JRcV7rTopGxvE33JHLLH3FLtZk
Zjd1NOzGAIXgNI7E0URMEumVoZMMQQBRf4KGMDQ/xR9X7vJ0GjDHR0weEEfcK2kYEtSZHDBo9AEL
FNsUy5hH/Yx2omLU1Vglaazxlzo4kR5oqWqJiAaGDPw73UhWUIryAMaq9BuJob/MPYhw1N6I8j3c
WUTJONwL9qR3yn/XqBx2FXDrauPFlNJM4+Ys9KWZ+Mmg3vZAoKDKjxPPTvEjCTQrQF5TgqXe9Wol
NfcNcOEHwqucqvD83ZDA2D2eGetj5M+w1zV4W4b6QNIZ1TffT3lCOzzta1yQrgWUvhcNSHbXYB8x
uTwVZCuYSEP4Wo012Tbi2Hk9Ur0bMIJBUtB06DL5HNEYcXZ3+ToYsKiWLobcjl+MuqyyjZfnEPhc
OQHCXms4vD65lQvmbtjzLFYdYuL4DC8O1e18Hwvr48GChwMjrA2ZxNogF1xFr4+CNdPkkvDnOiOo
KvBsokmy5R8719D1NNuXgpnQwUU7UrmSZBpFPKnPwb5XAAmZdi19inOdco5Ch4pD3VgbpSwf64Z6
wrIfjjwrSwHhbpvSKuM4a2yPDFyj060VNjqLptAYErc5pkLLNNIMsUcftzGa72ukm/HKh8zM+oB4
U9DK0FKW8UzBL9jjwM0T5frwia+XOeRBuq5dXNPyCFkc7FdF1MWzCDCXfaPAZhz+q4ONmiLSS44N
736cYK8CUA+BIHHtJk0UfuCpZkU+DC/HrhxQMeEXXPUiuDtbIJYslEeYInmSpDAy6ciof1dz7yAH
zwQc7YnYPZdfHhgsyue8gFoRVLmPZZeo1iaLkm+rem392Dn4pZvW3VptIMa+2nQltKlv8RIFU/cy
GFhVN/cJehgu2f9egmqkbg7owLJTtfoIl8i/dYg4OvPmXeGPRkQabuPUo0a+k1YvqrSzYtNch42u
/S0uXUrDz9cnjlOQci+73MYRKuJBmn6bgKYr+70BRFGBfBsDc6hUz4qdYk1NR+xmXqg75mln+dTg
W5FRUKg7YFBqJUfY5GoO2UO4l3G0l4Is9STTc/ugqLaRVTunjGOdsZtdC6x/7TfgcKfKIDbhGSuu
rogB31KQMRyJA17khjyXeVaidFST86wmvWMXcke0WW0+qA7Yiyx0BoKiNMlJFqHhV8yw/oZxhRJk
hOx2XKitnvRtsTK16OpKgrGtoRFlxKCE2g2nYIcOOGceAqPZjqVRvuMwgS7ATxmxxtMiXat3Opko
kU7f3EKNV+2yMkMRJVGsTAtWHDyOeMROwyZpbCHbVJTgwU89wxqicbsdkpsmplPeszY98m9xUcC2
e1TiAuinAiy5JszuYhoGL1Y3o/xe6X7SDkGQgK/p/K7/ZV3VT/ttpawcARPAEqn+izcabkmU939i
YeJS7WVYTmzOC0WQBmXYFVEL5htzsbtCyCRoT4Alg2UDf3loVwoFqoNlz+x76443hJ+TbhHQ9Zm/
AAJjhSbq0AF6pYLIHaMizodKD6DZQQpbxsdiXTHIc7XjCZqD050BtLChOa9u403KEqLwJgq8cT8L
HdtwLSHwIft4S6Yj6dbySeOmfL33YIvsF9qyHTs1FXMZgDukUQ8LBzhSgqPLrThR0C2gEKiKWhKG
uNR/NUERNssKNKEE1ZlOYZkGi+PuR50hTS8rJn1REngm8pcbzu1D+Ivb7VgyxDZaOluEU5143b6b
miJ8NFwu76d+VHyNePTe504LYcpAXusqmug4TRnN8ra57/wgM18qN4brfIBcLjlnNxk51H5PdG5x
i5qPXeyN9gBqtO6O/oNHz5WmYw/iJPB4vTgQZDjmNbhz76ApRzPV3C0L6ItLyL+a3YqvTOvqX0Z+
UwFjwWYeyhl+MXr589KVEfwLAuytkmfidBkFsOT+g0akE1PTlpt4hUPtpVEhlKVG5QfmdiKsMe/v
nDvPMmMVFBzko4G14PJlR+75AbXG34PoFFHgHuCVJYjsBYnx7hLbYk1fn4mHSgUccv5Bz0t4Vrdg
+anW3Ctv7u/EOyMv1SxqRz8hOQEG5NGq+nvJEd02RzfuR6b5AZAInwXEodZEc0fqH05HHuIHM6J/
LavJjQyXQpja6jUYK5zBjlN8R8zBFS836G7ctmNld2UkLy8EokzqSx/SHhzNyKWSibZmypIpwU7z
SyKIMH87+dNmUP3yZN1Yf8AD3lAcEqdqV9jDNLBatg0/sOsapIVgr0whH77AQSsctBmn2o310r6G
y45h5B4vioIfT+5tg/S3vdsWIa6on+pf/ust/c1sEfYODRUKtFqBhZVj4ad8YMYq5uuB73BT2ReA
A8Jm5RU7XDM+6ICwZW1N+UouBrGDSQemxYK/QnBEaodZSB6WPM6A7AyVkWlMEVHWBlJDNmyhoW/f
2D3ACRyKKf3ztRz2DUZsBNKCYXHORIBMrLh+z531NtjjG2uh7iE0ny1OLeZGeRL3ipBGbTi3wuhM
X4JQPAIZSCrmR97TdYOHbWt5YP/rKfbNIfqmUBtHo0J0MJtxSyL8OgvPoMjyU89IIBoHebt8acHc
R0GATAKHxWV4EY3bOlVPiNSCes0HrJbCOaoAc9fL/i4RomKUaPm/HTtissYf1HB90dNARveVMQJm
tplojRu/+tHfNuq4fnDmgRCOLY1RXr2PC10qbsXd6IQ1WD3dT6OkJNalz4SQbLoCP/QAzpcHYsvm
tiN11bfJNeKVzE0l4AGyoDEmLDdjsBrA6dpBp3kWWaOfiXxRjX2ZASPOCgRXWywjUhIdSrwqsg3l
CuauRa2OQ93X3MrV127iYK/Vi05HwQYDm93rXkB5Um7KinOxi9KE1pFfQG3Du5+TiSe7bMqgIu8V
nahZFrM9EPhqT17PRqh2I0nrQG7CwJkM10rlcdLHNZmQOpMlWoPpQTwwebO1ovr7+rLBDtVL2WIS
yOFmCndwe6iOjbw3toaJoTorz5Ih83R9GoFLrlUcDkelsrZRM0V87Jrn6xNwaFJVO2PdM+0wZsLv
ucpDFuT5L5NykktGQacLDjJBqJzi2eLWK1bkjkNG8OcIAplcYTPsxxnH2g8zwG/1OiVtH9pxcgEz
fLeRl8kiYnplVRqfsT2A93GStaRT+QEC4sQMEJO4rKwiqpSXlronMsegKDT0UP+ZFMPE3ULOlYh9
YrJIxJjTN0lkxdjP2PMn5g/P2RfcgZwSJvFPdwU8kLa8saagMGuSDTzeK84eWafnM4qzqHnFbUl9
TEHsUbHsvAWyBPFGycEXkT5g1NXLfyhFf6goFBYwsQtfChwcCNg0IcWkcqczSsnDc5tp6AnNMIaf
8rk92hXeF2EZTRrb0/jwTsuRdL+S419JSf3D4G6eQl9aICYLXCIh06XBRhH7txgH2nYjo6eb6+FN
QZztv3WB+eQEBgfkl7VVrRj0zKVKSeD4O1nNpe7JIO/LvCaR1GJtY7Bi2ykthUZQGBHRfh/dAwTU
LCVDLIl2K1+PdHXhnlKTBmf2FZv7UIQ805cb54eb2/toWUlUUfQZzyu3n1IyMwWShcB9gg5kvMml
jXBAvYL3HCvggNIxQCGWyaWx0BDQRwBTTmZgPHsWtQXvhyu0OQ4pKlQ9V7lBeHhKeiw7eemNFhrl
nJDk8FeSAzamqtXnKQFD1tvzi1Ji6ooT+1tuUQ77XnuOHvR+4b/lqhs01iyjh3ZXCw6NARWYC1r3
GwnEJbUONmSb/K7dIxYJ1GhyHEHei0Jhkv36iox5PPBVBlwY+MEcTinq4Db/+jnOigOU0vCGjsRv
VXzRUQY/ex7hnpHQOY4pSvQgsOkrgh/QSTywLtLIyDg4L+6EJC6hwkJRUW8W4BkwntNKjg4pfCo4
6asjJOVOUIeKue0DCAOzD3swIXPXErHcNBgmJKr4mkWEnspnGeLLZLW9BQdvmsmw/uY7bOzaENAD
muO4hyo5gV4TSUHdbfLrfzMGKEQpgVqZoZPvDYEsXAc7GH4q8btnpASq9ngHBVj8xNF1XAc8JFiO
DF9tLjlQWCFjSPv2DxyNrHMNb106UN2a6O5wr/x5cPM/2WQm0oS+ZXcfmmYCGC/q9okiN0Who4KH
4znqHsS+/DlRkQPq8aXxSlHS16tZQc3zzctPQhkpqWAdJmYmF9pUI3lqunoetSx+Js6IV8Tqrjct
hYSA2NKkfRHFmsxswTDKfFlVnApaBgzoRjZLlyPBgeN4AKC/Jtfit6TBJ+Xkd+WHlPz8UktkyRtg
fOWwjSlWkei/9/sij+Jz0EUU8Qjneht7CeDbs5pojBwrKaTKVLyYSO4ycoNDbMFvj4oxgmfxdHhl
9o5Sgb4GZPXZ7MnaKwFe40BKVBZRvr1E58+X+G1k/1zNEzsW3q5/DqJg+6JgFeMsCqBpf478BmoN
0loD3Q7c63EC2UYp2dFhzN7R7IIYAPl++8edXX9OGJmzqiFIRs29IDoafHl/uhsN6jgfnvHEF0TF
LCYRrIo0K+SoskSowxqVZvf36rTBDy1bZCGVENt6Ht8NuVVu/24cNPEefl7bKcFFEVfCnmi3GtTn
RhSNXW8McrWBblrZPD4v9Iiy+teVwfx9sWzAhirzqpoqyOPfADaI93YHNkDsjHSmpaFk7LUTRux6
RW+fjWgN74QSgd3W0HNJvr4oqeLC1/XguhO/HyOlXr8m+05pAkmwDtpSb7j27k5e5X6FnOghsIEK
4wCgSWBs2muQMbqExHIDraspwnsuRSvn3aMeNJfR4fIO912sm429pW0Z16vfSclL+7yW5JU0L06H
TTbaupdDkzQDIqSSKQGE5Lh1vkUzrXyTzjzLLzbhM49UYWsf2AzqpQ6LtZ/uZTZAMIXUGxalBbIT
lxowGbxGPnYln1TfeX+XiVXrJ9jq//m8roX1YSDcmj7x8F2XrM0/hi2erMMR79YCsxLVKBQarmYm
PlEDcp4NAkqKARo8Xu+R2DdMkaJf49c2rdxhycYHlsNpRMhs9HdKgNDVTvfv5+yWDyCpv78FubKE
Cxgo4bPddrINOztTz1m+3FLv3Q4rO18/B9usPjcv7cTPr2NBqzBLRRyCUXhHWj4FApHcmnNrw094
of5ROl+ShIVTxNdBYSh1N1wLB/FqzSVLhP+miKnNMwcXPxEMb7/0LpCUNGc+z6Mm5pkw6xNWWXq4
dOhaLIy9WqiAsE7flpxCFRX+T/K1feb0DQs1Yo/NFiBQW2aWsFKcIbe3im5gISXbty4IN3HkDhAq
C2YI+Oo2DUhDYDsalgH2pKkPuFiLwD5GyT5qDocboPHsmCC+hFdsTCQbz2oOWbyvKR68/QvtzHzP
nrmsUh/77o9mBWxMw7zpLi/NEfZuAeepE/EB4hqKwnqPq0r8nk05Bn7icA53x6v2KUkfOwD9gVan
WoMkbJyCO8ZEqUhJJKQKcCb8OQ1dm1QF7yVXy/yE43C0BLSGFAauBZa9QQl4jUDEaKzb6wVvqxwt
4JN/E3/WUDpxPS59PDI1vD3DtsPCEG4ZVomBRAfRHYvbGlr8kIcYxKrc56PJRV8XokanlasY4SSZ
8SRrsx16qoSTKIKfUck3EEZYO3Sub5lLBtiRZ9soq0toZVpbKIEcNS6ewxxl6/7SPaPCT4DGpYNA
oGoLbZiSrS1urumzQJZs6MjH+EMdcR+WCKw1jhKJq5NnoLxJWGzGzpfrmKzGmZvFDBaSfR8m8teP
ec73GekTmS3F6WDNT/cded4OKP4j9e3RwVyYKiiXiSKPTKz6BOSj5hUs/v+ZtN3vPuaMVw+zaCtu
eBpsILCllHwWqiVsIgqd/YFZ9mDhZgKB+YWx5Txka48vAGXS8csdFfgPN11tyOV9d5h6JJCuJRPN
8C3ngs95zwfdR1ruKgcK+I+hkqBzs/4ac+9AhbxzokNiUydtDSD0+VUW60jy4kfIVVTYjI933OKv
nvHY0YQp0tv/hxjbtrJieoC2i97SU0NyaLVf47kT1ptGemBnYd1czg9mlmIZoJU5EbgBJkeTGCsf
2ow7Pr2a5T12poOYegl3MRA75I5RLSfASIY3ayaiuzL+PwTs9nTQLE9PCdsB/I+nJ96Gdv5q9jFZ
dAt4ZMnpRIgHKCkuR559xYOiu4UDZM4qDzinzNtVKC1Y2aly8rbRqEMlgiydfvZ4FNsEWfdTvQBI
+BUtNLjzxaFv7O75EsA2lKnz4sG1qQAv/CmZZswA0WeVLd8AoC7m17zzhwcrNiYzuJVa3YMhl6es
8YCr60/HTmpuDhh1pIjNdTeUza69OiWQW7Hinty8FBK/iuIt0yJEyApsAp5OP5opQl6+g09Fcg85
oRE6w8o4LSozhLj6nYAo1NVZlPXSRQx2KC6GIbz0vCKYrgkPT7y0TM1UA3vUpGD/cUZanCCa7Nkk
EibyISF++XuTWhRzOj8F92QUeeGaSQ0aCp0+5keZmJK5CE3eLx3eVtVstWNpwO54yscJRKzofiM/
RE5outf18vK2llJy+hQrb3Fkm3bEbcTqd259jSaxIIIbdpATh4Gjq7CFYVpKDjpjRtteNnWZeid/
bYy0XfIeK/sjavwUEimtHXgS2XLO8zLYHDKCqctmyjaV7ZPMvy4ANn8u1zJqto9sInYx3tSxV5P/
kDGNXzusGkQqIg3uyZ6UVwJKgkzTcihgsBSE84DhreNLytfa/ImU9qVjFsztT7MepSNjz4QvnrIn
/PsUg+78Pd9VubIhpYTifPg82x+PJZ8ddKoewGxsBvgNF8+VRkoI6S7BbT/KArbjAi4FbXvbMzBv
Gi16y95miE0zWluAETph4zRdsg5F/50lnLdS//zUk1P0ezgHtO5ogv4UTn//PzSHdCTaWYobBzbe
OzmsMrdvDnqzAN8VpTBKRM5v2EkvLrxlCNzzG179kQqGTWM4KBWJFZ0NzKpVqXiD9gVF/xoq8TSr
Jl0EFlLdkMUWDuMB8KyTe23BoYEotOdH5+hBeLNFH06enDMoEnLRteh5Tm55Bx11NLfBiJR3oIaB
8wzUY3UyU5QdZ5auDpZvNX3Lt6D+wMXNHTZ54piuua2pjBliIbfT7Qys+EZlk6ZxHljXz5dClT2A
Bkg40HIgrqn4Yr6muP1ziCAfgiUldxzIwL1Aw8e0FHvVcU7IOnj+BaApw9rcABe3x68EMIrScZv7
nV/qNkaggsoGIDMT68k03jSyNLWCtmOipsWT7Gw4oL4MQridfH7mpnZjonx9tfnwnI769j3aZQ4K
ogxMZgVEpag0GPQLxGRiJeoxx+tSCTTeGpvbcd+cn1Jk1q3B6Temisg5VTtClyTtzGdxSIG6Bdgt
8TDffpRm7CNA8K4hWT/OL/IsM1HgNy7EiHBVzpTmz87sX/+Dk3dmrlBGRSUtl19LF9pQAlTh68Vm
K2ce+C1pwxNojVet7bfqdtrgKgy/qV+YIAEFcAqGtE8Ncw2PDsCsUStERZg/rfFq6qReoLPMJdB2
O8BCnEzGdGyyZzMvkQmRsowuacBtfG8mxLAPFCCVYEHcPR++ph3SZqA5yLPgalTgUBfQ8RPQk44T
QW/fSoBMDeY2QUDH2Us5AXUMIy0TgBLyZPgbJBm4sheu5w2EBnCbRvOixfb9dbRQ/PXioHwkZ/CM
sAq0JZK/XkQx1YFn30EXxtatmCgjWyUuRbzKMCi8sNRyGodm46I3qjw3K44/I9WIbexOmw5oZ2lD
har1JvxJ8NzlsVPubiidVwEq/sDkf4pN4QsmZdzsceBcI3gyX2cNCwHprfJLePPvessEjMirXZsD
wVMAv1vyXL1hQqRPMA5MdFR/UdyC/eoZGu8Wd+BJNGRyuxhOTfYE8WI2Spy4iGyKKSyb8kt8yCqU
QU3Ar0p5Q9Pnuff4C1fAZmWQTiMSHZ4GFqYrkyV5tb2j1ZCdIpSipOQrMLaKntwi6gtMaMmNg7LB
4FfSaK9/heeksvKhcS2yrg01Iu1WjAj8CHtbZHnE59v9wYysyRqivkG8a7ajXtKNCpAdxkLleEOx
lgq6VxPw+2MHacGLoxVI5ssmEt+19AH17tYs3S784iPsrymf2rvHRKwQ1Uu839cDNCtOMJPwg159
zFXt0jgAeF6WLlLEnB5oEmvT1rgawfwqaVTlgHcuLEBm8tJOpRA8fapys9pC4dGaKJUg08TWl1ja
y92QklilxwgbSE9bMBYRxR1yZ/JjAjmhc4CbPRUIMP7TlCTqq4kXhZvQ3vCbVx1z/qlkyCYEGQnK
Cgtr5LhXyRkyQGXgAf1sk+vCibsAVuL6MBSnZdPunJ1Tlz9Pg16rMVavBZrfWIe7dvd6CnX5HrY5
ksB7Stg4oQusg+nVqSxik8Yl2vMhWirQqySRt+mYqWasfUNWtEj9z0QLbrhe4ixcp7qxm60PloYG
BYNPS4N4HZpInHABMlX5+LB/ejhOxgqsZM03S1t3ylTqJNwpG6r6OzB+4LYBRH3mf1PKvnnua0nN
sxJuTPqtew00gPyngPMcKwzWriVPr7ji1UAogkqtZfG3CCMePQQtESXyPe6SzTv7HJgHrF8FoeY1
biFYV1mT7PrqoSw681fn4JBAZ/SI4ZCkQokt2UuWZiEOe1PBnu5EnPO0njQazmT1yI8f0BPxw3/J
9GAhuhImPOtc2MrLAsjnWmLEYp4+B/8gAaNy7Cr9X+UehDN1bwwMWJrRd0IXwBoph6lVXCvMibhs
DjO1nZvv9qeauuoGGZbRBaZvHeCfc7BsLIHLquIzCGWKY3rQCbpn8b2HW7GWUNvgo1egSe4/1fcb
prjkwK3UK4WJkjSdgPYbfwFvZSX4bx5rhPpsr/UoPtbj8sTrb5VE+kOVigIsZgUunTRVKTFRp3iA
ujQBX61VXnFHHb8QxMoXNOwOYg7ftFNs6S+RXSQLX9HxdXx79vFTbA4P3zl/JmDlLFD6pmA7dQda
2ZJOw30+Op28RyycjtORVK+JeN0hdHkKyb0RS7HqRUFv0QO39slZ4wnhPSz1Q8mZCGbINfH/EZ/i
Wo4NYEB7LQvFel5nHiPGHOVBeUR4k5n6CMDbJ3TPOC5+BO/WcjM+8Vq4oz2g6AQGik2YosS7+HUb
4KKC2XGLENsU/yR5CAB9ARtqRQttlCOpNM1ApDoX4TOcJ3IlB4+q+hxolxqR1F8/5VGZEBGcGFf2
3psHc8jzs6g2D6nJiy8meGGb0BPiwDGCNsyx1sD4EBjcs/MfNbVjs4w2lfqXXLC91YepoqvTzr9S
CDLeFNiyM0LxydbTgBTxUusQaLP6lOUZKcNtqHtsCzSXn9jfiNd3cxVqHC4xL2al0BA7hxAOLnvl
fDmymEY1ar4gjGv06N6LFed1QacNnAoU4O3cA4yHfvadQk7Oo/0TBI7Pj50mX0hBhmrSC96h7o/k
BO3715hnf79uO3V4ffUFoGCYhqM6eQwXONH9UkXJ8Huvsc5rnskNgydoQkaOCauLNqsMdnOmSqFR
zFd7aEuP+AOgz0C9vS+0cR0Z5mWmCBe7nSvizOOTdnh1iK/ccIhKjNt8Hc8QUDmCEhrDBYICIbGH
1AwETNxRyOXZYgeO4pnegJ38FlLGIZn/kzb1RGul9gJIicKC485qItidfiNiExNtCHpS4SSp6iIw
Soadf50CVWPF71OF8+rGabGzM7RsK18vBObtZsMexkOpufaxcJg0ijG6X7x75v3saEpIMKH4maNP
xnWNSQgsvpRBQ6tkk5gWwSmKkHwjD5B6C69XbqexvLhpCNx7fYwKqSs15LCeIAvFOQJrEl0+jYAO
jqu2d0OMusciriaiHee2jXqaiH9rjKZu6uOgejumZxLOxj5Qr3VKdOeyYquF6lDxMOd582yxn/qS
0/tEHuCKoPEA0dK/IelhcoLGxeTdj7n+eMeCtyD9JZ6LQD3J7Mo7J1KpDFhAFfXTbK1jq/j6Q7zv
1sv6qLVe1Hb1p3RPCYb+P96OLu3hFy+mZ4DFSqYjA1mfCgHcmI0juRBsHEdQGRVQnZd3NFnvEQUy
vGt4Q1FL70Q6CPwpsJmRfyqwsCW1CawrkQZlolxWdIqIx8YLiF2Atfta+mMfnbH6stRYoGL/qohG
3eCF5w8Evk9vfXu9wFIbj49fQIEnD30xWxk22zcASAPn3MX9ulDUD3Mr71sIhvYJxCnla9Xb5flU
j6qlBdU0y8R01JgiAh6ciUZCwBmBkim9MdZnVIyxknP/RvYUPBg3fIsp8hS9GKas9abA0VfFXWlE
bjI21sae5WB6UMev0z02L0saE4Ugx8ozhQUn6YQnX1JyFdflxQ54upxtSQtzYvPY+m/LNmG68LOo
GMn1aQwE6rtfpnrV58v7fi+NkDffnhidLpla0Ztrc836gV4ERlvLMp6jCUD7sGkcwJNrYQ0IfqyD
Z7E0k9cXIKCREQ8Vyf6+M07g/MJioVYSSg6QTTA5+lvRU8raZ4YGi4dZnzChbFCHK4LTGcv+5sHv
PZSPZG3Ov9d739r5Xleu4kP2v2fSqzF9DBz5jgQ29G94x0lKDN2Okw5WYMo/2c6JzBr4kLte1FlF
GalZHTdAzHGaXv3yd11IzF2lez65keGTTKfOFHSbF7FxzYqgWhar4KqQDMHMsNoC7sUZeiVpKCdG
bhZ1uJWWbuohegnLeq41NkvFnTPQXdIFRiURZrS3tJYuBRBODQBo31onNrP3OyG0JNsP6QZQpUKf
X68ZcTk+7oBZxji2ZdLPgxdvO5QjjFjZVRxCr2QTiGp4WuTa0Mwr89uhmrz1dDXNC0mrWMOMTikP
91HdhPQIzQSaY3xqsgEvauZmG9gwX1+fTiRwt+ckdLCkgMBX85ZBh5btfBmS1DJvKNnBWt7nNdX1
SxZIsOQs0DQKFbhJyhyNXG1C0qJwp4kB1Cj/6pSRPiPqIp2kqLUdaviPzB0F64wB3fIZt8Lodxv2
HuJYAXOxEdFw8KqonI2GNkn4l60cVDCIrC2je8q0ztmRir2Ok/lik1ZQ4bbVRsuNk4iJV22UMYRy
YfstueOod4VfTzUb96SZcN3uhLDI3J0kelgHt4R57oQ1yVJybVIdF1GzkwE48KGdvkVodXkrjhbm
Mi9tzNutuKBEUuG/f8P5x55E6HGd1VcAUV0IueNj6AuRRq3S6A2jBYfdTVizKhUIC2/gZl5+zYFr
39wfUwdPVFchr1gNozcIlzs2UHMkn+JXb1bgMTJINhdJbV5/IqcycOU+Du+vqvReN9OVNLADTkSs
pM6a2Vr7pDPvz1sfI8JaXFnHfNZS32v9a/r5PNn3QiN9Jgb98s957Y0UxSiGckT6Iv7xc8VupqFV
OvKCLyFVUNyTTJ/idlesQBUZck/3R3FKIsBBDpy+hmSPMUXiZhe++fksKRDJ5/M7rXGgDC9mguDP
BOHAgqHIftw/HbjDqsSt/MSvCPdp0PMLZiWWcwQqyYI7O23w6XFl5WOMYtUOxcUtyCK2VaDENZSx
CTr55Q+QMKNF2eTJTBy0byPttkh3Ymdsn8VoeyAZDI8oRTkaLiEvNcHr5E9V7du3BTrK6BB7/ho3
y5hnHNu7D++taNVqrjzQdXxL6a2zI1vK92xY3fhPPIHz+532WF4hUN1Ss9zxPdzh/wAwljs849Bw
yv1pcInki8sFYzm/hIT41HqOvMjtWUXHqicuSVS9vSmrJ/9njDYVxBu+UJzeYKpG5t2nXvtwK5Ja
OJhpF8TSvtzCz9s7bdancftv31OQJZyKKFIjIL1YSkAsOT98ACeymlKLG2RYd30c/ms/NvK6Hcvx
rxBY354yW7JA5v+KRucYKOhcoRUJTszgd/poiDfmvXNbWzR1gz1d7k4ODifFQoEpZt5kEjhhtXEq
gApv8oN9rtVjTuHXx1oEnbndxfzZeWyFHFvjih8rR7cKUyKX+jdEQywPLDZpNzpEjYeSre/K+jLb
yiNKNLEwWcP7PO1g3mF658HRxq7PdO0X4xKUCgvT21g0YfB0Y9s/hN2PU8AGrMnoaXFG8eEqO0SC
pZe1eSkEoRbsMLtdx5Uohq3XtDcOHyPV46GKUyP+xwJSjJ9VgQyoUVEv6bnpwJG0O4x311Vr+ddZ
bigJPCrtexXAfD2EHCWTnP6gQ9kufxIUIM/g0bf+s3MsM2nVxvEyySgYUykGTYPiqMmrCNm1/gUI
NlywrBbUoi3fTSff5oa/OwGuea54Jqnw4rtbm3hvkbtojdcbEHg0CN0144U1d5cRokbQoOJVnwPS
cG5MEnb0irA6tMaNm3eGu+YHj/A6Uejm2sK3JtH5qUe85ctkRYbkvENlB6PnbArZdhOtMu9MjLHF
o9iMn403nhyNAnaxe6z/9UQAK3Rafy0PNx/rM33kSrrXDHDmHR98iXOlJBLbyC48GethfI8mBjZU
7FxQkMM+4O5iteuCvwX0Bnz0NHTTqAkDqFof5qQHIVdJzeZsoTEdzhcfQGC9JCCKbzqws0cx2Xcf
Fi/FsRTgVX1M5IqhBKU8LaW1aCMbRImCN0Yw7UFctPakenqjabKAKMnwYUM2ibWytTrhl5WIczaQ
knD9sTECvNOdP+3u1ubhW0n3vnjpSWZoATUMBeVwBtEx4J4A8dOiQ+3BIZAwLmI9VMF700IPC2Be
iDoArpBjBR70D2O78Zm/16EUjrdwYK+j0sFzpAui8TalmFdimE4VPm4bRUqQ9mn1ckHaFZJH0NbL
F4Y+tdjlM4FAyJQiXwIjRcoGLTWOcaJE1fzW8Sn5IQipUPdANqDtqyvcWxtLV0KenVocsq5mhjy2
IL6h9TXYPwHSVqT+/o6n63TP84I4B/Z0iQ67RASNMN1ZqcgHNVTpPXeQORaZ9ATlkviYRA2eEAc8
8hm0bxLbI1S036dFB9oRbMHKs/guLW9iOdhwNPRHYk9hom8u+0alj4P81dxrowZUVaRYxZh+4xHZ
5HXr8cQJ7h6EYzH6KyVPe7uG0FLJhHms7W+ff8gj4DKh1ERH7nGTBy5SwKt1t9+gGSoyqjqyQ9x/
bvo7npWj1ASUx8KVJrzxI8h2foRSyyZffesY3Ji9tKZyagu4mKMsFk+QP+qDvWTynGLE4EfM4Tq0
I3BRk2FUZZvzTTRoLleUh5c1CZh0DV9L8nzcWkgJJKjjn7/N2opE3NWppTaMzmnAnKnYLFxJF651
L/LGWmU24MEmLPwrxjB2psIgEkBTcFhMEQuQaNYJ01JFn7xa1h2Gh8azIwrMdUsqrbQEweeBaJt4
9Byc0UHLVNZJv0QUh//BvCYm4jbLyanJVbPS8vTtUa9OuMiAhskVnOlkHuVBc1b1GwqtqHIYBxwy
+EvE3XdT3YBkt//oanHXObMavrj8jSdbslGWNgNue1Z2N2rP6vWCAJX3CcznnWBTu3vwe27zPB3t
29NoU7x11CAyQlhgAiRrSw6cTztocxksKkGtIYCMH8QHzx/Ptz7Ytul+Uc1jKfmCp+g98T4GF1W7
A6baK7TC/35qxAgsmAhCcuAE3BJe5+3SAI0hvyofqD5hfmS686F7LOn7Km8bYrSKntZAAyOWH0/f
XTYirP1eV8S7u3J5WtQv3aGGpsyWJ+f+PRg6iROfe2fFlckPuYQlGY86hz8PfqL0ZZDXKRJPFyVc
QilCgV1vLPc0wvaJsrGjiDJWCApyPP+Ua2BXRLW6pq7wcb1Hcskzfn6Hlz50YB95XVnWjyjX+TMs
u6QmIbn7NLxUETGVgKbBKeT3oRzldfjBvYht12x0agimFCFHEbOlYknzaRC5SF6w2yuiTTwwgd6p
59giaHxG9MXYjxlIOP8rnuieXyNWVMzR0WJOuaVfifPfvuD18BGPV7jVaFHqx6dNSBJ2Wl8fgsD5
ou9nKCTrDSv1Uyhy5JK6W7ihR7SpY7+VeSG/gFQZMGnNOP127sSyO1jm0mM0ht9jWQW8mbSN8GC7
qZ9MAMn0A1jMcQUQ7AkmbLWVzgNeULSszojUwuVvxNrlBjcAVHWCx45wyYhly5ULY7RED1d/06Fo
Isy4zY/ckqyOqkRBN9PsqwGmVw0TazyHrECoP6eZj5vUsTZCpFggPpEEMAVlAQzj/9BJP+adGjC8
iW4gPcWYEEWq9pmgbkY4TR1rbJv3SUDe5TbuqMSHja9/CQoNt2O4Lr/3fo5JE2ORVuzgC6/4yAUc
nesi7W4NRtdGfnhAdOGPvEHGNYzZknb1ot6j7ON6wYZsuyO4jxxyy+nyfAXMXjirzx/eYxj+SMK/
l0hVTCgqZ5S0AmUN5j/8jGTNHx3iWTCyoD+gbUlIUxTW2Eh9VloGkqiU97dXgK+vHqcw0MCvq6aB
qyYevl6d+3xojAtFAD7iu9Zft4+WIjbLvurt5oKAd9ZhqaNGNxIRX2nwIx7J7obxm1T8a2dG8+fY
MFdlig92RLHolako3hoYU5WIgur+/0cQ0CzMehELC5M+mmUGxANzio0mfZ9hF7kXZZQcu6FbUhzH
HZxIB6WHXbUXEoJ8nqdfe6IZfnaOVEs1aZKLULLaFTRIJOrJJmj4j/7rq93f/MBB/3v0FQ1oIrNA
PcB/FHybyj/P+TfvndY0nfF/Jedu4GCVq6/ZSSURQflD6txDC/7BNnwOnfUo3kkc2aYnI+aOuULt
0LMBGVSdYZr6xlXDsNXhNvsv3Boz77oYLPbxmISWDr/XWeaxdUCIbfYuzY6BC7X+tM9TIZzzFQfr
KLa07aoB/hLL5eca+EtCZA1qMAtCEufxW37TOHEtszQk+e/lssVyb+vsBhGPwtyWa3YS6bQv7L9+
U9iXgN0khnJ8YUo3Z2dM4CnajNryNa7627hCd7EwWe864KdazIffgdq6wdPwWE7Np0unFwsyfMd/
ByjA4V27/SpNoy9CNIO5pk8nIexGQ/C/3ceKXkJyfcL41aRYEaziTv/V7KGN+cLHyaJe81G/SKwf
wjAiCSk/hP/t9fR2+66Qon/daWIBmojWwtcKSe/UVNy2F1lTpA3OCd1LtON3Q/ex0zo1pmMG3Ooy
ePkrpJ3KvDUDYEN6zFMMmvQLuVppEz50iBvw+ph6vLGDThYSY9xXYwWFiz9gLNf1vwMdr33GiYYV
PR95Ju2bVUzu0vHRK9j/xZxHEFpbVP0qX0KX38ykY4zzyoDzw4oTWEGwBp4DBizykfZmVfKVFCZg
sk45VZ3PaB1ZJPj5WzBCGjaGSpneT5vQHresineJW0cXwgtdI7beOebHEakcfGcYH1y8ZcPwYVmq
Iw8+WMLrAS/m6GHdKZiBWrSbd7YniqdIgvWKyV0ikkfvlTGObIQ5IDUbgh92vqBdgoyi9GpfVN3M
4DRk//3LXMEx6pViB5MjVclpI1uVo81ndmvmaANkoIUIfkwkUfHerZ8bojK5Yfg14GBq5nuBfNst
cVi331A7z18AhQnd3d4joBlh4SnllXHp9bYrV3tKo3lslZeHhuGw0GShdxKRhP9nD8pF+LIQuMnP
ot515SEUvkP1v5mFNJcCm2HmjQqrntXGN7/KeGcLoW5SBMO7zrk4xXI4ROHqIozdsGE0CtKwS91c
r7MhOxAE4jz6OSei1SuDdsN5A/ITOcara61Fi7N59BU56p5lIh5ojKXAYkIzmq2gduChQD6qkMk9
tY0NfNuSs77l3eUk24ZoEhYWureuqRrYtGg4OJ6cR6pJeIb8iWtvGe9Y8+x71xI4g7J2xdL0Gigt
SikJTeRbrUr4RQs1j2MXcb10wBd/lXBuW8omFVRYIY/oenNeSpgBkcWvJkhMTm20omUp4noFR92c
4Hwy/48mURK+ad1tkbrHQcp5GfYAqzsrR5iItp6aArlrNVmJoj9A0Jh07GhCSDZ/vXYRRnrqyC+b
Z6sbfWE7WgJoBL1eRGSqBYaJjsbQHXFfvY6D3Bz88XFlnOjtWxdOcy1Wcev1YlZu193vfqWW+q1b
3+ULg50FyT2uFTQTaIxc0bTPobxTYO5SKiGPrWdVqHJ+Qd26Ke8erUftvi3aIFccNjAT95OhxE4a
n1H3ufQWOj+dgI0gXo6voJ1OicvQ10DZTx8ZrRQYC91t9KH6OMMjyE2WPQpEtSv+Pkn76uFf7rDt
I/6ZebrVpmYOPZx6PK7RaW4C2Xq6DZQa1XG3Erk2OV9gx4NqJKi1bCRAl9XynMW1trOukHnOxhbP
+Nl6UivMnP4Fdc4kgk+jsPBuXIYjFwms7iL5rDkU18E0Dmys9J9Pm84vA1F95CjkM12F81pbbcPU
vgaIygFdB03Pna+Ys6ykU1lVSxGHLTjBR1x+VqhLGpjn4l2+XMD2Lqn+UyC3BWCgsKopwN5gejQL
xBpywsrdoRsvI1n/XnJsE5Oj/ezWyOtrumd5IKDy2tKIyEVF9I7SbofSnR7rbAWnqVUYneUNvUNq
8GkzKiJhL2P+8zFC5KQdzUhaoJKHrj01B2CNq8c1HJFIV/x7/7iw7h5prbsSANTp0tUNXaguzWXO
KeTavN8dyNgw5+OhPaB6BQerJ43rin9JYbqPqoKd/IP2so6f2H6yBkNEmOG5klt8StQwgppFyPnW
nD52WhR08JNEWl/Pkwi9iCgs8HNCNN7CjkvfqE4EyTto7kHxVUtDlDaTcE0Flp9l2jG56VTF9zKn
e8uUS8Rt6FNdhfx5lT5cYLkDqXjwJJ09J2SS8e0bMo/0F7SaDLKcKuxvzeSApuXyokuJzNzx0WBz
YwbRDDXxQnSyC4bhj+BkfRiMhCr3kZ3Ln3TLVuh+nqqjqvoHLDFbx8flLOfPaquyTpBmgjglsy6I
mYU4BmsrNgUbOii6ZYSZCCBUJlxMY4iat1lCGLWfmxR2Gmq24xrIErYqJzkoImXRKcL1E4008QbE
mvoFKqtxXedYDtxijVBYdZqIYWH5AClwm0jXntHcd7d1AHAEQ+532kxHEIEAQH/AfP7hK37uKUl1
sAAsQIR0D1mbjtLx5OZeeaGHIe/zk5Nxm42JXXgFAJsrg4WRYv9DZMyzTclYQkt19+YhPmv9/5h7
KA0jGGDJJv4Dzcdk6Zh4QFXd4NkiVTKydON4rG/Gm6Nfn+5ktEfMCy7Pzon0Sasqt2Sdy++XIgh0
INLijIydAGRpAo24r0mJW6brH1mE5un5gj/CUb79MCQnzKEgOS6R59rGHM8J47ytXq1SRygorRC2
eaQilX1R3jGcn+V+W1DSM4Z8D4dk2KCf54l9Ppy2bmzCKL5hkKAtVSundEiUfeZeqEi5xtdU15of
8GCx22Dy2yKGNZqtg2OVv60RG2BUeTpEm6YXhBOTsDOrk/s2eezaBV/eepgk6vXUtYbZmWmHwx2G
Bu+NZo/INQpY4VfiNQyiH13jCD/eqoV698nhvE09xqBV5546uAgaCBINVbJ5Aq089G5+KRIFi6wF
31b/ud5FFc2+z6anbSuXHZx9k633BmxqbbJqo0Cy3fmsXYFkJ0lfMi1h7hGAqjCXuxkw2D7mCVhc
Ah0NDv4uvdT+neVsys2FbKkOWbe/LrMjednUQlauMLy8IWCNRp4meP34TMnGg3Vh+zFldnKnI/zo
eBmI2JDVIFtXn0mWbxiXGtsGl4U8m7HzN7o2OtnGBb5Ju7RDTjDBRA1X800e6bWNLrgB4v7hlXQY
96d99Fr0S6bP/TWjYalF07J8CA45cfq27pnACIwaSAoy3lp/qptEh2r92Op+y30k44ndlZbXF7FD
nCNw/vuqoRa5dPePnMeuMhgXeEmzDMVP3MXSywg3d14LYsu5ljVdnsrPQCHfT2niQ4DyAfhHCPYZ
FGbMk0d5f77oQ+kNMDw3cW+xOSL51+Gd/6h25nxO4QIBnV/iYHoAR7HiYQkRXarXsUULbseOgymx
fpEbPie2gQVBf+aAf1Dcg9niZiGSVR6LtjCmlciUuQcU0bd96aGfncvG2De0oK6mSSfYHypQh/1O
w1ZUoUXBWvWDFeVt2gFJu8V5Z2cA1JUcjrrBPdPIW7o89zI3F/02g583s00JlKOzoVbtkd2bwN4s
14k8vBHiDbqTs5F/gSlyUSVNxZeq1QzdPjI6Sxm/R6dXpbOaYoNBINIfnl3UhHS6cQy2aVd/zzM4
owcWhQ1rTCkuL2Sm3Jf6w5XQwOIXyd0ogZcybgJqWJ3fLdO503YRdVhLUm8S5q038rv+cpgsm5/+
iaWXxvWd0DmoKrXZPeTHcURo0LLzsClvgZbQGJ/S7DjilpRyR7v74gvcdiO2avOrQEJK5lkW1GAK
76YP+ZroAw2r8ohtWwrTZXMYhYFcf5fBNc7xsl+tOWjoIlPcxEUR+7xJHCBVlU5mA24aUEnKXCsz
4NcdB3Q3U5a7zt/AN7LEXCF467gkr2FQ6jtUFKiUHgzS8FK9WFDCvyJhqXL000JT+yiqoCNUeIYM
ISd7p03ZeHakNqbuTQyqHGGVynxFUAMwAI37hUkIClzIRTn/fkWwdUjmr5t3yZw/GVP8gy/aii76
SLXhIaSP4EboEDGWaMp0Cl5Jyfr2jX2hdBy3UBjgVw7Ax0KyhWL14tLTMDcXrtDdlvy8yUnyo4IL
186VNL/lzhVvR6hNynVFdbPgD2MuXACdO+Qtd1ml0lp5w6tKV05oJWKw4DhNwizO+8THMywo7xXz
c76qUYec2w7VzPmJV94MCeP/otFa0ASSKDTJeNOCQap4UpHY2UtzBP0ssivzxgexc00lKNGOvoKN
vw8nYFeIp/CF76efxMeOA15C13ojqgTF8v8zAyUfcWfUcir9+ArJoZO1EDPNaDJBFAU50VLCfjGa
U33sVOAhqju1eh+/sBJ1B9SKaP2duOihMIh3GeLTBr7aFDcULXISg/5ktKvVXuSjY6Sl8eqFuWp0
w5Vx1lajNHeb5XCcVeSoETh3k8fdPbLdhu009FckJgN3B3WXjJ7SACyktkTdHYgz0XAaG2TJ3M4J
Na5VLaYixHqwlPpeGhADDbzqxXehJPG4IdI+VW5gjMu1USQpq6zKJ+5RfS3dUyrSXzv+uqk2ETN7
aete7jzEYhUyben22uhX46ijk799VOMfTpqfBDggh6ywgzHbPRa4QAXuWwhiBlFCcmb9urG6JD9a
icAW/kDUQM+tqAql4gkRvTpkpckk3z2knoE8iQ5ourwn/HixF2n/LKd2Gpvj+mkuiEujiLk7SfZ4
hbLF9OD3h6zkxEafjVftGdos23H1LCTViuK03fsjyaIGKWCWsrWGvdzGlZJuHz00x+LsyJ5Zss4Y
xJKL2j07S4auiGwe1x95rItUo9MkBZT6f1JO3bmMDjc+Ten4covDynss+edA+DrkoxWdwzPHWGjk
sgBQ5xYHEARJ7VriSW0DFyfHldVYAyuvjTaBln0UkHwS/i66P2JURhZXxRVDh7cr4B6A62cBP3yr
s6exhcZMFCnkH7xKEexh0J/5gu6b5ALaU7RHuWE3u6hpsNHJeWFCtWAC3eFlVpKj6VXSunWmXMqO
4gmhqziqOcrByvZkFtwgKkQmj7V/kfbF1L6ZvAnuyCxqozhRDE1EpXX2HbsIjqBizegYCJQTDceJ
tELNJ8CT0zEgKEq8K9Z8j9qJ1Ib9i/LNOwPGA35RxqLgtvKWVB+/2ivnLOJo2R3jk0MgnfnacIJk
XSkDvsdIwHNaduuIfanlptBlgXj0o9N0xS6qqmOHFE5RtUWdZmm4WAgRI04C0R39PGBOgAM1H6XR
o7Jumm1dRvgDr7EFpP8CKKwziNFGFbGzb0XHETSfVj2UmjNIF+EfKI9Q7v/2QqDQeJC5HsDb29+I
CpVsslXanV+EgJWYyOf/snTmDFob2FD9RcnofM6Hb+9p1JnrCpg1K5Ju1jr6g5FLs3EPgRVsnVOz
BmOFLahI24xwbHaImuqhkv7+AAfZ7lB8Me5wOD38qDPFgFJ73X8ac59/u9iA6u6QuCfTPjrZCLOD
K1Kx5ePLlY951h19kW3uuI0PJxfGr6Hg6ZgdCSvqmSWwKmC6bT6bOKsudoqGhwdKJ5fEQjoVawcM
GieXVVHqS5rBTPnFPyPGm8uFZUdTrnLNK3B9ncZdbuidvbnAcPSVqohtCvwbNC+4VQp69Oy2qxtA
shd3W6n+eLVv1B0ByrdLI0q2LbaCQgTiJljhGAvFzhWm/V2IctX1Pvg3+zIBEpd7gE3iAagordkZ
UNGj8lF6SoewXAUi8pUUWDSTGXmdglvVAD0xUXg42MWbLkfWy7J7pv4oOMDzzGheUxlOUzFICgLD
awDu+z9kG3qr9l8UId/EEYwt1xDLmyi+YsDBPA/EsAMarCctsrdF2CTO9l6sxDXA8pZoImrurMQO
rYKOsBWDgH1H5E13+vCzao9CK+ww9pmPPFL8qukkKX8hgr8SlyrGf7MQ9tFxfSdl2SQ+TmwbQl8b
5QFG4ACsg3sU8hX5jkVfPnNxiuyAa8vrCuBqnOeK7lWGgC0+D0MyZIYjc1i1WKEMW19BDKmVIWEW
HNKFZ1AuV3NQKZL3ok+aPyj2B+5G9NeAUokAA5/8r8O+vjHb2oZmc/qlg3gHYsqkBE3J68nHC9VW
t6KKneAKOjwnr8ewbY7MOb1gQHrghk9h29H9H52g6zpQ80cCw/K6dnjxbcKrVovd+5gtABCa6KeY
nLz4mEVzEGeQOvSemKkRuTVWj8bIyxvQalqzl/PoWhTlZiuGMm7f6I+Uzx7v+540zeB/f54Qgxhw
uCFzGVlA/PUjql5x1GKlJMKICXkldpXAiNoH/JC1r71ZSX2VlouTGuGZ/2meByp5TNFFP6QbyBFy
Kd35pzjfJTbZpdGX1tJSpL7bcX1+5JmP0rMwUh6MlFDxig2UnUhFPOUQAppeUBnEK+14ubKIRLGy
ld5mHQ+B9IIhmhEkzwW0hzWLIJ8FSmVly9EL209LbiMs1+zuIusl1Bsm2k/ZF5XOt4p62/zQksm3
+PkVjsb5KSR018LEHo3mIhnZGTpUoaZ5z1hChJQRnkfb07om1DgiiP8JZXXh2tX0ZWV1bbPqfuPo
ixsVqFSwQ/6yBwFc6RhdGKAmbpikG7PB5jsNgDNuIJ0kqN5TwTIgILekZFYftqIeD+Yn7OgTlkzQ
GCaJfH4/tMGc4Qdy4RPMGxz/+rHKbROLf2Wbgy+tmCO3RamofRb15ozbtcJwH53cH+h5Y6w+Qnvd
dDGaX7wmF5LyvWKV8WjRnnMDh/nA8gS9OGRrnuDRqlMUZFYD1XFyuLM7FB+bGVHXTl9AhXBefY6Q
f9krEy6fcA6c22+QbaUdglpsOwSbnl4lBKqzECixR7u4K6LDFLmTYPJCsPqOVjdgRwGcry9lySTf
zmVsehgcX1x7c71Wa9AcD787sAGgzKLZXNmYbGmSjLRvyzErysTBJYz8dV2zDQpmklikZnpunxuc
OHKiZSDPxNC1IVQpAs24iXv9+zwylBf/KWb3w51I/QOQrEHC+z9bxBw4Qpw8N34mG6deVfo17aKN
l+aZ7GegNQVBTmG2kuyQG6VIwyNX0vIYrTjCrORfw0cHLarbnrMUL/DLaWLP2ttWGraagqRClSI1
duxZz/LPl40GP6yAnhbYXapV1bg70SMeWtXhZeqO5KZo90c5ytnn7XKsRi8/rFRhe4NXCfimpw/t
3JNi1eQu+TsR/b2Qt21AXd937BBWuKtlgwV57iG8KC1tUk3ly5m556kEp+PlI6kFLIjie9p5d5yC
IlgaidqWkm2T0inUyRFXjq/FHn+WXYSlbtBZXrHfU3vwRN+lWEH2lTwkvHDBIzEomWcWRX3M39Fk
pNFucu2TmPPBqqPpunqQI3+EY0krbzCTNarc1BxtwpBeHJevuUdAOWRAUwK/SI6spamXh5l6qAP9
6xawqKhhJqal+KXfaeiReUuYaU1yr/cLJYBOw2Lzvr43eU0cLuQ+HXo5sSuyHN9EgT7dL9MDo2WY
r2VJYzYYJS6FGS0BeZ+oqpoubhhIdNDAd1Ww36spyH3ukmtRkPPEWkmywBnyg+1U+cy+ibX8FH1q
afDo/RnDm6ituGGxTQ4nT+3crnPI9GjKD9QRL5xOtwEA7Q+ecTtAu44awWTit84D88IMhwDwLDSj
TFVBQEY8NiGhSsX6dasAWeOspUb8tt0Yh4/WbmlNpijPYRajH2MXBGD9sKWpshvkYAR0r3t6mReC
J/eFc463kZOmHQJnYzVkiGWwfO0HwocQyKEjxDQyA9BeQ8H0AXjAFvRnjZpC62KBqFijUBA/b7AQ
rvCXoKlcHqvKN1DBPgRab3wXGkJEo+WMgov0s5ub1b9M9tbtmfoJJMFEsXrRs9LdqMAXNCy6lfRN
UjraPjtGYQcPL/OkWNMvaNy/v20Bi/XFCNvYle+wnts8+t/TvZUTfAxBPQ6d98UspejlegZ0b/x4
sH9LwcXTyHtQEqlrZWbtiYwAhAGCu2bTh7h9czQTQDyldpVuIKQ+a8+hEVZUgEnCE3yhOnLONKc2
hi3aexnU93/xH+Qe5VgmkKXR13k6TFnoJLGmeAX8PoAgKgVmbKqZ86GP+oNYd7YvpBN4BStIauJq
qD0FQ8Ks2leI2buxx2QQ+dTGlPNgEZZlKymF96a50fUarw47HznsZZ/Dx4sQ/+a+LXRS7qA87/R+
mDFOcVU1HlI61SQi/ZLFRxzbnIrS0BZ5lZ3W9d+T5+aNRsD2eLbZ39a/YcFf9VQer2ZfoqY45Bdk
VxJUsg7D+5enVncmvmJoM2F/A1uEUsCXc3qf8jqMlrfu+252lZ+QyRbM93K5MhGx8QXHvSiVlawB
3slO9iru9mW8Kp1RN/mkkxnLwCL1i+ZB9AkwYVYc+6422wX30an/5Ct7ViSu22Rf41MExpOQoaB4
sis7WnY6wf2ZyssWV5Jc58UyPEvgPVgJwRBt7Sf0v5gQZsnJ1PlaPAGNACb/LTzGVctUWh44sXaz
+rw4GdaetUrGWYHYSHn86TNSnGz52jneeiEwP/jM0GTqphNql5nhgkhqtu8VLv2isAWFGy927UQs
0YJTwb6u9g3ZmVLiD7sbdQn6V96HU7453ODXJhXETEILpmuVGyldgR+buYiFVfV8Ln93n4aRVKeI
oQbVmGBGrcJ9TYg5VR1FWzirWQLL1P7gJd7gVL8oAEWiPqnLhrs9O55ardqlR7wsSs/7vkD3KLmr
ThTA4P54OvO9GmiWqPuK61w7/SFYGUDx0PIglLukRApsTwIeBBMScOtH//NuePi7TwlRmBQ4qYQM
AbA8v6Fw/CgdR52lFMHJmjhyQkqp8XhHxOx6DhWRtDirqlPurvSeApkBMlG165T8f+B9O1PmQ2D7
4ValGoRxLyQSU0hA4AUr8/yCuHl835iDAu/Rn0he1WKzCOPvRPv7bEQtmRteE563dCa5vNLLbksX
UzJiulzyX/2X9H7l4xBCpRfs14kMUgo4NwKvoFWR0+E5iiPm2evxACBHS5aUTX96p9R4+m6rKKIh
VqoWn2t8pL5M9MSsIF66u3tiCuCGxEBMX9uDtCOAMvdwjxwGJ1IDFA1Y265ULDsNfcCQig/Co7LW
AtNk9MIwvT/eUVIED5g7ekT8JDyyl8IZKPnKnsdmJ9tHHaMTerOlcmVyb0J76kB/4JmMUtGo8arp
ptixxtnE9folePL9RzJx4dUtLcDZDRGyW6s8Fqv9WKxo9v5CVFNnd/DZF1D6dIALgF11grOQnCvi
uwm10yQ30eYa8cbNX/f9Xt9CO0t0GmzLBzqz9w79Bml4t5Hwr0B5mKZxWoDOfI6O/5BVJh2NQNaP
043kNKZM1nfzP9BgDh+I5vvRk4BaZjmPmzoOoyqFI5D53XdoMtT/SGHTzPBEmhSgpSMJwSctjHNO
UXPXRgTKgoYxqtltRtsJFVd+oKDmfyNk8qvJ+RTVsIr0DAcCzp7jYOZAr3hFqz+D3kX+QcLg3Ktl
15yo1FM9TmIh7lZiAhmhVVJVeDzmluv8I6fkMf9qDWnuYHSx53DhERgA0l4oJXdQvMEY6juZCOYT
6caAHvq8Sjq75X71hGzSIwuFw0On64ym40SGBKQhBOfbMXyK8t5gBTyjchyuqpWQ6NvWwyQ+rfho
iwh9U7hU2/zIVCur2+4JF1JFDmKd/XAEs+NIu4eWrVvHTcg3/QBq/zu+h8WowHgPi0+0ITCpMpB5
ze5TOT0RxEFvdDh1nswC0Bp6+IgkRQDQ5RLwKjE6eKl/NZM9Day1N2ipqUsaKb6/AZIt6/FKNjbT
OYThbDfpI21AEWDPvi07WHDBNixt1UR/Z5ioKO8oK0UqQ47kxEGAyM4BzN+Jc3MwN6/rrMw93geb
0dKVcRqRXJTBOLI5ocopsxE0e8KnBmKJIWn0h4Yi7NhH7IuQ0r0ntJSBk3HCJYU9UK71aIZ8lSVB
Gr1Tmqolk2w69UgGcFPn99CmPEEL/FvJoh1UqDopeb6uXTEskkdVJ/xcOfKJ5cf1SyqhFs0ySNub
gtvVJJfn3pzZh5uDv8kg1B2T02QaBndAr9lgIrjkQ+NDgdo/NCr2uYToJT5HysrBhsDMfC1fEAZh
zO2dE8L/gmhKqSK3nRw0yRKVuSWdjk7EQE+Nqys7ecC4sPKfegbmN3K+4HkN4QQtH3OjyLNcie0B
/Hza9aiMRnjW0ikjbRa26/yu8YuYCihnr5J5PoVNUe1TvYQDZlw/sZHTHNGGJIT5cVrHMoqA4Z19
7/JHQJfuMjeKeS+pLIrBf3VhkJjCSssy8GCU/KzVWvB3tCTHJCWOh0Qr3IuEibWRR4cR1o4GAZV6
o/JtZ9jvIYuFGIE4DUO7omOd9w1YeNNSvRdS0zf1YDj7rUVfQm6sy/sXLoEQGa/i0gASxpIcWuwP
q8PBHIBZFmTA69nk3zTY3yj6xnTqG7nnfAHxWBSz0HIpg1+WlXH0xZUvOYO2fG5KF1nHSym1yisH
QCDhTa2yMfrePWZ9NpBIjh2L9aVm0YHeHD6+kspYCBygZ2Wx7XIqT7xmT82Gzugpw73sEV0zoxpJ
SENAwRpRed8gVBKxlGnvyBYlX9iGmxyI9BDHFZWBCFRL1HUZROVWVA6r82a9x+nO0PH/ZA0LzrUJ
MOXQRAxZJfe2DejogbJ2pjVP3cto/j/maMOUqfawdtwauovm8XJpCC2D16sgRx1mx2UfzOYKp/g6
W+I3vlgMPWAhWEfhTVsIU1UUX5PQFD7MdOVXaieugvqYQ8TpI38zyq0O+eNs/iUkgoiT2Oeji0vK
9HpzGIBC8h6BVAo9CSzGt0TrP4Y231ik4gLspXju5RMSC6Y88dRf75ri9HBy/3fWooZloqPTNLiu
MDqk5UGP+Weo7CDWAA0994zRfDIc+E7OCVg4i8ng8C3ChderhEyC/6uAGQSSBbfgB3tWHtjOXWPt
EGIwYYaQq6C+M29fxE34kpcRKVZqd3vD6ElK/Pj/q5xWh9+tGCgWY/3PAgd0jvaQ5d5HUXm5wvca
vGflS/XebUL9xUXrQT8MhnNyYlZOgx5ZoAOSpyXyJt3JsFCInVKBaKMG1sI8z8CZdWAfv66TVoxl
BFJokUHfGJDP5xiYcHkOJHpZGoaBMbnk+1LrnciCFl7UnukNhgHDHErKHxPweq3XTMjo1Xwq8Yjm
A4ngK8ND/nrmONhnkAeaaSLJ+OIqySyVsbHSblS1ErVji4fZN7q0Dv0YXhe51dwYWNxzIdTpcVT/
uG5DxHWx4QqDAjUY4QnR8POyZITb5VvKKrmOEZAfNy4M+nI5gaqYQWx9BRgA/gfrWigZvgbcxchE
5TT8Kf//tErTP+h+x4mO84pwalunhKuW309eVyfiXUBbMJJM0I205mgYobp2Jggw64q1be7L2Rse
sxAlXAPx02X0wMWpEohzBNFpaQPJIdqMBJnbasZMxISIBMKnNzxGbhu8GRtOw6lOqQMybDTDh5Gy
gNrQDdbVH0tKwXi5GyhQIYHTnNs5OQrBRjOeIUHyg9igYmCvd/N5lOCITuMWw2h9dCBWzVQUnfW3
CKb6ksRWSvqSOw6Ig+eysETbcqwv2KXkec1vVfRdz1XjTRmuD4kE39WpXlvvkRVHr4B4bua92w8l
klPbMf3jcD0wiGqj9cMUBNyOyd1g6RpNLNO/kC5i6cCBG3lYc6DBIDJmlr8ckUyq242wLRAcPgGJ
Jo5A8kIJLQ6RseTbF8zFiyCo1n4sMLkod+ewLmhTtWM15MWoi/0bba6B1l37zCcdj5DQgMUf3vzb
XGhG5pPHgXLry0TOepmSfYyrSO54NKg8ihK28Nv7fxQm0UMsSOExol7mhi/mHoMMot+YFAdF+OXL
ubLMQ5XrrF/buL5g850wFVYuU8xNa30oMFnr6qjGF6HFHjl1vPadcx7+I0Dk2WzGoRw8/nEbPMmT
3IZ3mumZFJmrHatZOeE/fwkRb9i+cqpjK6JRza8sB8F830uZqmwIbqGesMvlnh4VbsMSx+/twt8z
2BrdODVP1Mnzx8uzzaDevAxFYx13wa8JIRsbuGaMqt1+6L+rSCY3zSQutVo7kuMpWAU5XBYfYVP8
kVVyaMWLXhXBMMLxjY1s1xgRnyFKagS8ztSJbrftTBd9f7l9LtdxP5f4KCsLRRTGr88eAAydsgtv
ug7NpAhMSIPW03h4A2a/ikXwMWO+HmxOWSgpEGV2A2DYlsIoXuIMTMSQK+6MNJv1g/dPOWDntHpQ
K+6GYKC2j2mfOgRgjleg3yEoEUmH7spv8JGDEtkwNupw19hoP6TY9eaHXaR/b9WJmxSvugv68JiH
nU3v2sCDOu0d+hJA7LvOsnCnXxMJ+I3/esIhRumhSoAV8TfvoCOhTlh8ijacfaoqkBvr3I5tp1To
p7yZWW1F4/V2gMwd+mNuCC3ocLrlZXa1xMaxa95RfBpF9kB4ILNucGaFEhTvCfrq8mom9fFufdyV
2ZRFErKvqNeaK/3L+0PXexClGgpycX9uOHfxM+Tu8sE79Km25jKEYAtaHcu6aaXv+gTB9nl021IH
Ylay8U+YvalV76oYsy5FmA2BTrgoamCYqacdYeAYK5SUZ9rsbFFP+ta7Q+bRrkYhKrWvLFkAbfxE
vSzqyBs3NGFnXEnhqevBT86Aryqn2aAwNNSxUEd13OI7xWhCfle8Xn+DLmxptyAvhI2Tllkpf5hx
pEZmvNEcmdy8wKRQxTEFQN9HPMABbQJDqiMONmzvnjnjbSlkKHiO+NHfuFesdjQnpyawUYp8BsDv
b9arjP+/fNJEw02xg3ScVCPj0+TiOsfVGHgQJzIbAAcJUy5VLhcDc90j/ubSv020x7bh62/bUNrA
ApYviqHNoSrlZ/5K7/P/BW3LBU4AAU3IYw1rsYSDdNkxF6sQXowfHQy7D/nSarWGOgW5Gt9SURh4
U04BpV7Ynv0VsIJCvgMzBGDHViAvctddszfDT+JILvibxgAejxjFTOgcnyfGyxWVwQhfqpl2DGG9
T1itDfrr9sMUYTjRVsSNuxc8SyTFMlFEThJ7lK38VIuRqJYJPPdDoqWhuDXuZTOkYxezcscKe2SP
zMQvt6/abNkfSOT9E9zgVIgzx6hb5GXoGMsP3CGNhVqBVONBxQ9BDCg1GKl6YNPKJE+j7FKFZ0z5
T025keuFVMQMBNsxI1zrrTx2Ihupm+mE87FQ1gVWn4+y0OZ9xiqi6mp/mvuOz5Ugg+79Js4bGpDG
sqzwgrZ0QWANnqQ8DiZ88ZS7gVXoSUjue+EomYYfQ9N9Gu8t/gSTAhQdrVmJkF5q7ZDmggneh3tU
OfT8xlpF2zHeR5Qse2QHjWPSdGC+5zBhxHyLc+WR5ORswexOm5VlP2yAOA32WxStJZnFkcftxvvc
pGCn+TBzY4JHPSGHot2ir/LpWVuLzNfV/sax7UDZDIu5EBJHJA6NapxhM/e1sGMYahCfz4NSuyAy
1nkPwKDmwizTNMaTdoWuvwN1hAPk+OZG63V8tt8iHcixOUR7BkAH4+jExJ26skX3FYLeWjxA8fri
VkJO6SbxXqeGkhwCQ24qY2peONQZUt2f0OtOJNdH/MKVV4GqK/h77UNCtMgxFNNDN0kSSypDU+cF
lKVqU+Pp5uStYXY4t/0PKz+UR2kXCD8xRHGTinOyNG26pgfjqgdQxnCVg1XlFCuBFAfPUjVjB/MS
N0qmAPfDuIUTVksJ+N2pFoHP2dAconxj9sJ0tsj+BQYeA1KsahLW1lIYW2a+M2a393a/T0BoTPIC
o7cl3TJId8TDV8lkzk1Ew/t5zdW+1oVz8RCrxbAF1NgDaRRQwxUaqBO0xA13Le8ssx3uhqjHAkcX
/crp6iEZ+sqNStc8IDq3D4wGhC3ZOeqUkE5xyUQtoqg8Y7Z/PWY4iQxvcNgCls6KLM+NeQMdqZRr
lvoOLjn7KbNDsk9dvscNW1sx5PWywifqf91ZCz3lYpjoCGXobcnHbNtMe8JsViNZOGukJDcnnwbJ
KI5jKGz0sdHnBggZ75g5VSPm6GK0n8nnklN/jkfFC384PrnybMQwo5V6wyceGvLYvy0hD7OH4zzS
rz6w8ZgR8BRJFsoXUsGEPsAWofvqMl/qXIaOcuuKghpQp7YszCQboMU2Z8TPaWpKL/HA3kZxaGiL
ZmiyH0X2HHwvNuIWzjRIXFomE9NxXeDrmNF1YYrvqFjXsVIPWb8jO0Pys+Y0HInaCYCkxmquMdD+
HIGjH3wxg/Re3IY7UrzhduwfawbT4JUP0A206EB3h90J4hCYVTaOS8KbNJGDsuo5D+aAkZJrW3IF
w4ZMar+9YN1AmUtYqDv2qRcgT0kB12u6WFL28XjrfQyY2o5G8Q66xEYIksXalrh767EevZoZSHTH
UG0n7BdMC3KCaFYGARjEMF15wLmfAg+OyOzyalHEFc8MwqjNVO6WoDyNZPCnnQA6K7JKrjrtizhA
Mk6yGRyvS8bvPVXLLlT0rgtE+bpOPpfn/Vi8SuaTScfhFl3fqPD9aBafuP/wfCAnO73L6/wf0RIV
fxl1fdjbvRiyBpxelQuiCCKKW6lqyS1tPKuQ01RJKXEz2cIGFKFN/Paf/4s9hzMmP9U63qKVepHs
xjUnXDLv0INZWbTorUuWlnQyb52iP8vFp9ngkmeVlyeuOoz25/n3R8JXmCGaotpBbEOTeJ59dROL
e7P1YhspmCoGqhQMvNSEs0G4jVwPrUp8a7h0DOMw6UBruCV8lUBr1MK0J37XuHb355wOwT+9TLmB
JVRTINOhsqPNONJiZp+OpVpqBUVu3F8+EWFY9uAQOTo78dySFvpoBLY57a864/iajg6ME+dSZuDN
cfVH+SMiZ2EO+ZdHB8Fi/uoZiLL6CCFgG1O42a4/EibdNRZJM06OKE8My/SohXxNE4O3yBA3DN9N
0wYBATgJiO0ScQN9nFeIHskwAquBkrYE5l0K1bZQYscbay4Yu5DKR/yY2Issfgi2ltt6L50GQ1eW
5ZY5qEmOY9Fo+duUBIb3CepJRxnBZvU+1IAHaciWUh0qsnVFOkeqg5iPX23mWFarplUXpuT8yR7p
/pCrhHrwLtoAIdSQbqfnVClthWigcFvc2w83A+mCS+uP4uuoXDokrKGgRV5MJ7/UNaaq9oJTQxme
LjR5KhTw4RT2AwONQwjNRzTak1AaH77N+esI8s1x8oA40VVaq2wRAFXUPwU3BwBXWLTNFnZZ714v
NnuitkNVOrsiXe7HgmLu7vb2eHsAlfDuKJdhV0Q4rB0uVvpFDsy+Zkk+ldVrPXHLhHsKprPBb9Dd
25LPHANMfaYMz7jaGuVkzRo+KxbCl2JSZBf4W9CV8eOpOSmvEKJ0o5nqsG8Qjb9rqrE+WvAMHrvd
FVpmFdkO63JUaqe7XejWMq3myD9HxKGnwx/fzSZyxbYgBAJk8aSzsUjZoXpaJvSMWV/Fc/dXjc8c
N7HYuzyuifU/aS4h2DQCWH5apgu5tfv8kRv8OUKRWN8VQVlWB5ytIr30WUTOAgzeY2+n9OkaYY8l
cxKkrkl8Fuzaiv9Q426Dy5V/EIc4gFbD3GFtQYS9siN1J7tSOQB5VXkXVieTbd6k3DIDAYEI+Bj9
KuyJAbt8nXGa8CiZYoKcW3Bd9aj5SncNnTtqG4aEvMcyJr1GFbWHGGvirXqXibW/ONuow3+FkVQ8
+hkfBFJRI24lYzjH3OF/NNA7C40rtH4HfjQpM39Hle0ymXPZ7nFeF139OUqTOwlyfJUl3MXDx/1w
slUW+yrUD9XP9qCX+KhgE/DddcCvPhV2YVSb4iTsMriLzIH+XCl8sZY4kTp61Qw6juiZyubt8WV2
7QryjftfNCH5OmwdHPRramO/YfFVjtmvby/YYoblJaE5kWXabgfesZtoQbxAvZudzp4wPqJ6UzQL
diT6phl0l1M84gi5bgYPUu6m8FZioxQshdlTpXbQ/88Wtkx0PkAZdGwIj0VNlvDrRTZj7/eX5lmn
dPy5mWg8rmk6boNdO5Z581RdYXF9YuHJV4t8+s+uSpvoxeMWbW8u7JC06HOqIHLyfRWrnmHtumYx
n/HhusTK5GLhWi5LAUyM10Sd7RdJc8p0HOs+E6xvZ+fZNNZygR6raPIexB0dwqNt9QOlB5BKp8ro
OxXAW1A+d0GDPTpDbqWK6iy/tb1TWdsGgz8jEUb7sAc2O3UJ/CM2UXOxZeIIv0bksPbihTsf3Imk
7Lv3pJqfDDr91TxzYrnYwFA3HGLcVuZiPIk9iUpf/KAKMxSGkcvYmJ5fulxOB1Y9TgJ539Yg2/JL
e6lvaNMed6UUGcOlAnB1KWIwA02OH2UEpqeyLdi0srfwstZ5tp++mgLvByn0t/BM6ZeVD5t5CoOg
UWMtY6x8UwzOKJnfVRT3KRfOXD2n+Bd4a7k2QPsSk/5cIiSj/wSyNXMrQdPqrek8dUX/dAaDYAfR
445wu0YRGgo3JrUjRMc0W2qJMfFigYyfZc6kyDiRI4dY6JgI8oZDSPHVVGMh96hYCbAlCnIj2OJb
o2CHqyZl+pt1LRZmO4Js/EzMcYJAV3dltwK9RezmPGQyKq2JtcvcuhXgKF0DlFgdBv3vpjHxtLyK
P3ZShPyGpgUMlIWtzgWqZnMsn3pTroks5EjfzYrHbXDHVqHndor2S6vCm5m+1/OvJO6tLBZIl38Q
DTp29oQZdJg2nHwpMhT//tTeVrxkUo5L45LJeE5XM7rJ79b7gzSJFaGwcXuT56J1zijX5OH/VQcO
uxeSImcTk40HBYj88bdpR14J2mVyMz+V7I4bRj9JfINAGhI0b1aPYvuNuzqpaaTNkM6iEqpY0mx1
swxxaohPXpfIq3UDV2YEx/GDHPtaYBn+ww5Q6JiCuH+JE1IBRKUh2beIygiF+WtS5VTWBXstf3sc
XL4e9UbOcIiBTXyvkaHZEibdGbVpXIabDu74EONVm7yf943wI07dGLKmYBtQZOPP7WeIh9q2mClZ
NjR7r9qz6yzRSQ6o5AOSPr97s94cE+IPUypU9/DWz6rz3T3BsAs93PczAVke7xwi71FMk0iGmh+b
9BKS+ndXYF3zPISRz3/OohfYMJlLfg0KdCD9EnoYo/O8TeMZYE1xREMwFxGxNUkcmNyfDx5tlWCn
Kdwe507H2LLVA/mL3YmpXyIGGrii9OUilQCKAL+azG/QeXLLUsEAu0e85LN3dJyrnwqAidtM9tAd
J7n4kmytOtKg6BcDlNYup311iUhqQxj3suQM/JOWoiEqstIELyLzOFfvH9b1L1g6qTxOOLkY+zux
uikLr854ELH7wKBdcjUZEu37BbEsyeRiUMP22afg0wWU+cyugPBj2sq81EyXg3yeuoCaZcmDwfDu
NSFzIVmsQaYlOwnB8P83P7aT9E53x77iWMQtHyeVmtUt8epLBi3IlPWCQtpzhOpbd2sZbUzUQduA
DS6/4F43iJ31qLnOObib0Am8jYGBMOEsMdlMaujRPPzGfXZ8HHMx/iL4hDMBs9L7iXch9iKdkZUx
5YsWLxNmdWlkryr3a47Xpn2deMVRuOrX4MuCUOZXGuCCHKPcjSw05RKF6V06ukJXYu0iXLwli8d+
08W1qfxSFrdQrNAGbFx9y7lSnhfSm/OjAf1lA5cdC0fP5kK5CzPwkzVWKFnxuoz0BTRLj4ue8xpE
2LSeLq0nFLywyvSJIfj6dD+0nkRcfj2/V9uXPK9UoPk8qXcYqO8F4xMyxJ3fNQQjq13xRImjNTzU
KUgr2bbXBc9Rt3G5BWYoyAKMeSRTbt4jC5bzKpMXu74+rrscAHlAEd/LZR3hilHtz8wVNOxPPxul
rKuVd22GSHs2p6V4yvjX/8BLhITyEdYLZ4LBb7XH3qTURkAUdnS4dTrfnGPm6k2Vejgc3uW9nvSd
ArZjFLKTy9X8kvVQF9lJMd5kbDfVRrEwc26V62GuwIDE0+T6LEvKxpYH1SrLzI/WwDsdo2rRyHUT
Ipv612Csia1qzANPxMmrQo9Un25dmTMTYPyYE2Oragk+E9b4N070QDGwn8XFo2CGKSxDY+DGjFYh
3bux5yxcU7ySqgbntIgggsRHlSp2DkfEM0KHdjqAqsBi2Lo6Cmh49FTA0DxPKRGJ5/Ce4kJ+hf87
DSCrkzTaky1lg9EMa7YMmNFL9Y33bkOAo6wwe3AeQwMayiiK/KPTAE87szv/imWH+AN5VVGt0xEP
Voa9JzQVSFF8aFcLQiVHWRhf2TaH3VzyRT0BtaYhj/n/kU5PJtn8flQCt/d8/U2/S39p+Z92iS0T
TkeA/DdFpGpR5HTTOO3CYAc3Ga9FEMMSWWntzK0tw+uXXDuw3Q60ySy6oFs3cTQLypkfUTuaxJRe
BMsC2SQrgjmjR7DKDORHrheRFgBUNJO5W0AZz1mwmVxCS2uirV/htxQMpm34RBemsvI6RLOF5dtk
ksP5DxuhJb24GFV16Y//vtmW2HuBtgPfZOhxnrgZrfRRdMd/9Nr2a2NOO06Vzaly6U1fbTNguTro
PvE9drLuSySh6kTX8dxPDAiX+nvy8IDIqWOVlSJwMOA7DRn967hTvRDc7rXchom0lZRYOIWsW75j
hN9pEVczIPz1Jitux27x+zME0DiCDSr2/n8ez0W/1r/y4cp+rM9iiJs0qorEh0B5WQ0npBJKu149
htYfMsSESKuswRHdBwU/ak8v1qQInPhSqLWzbi6ayY0QyrYQtz5hI+/aBz9blQ4LisQv+kygRQ5g
3k6ebwRoknr37P+XP9L+6GyMdcOMPz2RdW2DSYGxb0iZHQJm65rbgmvf34jg4uwd9qPKlBd0ciYf
7xBNwBMrRFtPzOsewbGNvPlpjo4N7b4KIVDh3HlZCDoSIab5OspYXb8nS+FH0BItsdQgtwjUenLf
Je0YFalnSCg9AxCit6IUDtIl3PzKKx669J+TD8uGJHJQ3qzbOYpeqT+ssp+qHmpIwtf+xJ9V6zB2
x7y4rEymOFNly3B5t68JwrLj6DyvWwJ936tqdv6ZQsFK3QxQ5NYDy4uYWtk5XKD6GdTyq9LmGfyl
67jndU2otY0ReijgjoJYoDs58AuBCHgJL1ua6z9rC2sxtEpqjxieZRw+N+mr78dI8K2Hn0CzGlP0
ku5b/gCihRllICpr0kD6kSUUnQ9HCXpHEtkf7LVuz3kiauMsi0afAqDF3h7OJFPa2ICmBBlP2ZH+
Z2Nkd1tYvxh7D9EIulhSiDgbz/GAg/4LusMu7sKD/KwkmdUZQSp5IVij7Gzn4w3COk22IydcM+W2
JQsCc0ZjY9BBOJYC4Gs9XszRcYAuo95seObS8QYynKM+lD6o3MuRrmJzD5+RNIYUfgeIEIECl0YN
FqoIz9O2dYa3OlAlc4cWFWOlgh0hSAgRNhLQOXdf+bbdiZBtiLyt4bDAczzxJ3i2/1Up3e+rvG+S
IEeh7wiQ2nBaHDBsj3qb9N1P3nZj8MR+XEzUUtg6FHYDUYUUhx/c37waXWL9iCWonOdsEs+rs0n1
anbgVvWVzzZJBSPHgm38n/mzkXCU2J81OYk7/geeHbB8reFlmsHE2T8bZDsVV6878izoHbwPm7/d
CrUE0GqQJ7A53IDucv5U2gMjeHrmegXNHszTHid966DLHsS4Vm0UzzQSSfAHxWZMrdoPC7vUx6mp
5h7EW8JClsrBf7OHlGkhYasoEbuDy3k0xTFxjJ4Cl0zC4f+RJOfdSIl/Lg3hoKOevRhyCDRq/BtM
WRG96xe8cyBgtcp2SrbY7D+SVOkubuWJR3+3QtBjvDMW6E9/JVDm3DWXWdn3IndujcXqjaHE+bad
2VxbznfSS9r6iqPTtv2UzUGgW9VGZacebcinE1oRhVNwShcebmpAQYJRIG30GxtjkUPck9qT/deE
JbGR2Ku19qhoMybA/0xUzi9j2HcHvMlLxYHL0/oTXATWUaUlDsBjTN3sLdu6vAh6hvTk8tfYThYc
3sg1ODQLQiMCHKtFIVT7JckPaHvMirHVn45w/tIpkEb1xvEHPxvq4BXQILpYU04eKs29sVFr9hzy
5OdaCDmIEYMdEnFd4oR4mq+epkZwwERrK/PO+waS+RXk63FC4K3FgYi2IeKkvoAXMn1/arGDXigf
3YL2v5iy5QldMY2YvTa5m+/m0MqxcG9MlO2NRFIZ7NJ4W0Gd2CqhKw5BExMVboZ3msayoTn9EjnQ
R2st+l/Br3zO+kxYcFKZAF825RpeXtE9JSCIzsYoXnwptcU7LOqm//oqBUODp/znwsLL5LbdWAvx
rXbp9DXVKh7kMRWHL39wLBQHPLG+PlxYb/dryUniauxvoH8fQ3Wre7F/7umSTcbc+TBWwiLqQiPv
KyVlbMutsok268En5z2N9RrvQFkQ0it/IFDy0FPSRWKzzTT/NGo7bnILGamHlNT/4TEM188ulkGT
Z1PxHy1taDkvDwBN/V2k3PNzRAhpVN+j1ETapVcq4E6Gi1ZyyAF+v+dpLfXfOpvvaXryVJujHqNI
w8CaK14LARA4N600UuZxDLKDlpxkxYLjQdEHQ6GVUJG2GRGwts1v5aGYzSPBPncgcoaXWiRfX+qh
IaVzy8oNnb3Zel4FdghgAXrJsy7hH14rUM4C90qppSoGCps+UtmjCZ0RcrX5XHibotxmccxk7zEn
Lqe/fV4N2D/HMm0m03AAXg0BLdPez4PTMh76FbCX7zcuEYO9rNeQ9tQNUBjKLZCcKezmsZ1dhrAX
G0T7D9oLiRyTPAIjgv+8PtBmp2fhBg/uLpoHgp8k4EvVhzT2CZwnZq5zUnGHj6QKI317oSqQ4XHa
d5xlz9XnU+HuooMZco5qUJkI3JqfNh+ZwPlZtX27m7QmovPWIggndo5mRNmDuiruo13MZtJ01gNE
bkaXfBVFCeRZlsA1RDd6hBv9G6PqSS/RlVQ3LXSzeon9pRVui0bsJBWv9K3gqEGL6pBfjYt/PgaP
KDoJ3kc4pHzRHZZxofdgnhmkIqlL7qbE/6tQb/nF5UCUEtSV16N5ap+FZSu1wHKPzFn6tlXJQaVg
0OCgqOm1unah4snUzDd+Z+a0KOGjKViSBqB0YrOKMPyh/PRa7w3Ne3LhR1vqED1SeQMUroIlziYm
aPYLhTQbP0DYOlbzTLySbMXzCS7nUHhXiYdUlEV3VFKAhfXV5LkB7XT1l9F+WRPSssjWty0D1zVC
T9Sk9G5e2ZFtti8Sly7D1oGzEcowWyLfNF0AJVDS6XIpPiU/vAT6HFzVowAeddBxB5eWAZkeTTin
94+zC0XWApEYNxg9AHmaPmAJbL6thP7SacFjAgSUm0k+6ZAahr3AVleM5WugOwDXUuzfOiSR/h3d
E7pSUdsx0l1uVmRdY5gR/CmzGARx5aopQYVJVEnuOrFtJTBy8qzjMC/Xj4P2x/zLTkjkDOf3sARL
oGO9sq5YkFjuAaBaUdcTtdLRiye2I7d7YSYIfknrUq/L9h2HpqpcA/7rOAIr+i8LIyQkmRENMA7r
Y+hFcaF+cBPSYPWyneplsaaj9jC4AoBrTTTo4Z2oEKrq+UxOOgIzO0+HshkYinVDu1BTWJuIoK6V
gu6EKxAO4naCOjdjYRtgZZBccvuIeVVftt4VzSIFrtWrDlyjPFOuRb4eVTBDI2EZ9FW/H9MFmS/w
oL8tLRP2B/oaQr2VzhP2TfJjjdTlhQFivOFldgLMxF4gQ9PmbkC83GbPOY/n4r86vOFUwxxuugmB
HPl1j3q4Hxh9SehhAEjNV95FeqSgNN5MBxy7URi4/VmHgwve9tsT0i66qydkhAUH35iFbcI7eJl5
7yu8sYwN3hDqSside7jtE1dctr+BzmEYjrX485JtjDu9d8hpEXAi5Ed34PDnjW7MVh0qZ/DgacRX
JOuwI9tki1vvwFdPDpMlttsYavleB3yLHo7AG2foTKMnA4QQjQtups5xLFSbrXxSSYGKbaTpfVy6
KEShPXNtRrXD1pJdxwVjb/430XY8jR0A43+pU0hr9z/XKOOcFUnSNBe+t6EXQZqOIr+cd2Wj3mYY
ootOdOGcxiRcN0oDdUb6JpQy4LaS2gJgsHztx4oHBQQwTcJoAk1Y0YZOoKpqZ0L4ahOHy165dwuX
z6OXcsiP1p0cf+SYwLgkBlIttH+FLdpfw3hlPX3FgtkOuLEcO3IEGowbbJNSyY5e1oqrXBrMLndQ
N/NZZ/bUa/PIxoTKBaan6WzOQ2gJDaLUy/J9r3iHJQMTUfw6PzpudbzTRmYyCcEa2KjI5aUBsqj8
z+nPmeXtvCSESp5skuVXpp/NoP7xwwj/Pp9HN+o0tMGRBZWgn3uQuoTd1eC+BAFsS/KkZnx4I7Kz
ImqHiuzylZjpPjGpJaYptfjSG0i79Y1RUyyH2YWASXZWrAuJMim73qU+2xl5R7uVK56u+5pJgpQD
umWMX/p8Jhahg3e1VHbKqFdNDKyBV3GU/SZw5uVw7QdhB37mG70mnP++beq30I553DQ7vrDoAzYg
pzbxHqiQo0YTRNuVnCB3/D2+qUgde0Ow19yY1EBYNDs7+XqqCbRuEieBBr6xR1ykOWji8bGcM2TZ
W+BBjdwFMWVxuY0eMed85FkZ68CMMrhD/NERbtNtUowq8YmqPImDR6HlbKnKtem49bFkQk8X43mC
y0euFAg9zGfcVK7J89aw2hgIVmHlTWgIEc1uIVAAjgECjkPOFUaVWOboJw8KIFAxPYiEdEQMB6XY
Jn69V9VZMAEa25eOiXzdMiBiQZFu6GOpoIfw++GYjF64z6e6JRk0fU+s8XZezUAPdqm1oMSk2eee
MaRa9CerOExyOOq5eZup3PLRlb12xQ/XwJp8q5ioNsNWIXaV4Fdmsmbs9afuzr8t9WS8uea9eR/b
ZB13HJXyfIlXn/8B+XqDCMCrSOmizLD+mrkSUTqSsxcBeWCqU/pSO0iJSsjnIVoTADicgrcj+6vo
xFRPE2COUm5fgdsqOXR2CEDLd38rPFIR3rYYTAhxCaom9+So8m3suds2lICckSV0hcGMqoVbC3Mv
3C/d/KcXeRRtJNvBXF8tzYNX1iPry1G7QDqR6l8WOmjkfkIvIu6Z9H0+JQiySn/gyprHZsF3f1yA
wtHdiK00p/tl7XEuuYj8PRrueNrDf0016iadxWL1NDgIwMuUK3vJQ69rfGxrC6zBvJtBRIZvdTqg
pWY/ob6Q8UuQsllb2caQxgsW/TONkXWsu34fHX77P9BctHbhuIgn1tWxCrLRcpdH74OjnzZEzMmZ
7vYyO5jzN/kf3sAjtTLhmoMF7hTwXA3YjA9gpN4OhSyAvk2Xuxs/1joX3mjCLYHauIGqcuQSAVTL
FzCDv66h0GJyLisP6Enq1fHdcvLCdsJWvkspWN/4CHKpQ7Za4iqntQy1CuH7ZgoHpMWwpFCrqK9E
S/+SjUMW42G35oqSkuItYcDBa519t5nqDmXM9n7DTtFlU0ykvyx7yXMtj3xTkXZX4HwUuLRL46wf
VdZNk2uhDHLO3u5updeQkDRRHfpXu7XmPdI3jUVeQ8omBunBuKWxa3xhmTb4Oj77YhjVlTWNaWhZ
bvf5S0noX5fXoPOdtl2gaeTLARNxaZNRg4EqDlqBsWvaX5OEhFYaTmvqqtSTxwp3UDigJcCqfmP9
v84DVOWG8c0QlHVeB2E782oWlkdfw2GOemyzoVNZFAA6vvdTOdRf2DageTl4dvIKQy0mchbXhmQI
w1OqejLUCFG7jHZsxm0qVufoBz2zavTnwwOmVJHmjfUMvpvYJUnlB8Hf1ca6xk7hBdEtDx53woq8
szj/DqEshOlRzhNTXg26AENy/fFdRF1FzDS3vWSNFUuiCT9Rk8E45TMn6dIg3cjyZo13Lectk3W7
MR0r4dWtV7sNtRDYF2LEw4N4Z0eosMHkFrTZm1DIQYIoAww5fftO3ZSo80DGnjQRTwmBsDbJX/XB
wnL6T0192bs6jpdTfs9CeXti6lk1ZmDe1DowNFee//mSAIAI8M+vy0pmsl3Z1kRQPO1P2r8vqAxI
6SZclZ6yCGulkveZblwuf/7DnJjWduKZlB6c3b4p3PxLmu/8NCFNMbbzPD75NciRFWxUhcFExtYb
ie3m0R6hPvAu/jl25WfeUqJj6IudtVD2DfF3nD4eoQY0YTdTPm9J7xBe0HkQTBJqE+mQXgcCrMqX
tewDNo51uY67w91taNNSo68pFFVC1sCqSoIdvmKMzpuEvNMbMZNrU/GnxpImpQ8rwekYlJRXqq/H
5YZzMFzjakmfkEqEH07sYVq6SKAfSDDtX9hcwkXxAhsft7R4LcfwBEg9hYVuVaVUrcyWnipqfrGo
K1cuKBvmUXQ8e50c2LRBqs2EMF/vWSUPnR1Xxp0W+vxJIs2JBiG+gIgOtJrfNUk2PnmtxT0NzeHc
M7zGcA/yyNrgUjO8UbTjiNKEHtVmTvMrf1u8tG8+MijvJwUBSqqYKvRc3YkELPgEi0NVN/mvDSko
ItovOviHLQtm44le5aI50LSY8fnLj1SeeIlaexw7XUE8Gwj/SyAqT+Z8tzvtGDDXcDczSwDDs3A1
KOltcqapXSinvGO76/x8PNg7rWlc1ftfN5d6Ol+vNoDODnzo8pwyFFBg6XYBSC+FOFCocFO+5uhb
d7wdstSijVAJ8QDCsVp0LzS6nbMKJo/5TGtHC6pyA3xqB2r+SmGnMRhaoyuL8493ekupmi6mCcwF
zte4+6SvLtkLhDm7AqJeGGiNIwMuFfPh1xF0Tgs+frlViHkzhPavwm9tzhWNlUFoDFhuUlfXEKYw
YFOzEr/KHU97WmQXp4r16tk5MHUdEt4TSWNPtCLylHmn6sG6HMrwLLktJA9OUHZXVvCiRHrh530g
xyUgNhwzMdvwXAhNnZdz2+8AQUEt7ClgBsV8qAI4M7TDrbgaLk8nMFie3c7ufHEwQ6ujv0YRA9TB
DM5KGLgOlwl0ac82X57/pOcbC2zvx7IvXTV/Zaph6ye1pky8+mvb2L4QsrsZAkHkUiBI36xMV9lk
xS/QPBJfEIm6+xOmnyoaV4Adzob6mDhMKlT/+B5837fX15iKPGnm1ngcyQyQcvQin8dhZSdeuGo3
R/X4XM+4nt+IMRYnA1x/r7X6UMbQ0qxjRlqfdlwTmwLHcV66nIQxCOc2LBj4i4KJ/Y5ONJKZ8OjA
vmT8NjUxsY8XDLuzDbBxnYiW7BNhP3yiI0wv/M7fExrsqymW0Z3V1NK4uBQ4xusR99ng/0X/hh3z
Q4zAv5wfLY4D+NSfoVz+ichMhc2YVKlkiPFYq66dhyUcufZHcrPeEu8i3ujpsAlcUOJ6/LLfS5Mc
tRVWM7YpTaogJJph+WiV544MGdRHYMbMo+mhm6TgWopW3poFohNWcVfKHESwWFI+OslP4F++8tjM
UaMNpynT70ySIOpBb2WBnAXWD6LjuqnbpQmm71J64aP9rL4fKnHClyA1ROzt256QiK+JCItBsdg3
5W36UZ7LdqmRMrSeG/cJJJP8R72+f8VX4Dvhm0hIVF4K8xSSLCwGfg7VYcPzm56BFvaLgtYwroIW
1gpsQ12wzCnybGU4I04HPTmWLSaTaYqJy+bgcvoHvxlOG1xyzBpaAsOX5C5JdT1gUeVANxa63Rlx
PE/RonQ6CFUxAGQgKZPC0gK3nS2j2Ttdpx/zTAe7JRdjXazNZde6s6hUtvTpbV7244by2gkmG8CY
NLe46/gjcxvSWgIr8bVlik9A7QStY+ByO0U8/CSSi4ZSxXFXciNsDlwVPXjBvOpEJ5GEjr0FewRs
vXqEs/rstayUZC5QanMHYPbZX7KV25hjiQkd0K2i8Ox3Oa8tJ/lKUUVQa5GeY3rDBvBnEMz9FeDL
Tl/3AezgAop0HFgT9s4hb4oE3NlufiP2+juBNPAQ7pLfBy3w7puubd+dxQRivF0iErv3709wQ+Xl
sPD24XBtZsNFNNOrhkFdmj1b2VO/2Vu2SKEU39xvz59GQkak0w2pUpYhjo78XkKi1tnx1xWd/m6q
NmT0xqAoqKYaXEGT3iy8urFSNvJrnSXgqYR6s5Q9bPEqnc237oU9i9ZC3wxHtsC66qJ8JObW4hAT
z8dKzjo+hMRilDr05vFWHUS7xA5eo3Wt5opEYBR2KYXT/euG5tKw/53mDnT2DXz34Jl0fJcq/ZTC
mNg7mOr3/cKErb+RNFOCiijgo0/rXtHkNWd5FKoGC0so8nz1Jhh86WNJPLaEHjApuknUzbq1r2UB
D538/YmgaLE/XnV5TLEZJauy3RNelclUPrFKd9S7skfFeFFu9pSryRb33ZMJKA3j/C383veGVA0A
lOb5fCTfBJMgaoxqZJTG9+R7KpH+B0Apc1z86L2Gff/jQvIiiwxRaLZM03SlcXJdBhI+OhrbHHea
G8Fqe9c7So8CVe9jE8NeRjYbSAp0hvwVWq1U3tng74sUqmWPFRlR4NC9dDgWh4t0d4VGMHU/mvbe
HMcXzAEdqQ9MNtH7tbdaSrHU9jPqIBrZHBNZYaoN7pbyRubignXaaybe2pcsz3PZBNDrcpXMxb3v
lg+LaAKDClfzWgjiBnwrMnu7wIaBnQ+YVc5+yW5q5kBRUm4Pwep9zvTK/ssqPqVQ9fTArDfr34Cj
Ywjds9jOMfziE9ZNqkc3wS5z5F/RUgJ3gmYlkgPnuivKe9bTwHPw10PSUQPypRqP/QYkiP8PgpDE
4Q1gVi6tAGKUk+ZT5E0lNLUStHHhm7t9J1rWK0vyXemfitiiOwkln+2ydoZA8MrI5s06V1oAxptz
oq0bBxfj6otLHudgBO/avKXj6+6LknaCIJtZKkw0Kp5c7SrxreaOIwazmFOOYvtCMkb7cPNm06l6
CfQt2UsAwbKAxqkOrL6MeCcAJ7R/ohsaCs3k9Tig9sfau22qpLLDy/AvXvC6fNKhVPXJJzegIiMg
65T39mWImh66qffFW98AU1vW+50o8UXX9Yr9B8p1sVpT39RQXtuM+kw3iSjdUMyvBtNk9x7PMGtC
fcNl6mP47o9Ipgbg6BfbD8Qukh3etCEMbGeGcMjrpqiP/T9N2MNEFPgWaBp49NSviazzVrDpNAIg
X+hsxVB/Ak2PLDUOCtJAY0pmSkTEVxSK5uzPWyKhGEKebFeodtobS0/sTP6J4HVHcXNnQtHeq07P
M8BAxgKgP6Ha2YTRKxBOlAikuJoAWdhfA3PhoAosoXFCted4F9Q7Ip9NjngXGzNxODrBO9xBDVBu
G/hoRtVhMw8+7sOyZ6WMIiQfYXyIKJzLprVrWIQ9eAKgFjkon2t7AyUwoKBg5pw6CUU5FuZbXhrv
DvTZoyrZDBNclCW6sgWZQdhHcfmygTvPXj1rSuqJ9e8dsd359gH3/MnRMrHvE9bkcyANuVRPhAAy
cc4NXTPsGJTAhU7UBsjZLnznQVUxJHy3tXec2D491J5Jby11UB4g0nGxCVcbF+lQ/wsxqa0yPmE9
DUJmK95f+38koTUpsdY1rMQXwH/5BI1E22xrdMYQxXJ9uzVtrsblOc92DQds+a9dHQRQBgGW0L0y
S8nhJlyE/EchuAA8e+cPHJxEKutbLeDkH2hVIQPe3Dhj7sTIvx5FCFJSDg0tdovRmyvHMByZxFZu
EcRdrtL95sr0vtf3ljmNq+7mTxw0m69gAhfp/c8PMNHDTPA8SLy0O+Olrm6ZwtpHk0B/cN5A5BNI
XCk0qpKG5Gm/EJB5S1jXdoq0GLPfdSrrbB9hN4uV1bD8yJDsEyvUZCMrCXghE/z1Y3Xlc7in4ao2
3y5x0dUUm5jNyMt1EH465kLR7Fal9eW9cmBENGKmbcb/asJ2rlwSLYndsScLcMsKN+EF5imkwZM0
XZK3FmoQ4n7K+xCVAXcdamp9y5bAq9nrWwrknbJO6UYwTJ53u+OXIAraWQCuNT4Xry01cP4CtafQ
xZ3K2KQYFDFtdQR/0W0KUv/PJf4n0NER4YkIn8QjX/y8eJx90P8XMkrhK5ehQ85AOGRD7y+RDvB4
nl2a+JSa6ktzijoGzEdibbTU9A4EwVwaxlPwxuouX/iaAEuEKrcKPKY0IiYtK25OT95v9tC6AWX+
7+VIIjIIMf+SjT0xxFXqLGWROydJ/0SqFzUm6rh5GFx+VtW+rxNkFHMAVjDSZugQMw4EAkhM28EP
pLMw/2OsnJeV+vQ0OTGaTP+boMXC1a4+wsJT/8EBmOFVt7K4dQQ2e5FUbvU/99ewM7ETo+WC7UY1
qFTpwK7ny9Ciqq3nsm5sR7hskX0INT+U/Tzxx7QtYeHlo8SZ1B4x3s2azAI0zt+vKyuCKbU93oN3
BFDH1Hy17qHMmyxGOiA3TbS+0WX3nLe70jqCxDKV32FwLbjdVJIsqODTxC7EnBxAXE/T+5GEMueb
R5oXy3mFhoyIlq6qkrTGoNyLzWdrooj6yIegAxT7XjrNBk5wUh0h5mR4DmQpi3HLV1gtVKIYSe9E
Y2heZscdoxkWeQ3y7V444ux2Qe/IBbtOJX5ielEMh/tXUHEe6ZTdjrE0lLrOM82RBMYkeW3wKnUg
tAGJ8PJzGeeWDIWA/opbbWQEa3jVOuudAj2YCpWUVKMSRn7JB+jnrHnTu2yPcYOdsc12JtIyqbj4
mnTIQadeqZvOv09mGjPHUxLVIms+5zL2Js58HnHK9/gfbNxnX/HNN1QXfAWkF8UsRYGHZEvRReK/
fhl/4HI+ggM9pb1sPldrVDanc0JucCvBgz+3PNyo3XzFAjvl5EtH3VR00MzTp0rq+A5PbAWaHU1A
FXtm9Wlr56wA0Cj+mbFpgBjzukocRcItQFAG4SR/9FOvX1dUw3JTKW+3+ltA3rzmHnLn/mwXruWA
570/dMmFPz4bLpYhbAUigdYxUkZoUiGN9qAXhClM2VJ8oT9PysW0Cfk0ccyW4JnQvC1FxroEO4eJ
vr5zCB4/Y+/LSi2Me4G8ZlgGov6IRefMUoQhgYJQ4Xf4zvKM5aSGXr99iZfw0nuvnCmMvRpSU6+c
pANw8IRbPARkSJMghyHrZNC9xnLJTJeiBTmz+r/x95RpxWrTDQJkumnXqX8d6NHgT6Qd5lODWOr8
q3OBcRMe39o0Uyxnrs71nbH/ePCuuwybC0Tkpn8DfIb2PW+TpW4qxhOXDCBW727Ignk0vbxUfqV4
l0EPC890BwdVbGTUIp3kzEiAyID+1fo9Pc9WIA8yzH/OGuDE4U7Fm6sqmP9qvVxr/3NjxzO13v7k
mH/ggSeCONjCEVRVt66yWUi08yIl8aV2Is9UH41EaO/XRBf7WiZ3FF0W+XmYHSRNWSMI4SW4OcDG
PxCNl9zjJ2MvvcAGahFCpu9gQ7EXxH6Xevw4u3pyrpdy1Kp02Rza9MQff7Qso3Gyuk6bjJxtYZxF
sTXLyYVTuMAMv9EmJ5NilCWjIn2ASbN3YoHnJ7YIYmH+1UVLvGx+VJ90Y+uoyYzBUUTGvW54mWFR
BDvZA/zOBrOpmaMmKcNn5TxirA+5fN3g94UzKKZDNQFqMdN/vP1lVwNbdc7wFB9WhmKthypla+Qp
ALfJWgXPBytXngMBjXyvmWkCcui3Bg4dDH9m2n8w8b5VTfJfI+MP8GOGC17sZKq6ocvGcyo5eO6y
0/rdX+5EltlQs0YAl3nxVHju2RL8++1H54Gt6lE1qfhecgXSrJjm/vdZ9mZj91qKiZNFcA8+lA37
5xLI3WK7qiAWfnQ3+W3jknMTKjsS0weDQ1Viyj1CcKjUmLyRlPeE8w1fHqZp1NrWNrrBT/3Midwl
vhl9tTOalc8EIZHAJ5TfynjGWiwS4my2uywve/z1g23HefwcfFAG9ATCdKa+6Ot3O2IQUB46zj16
JyVEtT28cU8aYbrs4xZvDoHkLE8FA9cHRJj9/T03QI/rWFdMSqWGbGGFpNOhr0NU/cFLgRClwIVl
aYO/ryZqytfenCXZYvujm8QabBYOvJ807uWo79kdnq/qCMXSANX5KeijEyScrUi9EyGu4uXADVMs
fWJQwqvc4Qw91s3la6o42tylYYIWTZUclqFqIfTGnGVvzFeOEy4dkcl3QbAetzegXXbY3X0JeuUv
hRHUUogcwEBYf1SJhkIZ9jEmeeloeKpWhRh/pxelJgF3+p644jPZAfYlD0UWNl0GFZAUeX8tfxZR
t42LerLacI7qG8zcmg+A747H42A6wyN82MsGIj7YId4eJfWq4SFtdF8UtByYCdYcEURe5xyC6AXp
ZDniAPue222GP9CmUW8dBI7K+cLLldR3NHCyR8uHC9L+Rt50NtUBGJDgCrL2CSf7BmN1W9fpl7rh
alcd9CEXmc9LWyjW4MPRJILvlMBlMTVoWkppVMUeytUruVHOBa2eOQubZwgSpbj65Tff8GnOd/Qr
9CQwry5Z+qyFE7uswrmcP/YD4tSeh5QW8++0wscQVirvP/VsnQc3CO5M3Hq2I7k6/R/OovvNwGXR
A3Vuvn/tMZVorffTcCnF7tunF1aX7qF7zl+bo/Cp0Om3r2UODpfh1CL9BrwJObYi7svBMzN0GZUI
s8HwgyE8iPCkuqDBA+G408mPFwyNUP+vkmbAg8DvlvCKQ6OG/d2hpoPr7Dg0gs3Z8/JdrqvbkSFl
pHb2dKXyVYM7cZ7RwzVE0p/orftKwCUPItYxTvgEp+DB/qTfC5MiVljKl1vdE7AOf29cJCH45cyh
kDsCpgpjoxUV/4hSyiFrlHlYUC4DgUajVgalx4Ddx6p6l6UywQFdTC089jOB3JStRlvUU0vuuGfx
qHuxa1Okteb0jm7w6GmcRivM65Tf0OslOe1CNzDwSi+pFmU9foCZfIuIN0TG+fGFyeNPQWp1h7/L
QN1QEe1V4b7BwSbcwIFkuOV6rjC0WVjq9rADEmZJhwmEXL+BM+NoZuAYvyV4qj4jeH/PLd3BGMMY
nvHHEhnsmd3QsrYh5rHaFOqN7BfI3fn7l0si/43NLTIVcJmGmud7AXwl4RKLX+dLgqSURUNuQT+9
wDmDE7FV8zzmObK04jAvSKVrPF1mAyJJ2TforYQVrVFjIZgnzoU/DoRjNRvSfU1+Ejc7CwtIB6E2
1WJLqH6ZKfwnNv9++J2yeDb2lw5v0TIdx+O4kQp/2gAikMeUlXbQXWjw58hHZhX7fOC5Zw5FkRn1
9aP6f8/IpuWFUTImlAM3zgpInugZnXPTW5NX0W+tg0LIvFDeGvqz8vznon+c0P6kdRAyk7D78g6Z
bJUAZQqL6JWTCqLOSbKrujMDBAohCRgoF0Lp+1UMjsBVk7FEpUMTRXO/BTG6AhHtXF9204Lo63Vh
wuKCW4x3o6h526Y36WWveyf5K6o1+PpHaEuBk3O8H8Xl3Ctrgm+jNPJPsH3XoMjtuov3sioa96SJ
qcGsm6IcTgpunzoCPnKcElCITxFm1+q09bfXpVhJ+Vi1mcd8I8uNpqEn7MQCkZEzk0vCcQwse3Qq
ZM4DI7vlmulkzNjSM5CMi+rt1Q4Fs717MzenxNOdnHJxJXcsVG9KQ2/HJHcRtio+IJfL4rjOWJdC
44wFSf7eZ96fWj0l4bqsPCGVTJGUr/CA+4mEyGqbKYyPWNLSBKIMMhAWJJSfGBvaXBT1fPnaE3om
Dgx6BGGfrIkUDYfzeSfjKXanONgXUMZW04RLEpbmYzzj51yFtcYF3B0k2AwrHcmkt9GNxiFwDwGU
qFk3eh/59iQVgHa5BAwRRpnVMpxTmKbI5luKxcFzcUWfqW8eX3j1mLYfCJJ0553cFI35B/oHOjng
s+i3ygowFlE+o5lgL/q/sJYiiSFt6uTx5eZtywAVBaKbMTsrNeXvo5T6C5Yl5/Mba2neM8MgF6tm
pZC8t0erHUjd1Qeq9F0yEz9da2oTgVlaM/QFxk+svCpK+7BCHziQdFinoa0tzj/s4AnYdwmpbF8M
TfUx+SyyyIvHtsHvozDaGou62fkiUrs04uJ76dzvc+uZX4i35hDNDjDfHVXochDSEO2NtR0daHvv
u9vVkT8iX8IQZNeS0a7+KoT5ACIQEeyM0//a/nBVlCoA6hsGhYInBIH7FFRrCa0npZFvf/pGfGWB
+ReAyhqLoKGXBqFt6nl0OQXmwBoV8WIvUU48bHC7qqRuboYf4EFrg08wFhaHUT+62ndr4SX//BKN
2pJ8iWjCZliAqTBD8qNhsqWsoY4yOzfJx95s+yJPSEGXZIKUpchVwF/5VcbVXIwNSsoN3zd+BmZq
7k086gl4nL8k4ctM9tIim8d0hiinBneVrFx+8t9wdeRyyI7BNtkAyGRYCQAOXTyNFWKlB4LE7dsJ
MlOh8F8GjcVe1JD/py6an55YGHGR80+INZflr0c8HJGGvmWx2o9QmtfRS6ihfg036SaNA0wRAPoj
VVZjyrQ3bEuFBkOMQBmyFXy8t1V7y1/lLoApXIiz03I+Cca8hE/i3Wv86h+86suGNjUZv91QWgP7
8Y7J7d3O04MUBevbtlR/xYVcGONOSBuJ/9+5ClQXnQvnJ/sDONeGFMRlijacVnctDwdEGfTcXfaP
OZ+lz0DEYvpYv9bD91Zx1KeHPDa5RSOjEQ+wUipnRy8wbI4jADpbmYHR7yNYVOfubcFHW/rU1gdR
8NmtveM/gkv3iay8fddxFhBAs4yxO43R9qXpWaiadOOIKwHcZEifQcsnUw4M5J3eXwHRC419ece5
BxheG54TMN2eAwQOIZ4lJRzp3cHydqxFwe5/rSJS2XnVkFuNywWEMQqQzzNcruG7Fqfw0Ot0hDMI
x/jGQ6WgNALznc3xho8jHPOklzzvhmZiDxkk5bFbsl28dhYlwEMUMhu68ipNi7aaifHLwFkPha3F
4BR+7asr/3VNcMB7HIoTdI38txW0PT/MpWH90zREzFIYe3WAMcFy1ajvqwWzaMl6/KlK+Q3zU+ZU
S0WUo1wkAc8fihYn3jJwSnF6GisHp7uC9iDPvjvzliQhsLgEHekNsWR4BSoriR/5nATO78birqfl
blfBDIstGaOPHIyZiWHAzZEFpsLBY2nmA6rlJHo7tnh/k6bdaIZNY190FZsI/M3J5pDb4RNYaE/P
U0tMuIPvjaEKW6d9REGRgit/O7eH5Yv9Gm847w9aTj7B+yoWfIyDPLcKVd55e6L0+DbeUzgXD27S
jt3nk19y8UYLQluKc7BlC9B2gRxdGpdQ1DcLhM8oaJHAwjsFXXc8pZp3D1ls3W2Mn3Kb2kXOVd9z
QnyxWuCz6q/nQAkBkQtaNXSbsWAg/9HYFVu5mFte1I+nAr+Z4QU6tX6bDoTcEUTflHb8JPi37xD+
Srw8L971rGE+rOurTKNWTUjGAQfROFkKMZJSHOBmcBsy6acVAV0ZzF3Y/m/875Otodi9zxHQQkSK
MUNrf/d5efVCbhyIcN+UsDTxSR81Z87Vj43QF/FF/nj9sJIYWFhTtxwRjbRDTkzT31fxdcCaKJaK
oQv60lZrN9K2JaNrP8EFYyLfL4bgE5Obe1B0t1/xhmgmvL/GzQiAizKkD8AGsNpx/d8paQ9KOUWa
y3pspIdcsVgq6LKpMkIxQ8aW3QByiMf6fJK2zNV4JPloGfVX90QLx3oA6FyT0WAomQxbLI54/stm
kEFUnNapUL8wGlel6geTqBdP3lqslXjFMYmCq7lrlF3AY5R9NZ9BWyxV6WM+nIAlWbBkbQpi+edq
F0fJCYiKZ2eWDJw1Gx1A0J//VEtQSAoMpM745ku38mh+rt9/iT/aSqzFYCsDRdyTqFXnERWV8/7g
T4NtdQGNvRw/4yvfkm2rA0zX70hN9Htcv1VxMkNE7FAtdKfcLv6KsmJrWjkChCxEqUdwVKFJ3Vqm
cTGdyxCE+PqwpDXl7lufEwh5lVX2uLlQ7DbQQLINapccAmlgz55smNrKfg2Ze91aEs8c58blb00E
DnP66G4rqWT41m8ypEafojFo3/nvCY4gPoET9h2Ek868/GMArInW2G/SoxJeFyY0f2jsJdo6qrzC
+ChL2YaB3Ip0NNwMXjJsvAV56O2/ohNzbyZV1tFIsOs94DAJcU6SatyZfo6LRiIaEmXTuI+QNpSM
ztgoT30FN3P7abNiCdWHjuT1RvRZxDWk30kMaxJ8jrRyNW6p8IvR1iy/E9FK0waYWs2cloUCdYJa
jNgzl+h9VZo4zbTx4HzORwX5w3FS7hJke/+FYEPTOMP5jDn65lKeIdwJtg3bgt/92h34yPgee1X2
fVOb0LD0EFy+nC1f9NxCU+l+pG2eGvGQ4q/QtXzt5nfriziQk9QqTWihHqg4iY3WOLoZzrBq9ye1
/Ky4EG+NPEhq0+xJS7fMtweXACPkZEcw0kOks1uSw0LZR6P+OyJvzzScHhaLDzPt1/AmFM2rlx6k
znN7kNRMsWJvcRr81fMksEATVUbZk7pk8Py3YgezoaNDRhrIyg5NUuw0o5P5gk6tUKJpSsnE/o0t
8Je6Tlwyu3zc7malI95qQmlslBom2MVin7lwFiZV/eI5swlRKB+l2CIt1bui/nA3hxldEKqYeplS
mjFY90RQ6Dxrbq3zb3otNTCJvOZum7O2Vh7WpqLlv0yu2F8WsOgnqJvp99FexEhHAdeiAuZIE34+
7EjU/22/xiZ9hNg2S6jzOx+UB59rLM0Wu33TDfv/g9niDdZJbXF2ZlYuDP52/iSwnRvTsVp8K/OL
kiXYPwY+oPXHiCn8lb2l/xAIUuAWyta3wRP6Rjh1WgcyqsIciEDM8JReTwE2nN+Za9de1RCm8AfV
WYi6J/hPswuNReLv0beirV7H3w/9TB1NuKbuCKFNXhPeBDXb04NjjHZFEAPGrSXOBj0BhBn8tCKZ
7JUOgSzizfA/YB0175UcAcAkLpsRELe/3ku+6vhzYBThZBlLfLKxSUp7UAGGTJt85g74TWe5Qx/V
uB307aad+6Pz9PfCap2YsCFT3JBccPjoLy9yia9YFG54p9P7GzZjH47/nemM8kR6ChCLl0brHVH+
I28GkvCey0dEjQqjZI0RXOtB+0rSbSQITi//QzItmKVtwKwzHxfQ+L0msW0a+9W/ny9HMfzruUwP
50S+z/VXRX/Uryf7aMoFu4wpd9ZSVZIO7LK2fb0Noghtl8tFMAWHpSxq8VLoW7AjGSLJtgEKUGZN
N803Mxpn+4V0gVI/UtYPfm7npRNMoNak6eOQ1CUjL6zgvstOyhT9OfCLEdQeEM8EN3TlwPR8XnUF
jNszLqgvyYSam0Suq3Lyp7xSn/gMJq9xVlNJeRCJQUttaxC21u41MMOcbbtgn5GEnqyAUNP8wARt
feXAAwz+5wL5fhBYz/ZI+WSk9cKYF4Xf4VAZmNtnE3D7RH8Dljv/eIzuoIZAVf+NYwzmjUMg5br6
IfyxfibARd686cZJfw4DBV+knqb4fnWjHI9d9iWrt8XI9rGB4udmx4xgSZuFQw99SSe4DdkOpJqB
JfFqKUTVLZoBQCHiWzvwF2ZSNU4moqAtXe3ditlDkDECdEIksd6nR+zJixj4O4erzf2oW/zbf1Ke
1KG5z4guJRoJN9QxFpqcqPcqwCELJBC42kkHJXhFakkaiYpMQmNuoK/q97JhpC+kFhwkTSrEprjP
/oEztrFUOeEqDA10y5Ia0k3pAF8m/i4xCIjg+ZtVtSSzI1fqB5mK9724KwcHWZPOnewTaU30TqYs
ha0UmypMhqGpkwQwolD+1cWb/QeiCVBWt4raq+xx9hiIc3YX1/K/H07hGnfzIS1PRI28wBypThBC
lc4dXgDckK7Uts/glHDUvMudly4GKWUqrRlEpeyHf5QAar28+Kbe5KLQ8R+9fdcJGZd+thj+KBHM
xgcngoXj1L5b0No2R+HhRQjtzK9QGz4D9zf9ar2tkdFf9Row7hsySqVOkijVFGP66OtRUr5q2Ny5
7TjOAgIzMMaYo6KvvjOjdEMv1pNmr3bc3aXK1YF9w5YPYydjPnv8bAKeBLtR3ztSvhiPZd156EIi
YNCS1waOJ1B7Y3qP7KIqK7bWp9xoZxI1Hua/3FTSGnVofNWL+MGoRrAMmPC+sUrNgWDlPsPY5WiK
EEKVmxUZMO9smlyrDP3d0Z3avyZww7lYvD2dy0YZVYKOOZtvnF0oiEwFC4bMgjc0gwP7kFUDuEFQ
EFP902uzr8AGCJKkGd3bwyLZ9fCycDH9VEGtD3ydqy8vQZpZDqGbriEocbbzNaSH7sTDvoXNjHg+
1ift7Yz5WGfbihLOYxExNZ35tw0OnR95vNU0NWEeDnS+Q/g4wFxnJdmBjiA0kTMQcXRj1Xjq3D19
9HRV6KmvAaQ1ikM6pTAL3lDukyWWfYMQjCmsrIM+frQWRwI7AKTctknVh+BrfoRJel7iwDa+7dIA
uFezqA4vwM7gwLZodl6HvCPcB8PbusNFxXorPC5Rnrwb8wyt9Fg4l9R8cPOlF34wfi86OSWVPlim
igj/K9z077wT14byi3ErpRS06Dvjf+g80S0Mv7ZV+fwNkzKsVEE2r+OzJuyVuI4qlB+BbIiA/6/z
Z6+nwULawy3GtBprCq8IfSUFd4zqtndWAJ+DgMz9vq6LyVaZ421zY0Mjic9SOC4CZAvpGm9aGMR9
UkmBHBJMuN8gkWZkKE7QMtvesrfldhse43gkzcl+/iUW1Ad6mQSYvkBktptiOhQrNLNHnLkcaZdX
b3Mo5qkJvugJi3WKuo5ehvKTWEUw7SJ6USfO41HEH4D+Zn6uPj53weAX9zo89YaXv3onaBA2Otag
nWNzBDerqiyuuOclYZn1cYSfGPdVg88WYQQbZ/LcYvK3JMKTKaaWChCXLkd/plU+KEq8GCjCwa/Y
7Xb/V06v7G7INEK/7h7dDISF6kl3ARmE37OVdnSWEDCzlngLi6xAVEzU05TuT+0pwcX2tZlSVnAt
Ef9/bl3PRmAuz2vrNXt/sI2iZNJtT/K+nkLAyvYpl3tdMINQR60ma7kUwCi4g2kOayrVxmKJ6rOn
v+sJbn4BR3QcXsjYVeq/CiMub6T26h8jvb1mqXCzlGpfn+vbmJZjYzMxRWydrf4GG+I3zReRpvVO
pyazZygUGVZXcEe3NakDCRyChlcZAs4hJgz0kghKYHkKV5lqlsVXH0PcR4VAebGiTu9D/Bb92iZe
K2dgu84cG+PMDmDQ5aE6LqWTZVMYM9OFhsXq8/pG8V0sTnvvQbQGwXN9FGrDYKI81Oo7SbRm7U8V
cO6QGCGxbkWxUiy2U9D8h5XTpnMNTBZpqNn/JBrcrWjAgPbKebFQXJDHRl99Gx+x48QWKtXn5Pyx
iN8fm/pOkIOKR9v0eYWdujkI3ycVNOsi09aTTKqNoU/0if+/w2XINbhi3xSoW+ftYwHzfWBnwf6U
GfKrlzYC7BPhfQJqVcymvHCMUzvgeGtl7qkVFZvLp6zndCwoybwAfGFg0am9UyoGKYoCOlL+6ab+
uthEnZqQd+ZKpFqo/CO9RAIOCC+42dYr7qtIl1Xp976fw7LwUqBBoPaM1fvtF0iHWjk2JqsJBWyf
38rEaE8tfB9IzOSuMa3VWrqHeRtE1ti/AQSk4jM/A5Ms8SMTDNskirLNae8NH9jpeSwapnDUFCH2
HeLnXF7G1wS0knflsVPav2mCPX7uy7xSWLAETBTC51Tvz4STdFxcjB0Htmh/NGZaJX3vpnNWBQNV
Eg2oH/DgdD9ODN5irVzsGNvVJaOIlZfvbRWSaExit9wcm7pQa0PXIbpDdprU3e1UJCFlz7U8Zeqz
LvgKpDu2J4LZrOzKlUxZ0WUt2ArPFMWAOykb0lrt/xVDHIamdzoxeYtvysUQ+CcXhhomRMUWDnkj
re3efdNUXdcbT+24HDuZGrXSCcmNLBh4UwoA82m7KPs+4SzMPSZ4rAFqhNSdM0/CeI4JAjft7FSt
aqqPLSzsiWt9F5leguZtZto7t25k3G1qmDY/+MxBx7ybKX0Wvq5o+Y5pwKcnKO0v2/Dcjx3AWdhJ
TQ4CaNmLRRZW5JdJOjUNmtGdd6Nixd7qpxpDOrZQn1kZaNFkIdf9wy4iIFyodkDpasNaRzw3w/zn
PSWu2CwIf1cZYKfIX2lrn9DQ1rfRt6CV+H96Tge52U6oLJshKtqQqccQtJN7qIplWwIPIouLQmP6
GtNIhh8nWiNto1rhg4pugDrwyagJmOjox+ZlcvJT3cd6PQzhWd8bdJdGfl4SFIMifro/5AcvjPPB
MiLMOkadOwJpEnCNBT1WfHgIaXjsPMoEMG6UKX+iqKkI9vvZ70JwEmU/RJVMCVlSXbWq41GdbQrd
9uMRa8ohxBaZilxIdEaniA7+dvPnzZdbtwpHapVOovZ+LRI8+4QiInO9Nsok2cR4Tc45V81xcHe9
hPlPePsNVbU9fI8LTKUg8ov1nwSHKx8BYBP2vcRhyG23gasyBdvj2iVp6JKRE0N+LAxPA2I6vyky
42/S0vwysKDlLdEzpnALh3ASR9K8RhRYgkE6KaFxGPrqi5LrzkCQWssvnmCyOUdBZheCVzHSke/K
zxS9eEklbSA1TUttdFjE6IZFVY0Hzu4UcJ6BAbSiN08nALruAfLeetiGrIHvgRz82tVFwvZglob4
Ku3c/Go4kAxnOOP4TkkIiCU8M3bZKm6jQXcD3V5DXUKRnDLvggq8+qmDM3GmpjISCcSg1bDIQcLJ
zq4jzXNaxGv9/Yu8bBQ+68KsLiBh0RLIPNPI4XJvStSuX34+TZ5LzUgyJe5maSNb5AYmV7DuwOYI
RWJQyqzIty+osO22UmeVPuMwrtvLMGV8Ppi5ZlJbEBoYXK/doN9DLk3LKUBkxCB8+pHobKGNSHtE
+ONl4tZEiN561iwscsYCgc2y18eLD8v/JsU9nECwKDVJXQzWd5YDGxO5upnI+1Q6UpgfFizUjzWF
urCLKVUp3C749llBH4nT1Tvfa/dh328TD41Hi0KgIhI35p2AmNl86So1/WxB0l2eXV9zvXV0qYqX
TDA3qH2hrXdi6eknqOMEX0VCRcsm11jT4LNadZLblx5e3DsuXJW2T7VwuqnP9rxpAvNPD/pdOtuZ
8a1IDzi7Y7USrABY6gZD6MmA2U9VNofXp+Yd5gxZEbn2EDUCvH+twyYlC8P2zt09dOEfuEhwcGxv
/lnvkkoUlDWp+8+3j/PTKF3Kx8I259Tl+DbPCJ+NpAfMGQosmHIdDr1JcKfq9L2XoL+lTgGUITSb
zBuyZCZ0OWSvCZWn1hYTvrlyy0qYz/nIZwjZPoXyyCZtWfpB5I0cpJVzjoAQMaiumuJftiXsahXK
gYKHsjvxtOzjlz9B9vBIcO3xVrXeP2De0gCK5MynOu79c7nI5oKGsSl86+4Yt9zc2WfHBPY602Go
fYT1VrnZjwv8yes/GDLs05ess27IOvdG/pUFDQPomEYbPgsnJhTxd5W/dyS8Ap6V/DNoUbTcG/wc
lXJO/tSz6qYij3VNfJ1CarNdErcJvsnutFMRzO7TlBD3FIU0pP9+PZ+H5hBJ6O3H8tLc6ONPRb1Q
jRU97kE/MyPH7qmBWztvBNfxl74mUyHtskIRXFrqOLIgcwv7TnOiQrmsKXhpg6GbRNiI47WYD1Dj
0zqEH1/K8fAK4nB3wS9wnVr9MkiND/YQKwwQXwHPQy0e08HPmu5Fk3d6Cwkbwi2gv5t8g1kqSOou
hsvutmwL8IrM0aQzSAstCiLjXpM4zgocvj8lZNZ9117+AFcGx5o6mWVZyWPiAwuk2V8f3fw6Pt1K
7cFYHeTeBHegdDMtvLNySPz2pqDU/KcvF+bFLT7WquxPYaAXxL7cWPdg3Z8gqIhBUtjBvTQ1C5pX
LF6QwV5vILydhC/g/fJx+Tqv1hib23xYAiPjWmsOMNtTBOBWfkpAG3N/UXjL7tQr26xJ2Mtyw5qR
3MTp4KlGO7Gb48cGpG7mrCwWUcT7bL9mwSj6clT27FtI+OLs4zyx8IEWdYSxGu1Fkb2qUffzLlvh
mFKuHFAS+avtONbsjUHZk9hOFp5TIc7AzZNn8AgrpbFFRP42WkxlGnOKadPf5XJgpWo06jVy4bHo
ZK12dRU8dxWOh28Q20hIq0KrsBQhsKlsCMdLszptvWUzIoCIeGvybXclmZbFIqK+A1QrD8/voDE8
sS3120C8cdMhoiHwII2hyFXPI8A72RZJNeHbQrNpzy3kG6XUvi35uIZWSJWKfIAlAuZm0fQwgbX2
pCBUd7OtiRo+Pov1l79aNgyOVMaqAEWOMvDZnTkfei2TgdZfsKl5pyJOgqhvaBAJFDgBPTAlU6qo
/6iw3WlCOMg8A9p153jRfvmXvobFZ2mCzP18gsf8XjdAwTQxs6gl8AL3kpk/YseAoLCuw9kPP0Uv
qM0cyCNzjLqp9AUFJOs8TNi63SxM3uhYabSWpIgPAToXgU3iXisTZn1No/qJhwgD8bBAF9rS7jt7
D9Fbb2BsHa0D/XU4Wldsa6kt4svWDft8YYQ4gQ5uy1sQVIAtY/J/78h+nbfsOw2nd4Qm+eEP5ppf
now97P4Mh4LK0rSHXB4U0rjhChbVEiGjGnw7/LRdHrs9sEy9WQLx0moQbrISO7/K4vKPeVv0dsAm
OjcFj8dAwOXVeAE9WdxvyMsgJEVvqN7QkRYhGVDkIuDTYP4AeXQkAcwQqrIShOCBeMGTDIluLadx
M7+N2x8Jnjmwqjvaelvs4Vo2i+zZI4WeB6odoNvD+ia1CR7MYe0RB63xn/iqvHbZVrFzueWBdbWt
5lSlLv5vrhRDvkoRLCWvFgBxdX4eZbte8manGl5d/7kzY3sUjjtdHBN9gZ6z1Q9eGnKLOMuqYQZc
tOL4NqEzKiIQMhR/sN0dXOjhux6NTCOsvNQwpEz13Eferev4yxaBhljDqOZDUs3YSTS8arHh1tKs
Hwi/uyrSJBs/t4SU4fJ7GSd/1ShvVU8KQ9nCccGk9EB0T3Q4kpL7z77SnUDkGnipdTzO7B8Bk1ba
Sd8xL3bD/pWHbvJ2gAv3wJ2u2Jc010Y2pSs5xhfv19x1wAqi47twkxRYwRUuxYCJDnq7E/KhaXkE
cqdv2BckvancZVERWTCJFZFb9EIyYOd7Oy0BgoniRN7Hayn4QqAA649xbtrfxuaixeaCN3VtD+dB
zO/o1ITKDNhl7YhRDFt57D//Cw9/AWyaeKFeXZXlgp/JijWj2UPu93MPX/GhlcB+lxCAYx86a+bN
yyLT8iTc+9AM1QePyavLaWwigsHJ7N21VT7Abx+F/SSKLqnkch8Mjb6cnd3qsurQBVoJVQj0N935
612qdYnC7j43A6R/WSnS2Jy1/s/UHNXA2Rz9DybzeBLjfB2eL3FPhOomLysya3aym3Dlzo14palQ
z3iHTPlskaaFRj4sxIfc2j7rnBQ8I9YLXl33ITHth8AX7mjTNu5/Gq+ydzxsqkRo3ewkEkOggOwl
mv6MqrvukMlWGALxu//bXuU/LiZbxcEyZuAe5F8/4JtIXNdoLFFHbz5NBrd5O6GpPFFonx2EcOdE
nQ0rGwxpFqNwXqvZs797z4ZIg2GVv6HxQMOc/izSDRKFeSeHCJ3FiJO/IDr77J3YEzwDYdlU94Tx
dfwxPOBMaDBmyHPv/Z+GB3CsJtmdrRmZrAMa1H6y8/TjZMgErmiDGh1+ywdoCFmmK2qUCIEJsuxz
6447z3WcNVi7gXOn5zI1SVQg0mcqJapF+G5ewoaWxzo55aBLIeL7RidOFGd+Sk7ENAw1rT4JXsH7
tP9ynTIQy2CiFZvE+I98V9oh3jfREH0EEVto4RfCyUWkrMluVkMHpw4PXtOsEBHYM69N2v++J2zU
EZqDaWOS63kdIO2/zVzRc+3eWRSVHtKhgwtyH+FPXK+hR6WeOovPzqU0Q/4OQqpQtF8B58rpO0Ns
TmMyRsxcN3Y9o5hj3+j5Nr5Af3Cne5d7LYlxeXNvP3U3T2iCbwjksng9XtHSXOp8ve7oWlYD28+q
FAtE5zw5jUfgMMEiiPiefviIlNogBBqArTT5rKTNt++JO0IKoTi4I3YOdNOySOCwVHfTxvEntRVo
3ylUQIB3X99m15m3mOdcqdkL1vziITgT68Ku11y6qdk+IqpNfPLcVx1ED8lgrN59X1E5NQBKV13V
ZEEHymus6pCvrfck+rncBTFGru+MbmP91GjBAN+b730LAf2EmsERA4h3isz3yz/rOP0O/hWm2hkS
QkS8rYBNVG/I+lNj0N+wAFsTBSRp0vHnP2hka3O+q83FdqU8SXXQRDtCVeu17rC7NaPUka4tAKLZ
M4LymeLGbBlijzYKrxFkIGRMK6uBVYtmRf1aJt1icrI0d5WUY71V5v+dOpM/Cd+vCt1mQK0zYGKw
3/83TUoyFngh+g3sIJBXfZKO9dnlXtiyxZTC8zzvOWPlpZYJzXhUGuItgGGMd5lBiCRrL0me/e2L
TLajtWiROjPEHHviuZm3RKCDjMezEz/YjOPI4cUGEpEvH1qs0n7crKk4Pn9UMfHLoQSpvpdMcED1
s8XtwMbQ6QCi8LgIm5YkpGs8vAXAlFur3TrHHqjrHiy8cYFSUDKtQUd45ven7iovhNRlEfCrEvp6
g0AH2VxTZBEwBwmkMCP/7DtkV8uqRMmo0l9HC/NBOqK1VsvwYk+tKzLSuljQ3PKD871lpHIPisEq
zpjBloK9fCO5Hd1aWFbGsUYNaPSU6l6doc3WU6dwIKE8m3DiM5XxgJYnsmNMD1iaubiWXM6/AF/6
NMdnRiF3CLUWSTIT7Q7JxFURMqjKpZrFVJk19wpzmjRYfRI41OcsJUR6C5yCmwVl2YdFxuHn2l2W
gRRpaBPBsvhwqPjrcwJMsBKcKxJQMfLO6E0U5Lka9PyUogXLPGWbnTwddR4EtXId2Z7DnKOJZFyC
ZEd5b/q4hE03inRj532fxGgx0tGDHPbcCT3cSY4Qf38xNUoA2pcTcWv4x519GF0UYVtj+KgWsMrN
a/Cguj0/8d/BkVWNZLF37HfuKndgXcj+WrAt8l4Xi3rjgvQky+pSRHg3NOI3+HOcTKKNyEQfzoK7
SrQ4mYARW4wuFmKp1G91n9x5d8FoHW1e9nfxznzi5sOP7jb9VziJxtgnfpRM/B0CueOq1XRonp25
QmpXPTdi78z4lKifN8NPz9uyP8ckLyKluwJeCx7VX8ynEdO4bAhNRnOk0wd6x3e9t7pM42D8LE/5
wBIhORAVWjTCUpWQNtvhPwFauFEIMThfOoit/VEyGqoEjhiwCYJzlymvvcGmQ/FENrBBSTcfbbfT
AvOiQ9JP8C57cR+UudKcEjvDCDKdA2VepJ0uHCMLGtsOdBeRnwcdD0M9bYHH9dgcYWGAcHx5ohEJ
sN4z28x77U4nBL+MQYjcwaW7zKTimaREp1gmMW839mGIVogzqkot3zNoR2C9IKmwq4yqoXQ6Mdk2
/AiW2deXCgr4F6+6Sublijc0hfMj2crM94BBAgd3VK3vj4IVHp4lpT5PZC2ISdqRRiPh9g+p17nH
LQxZ3XLEW4YAcgG9zA0dFm0u48V9CijYtISSGVS6/caEYJ34VkipqSY0hKmMwXLNiVw4PiGllxu1
DGjFSEFcxQRnA7Oei+hQD0Bnk+w081YFnnL2gy5oAMX5MmmtBmoAuiKIVq8ba22DUJMnS8M/0rKA
iLf+pjM5FOXYStG1bgDx5otGNFSTELPtDLIh8XIzPmq10bSrRQpWF3N+hSTsc3ySLGiukcZLna3+
52ur3lr5gnt0cFnAm9fpk76tMHMfsKeBcS9rUN3RS+VM6gt9IdSnGgSbF5jOEu+KMXB0D9dJW8Sf
gPkZi/J2ocrGw1iAWUUWclKAtt1bBQGuA3ITQtAwuGfxAXSsV9GVTjU1B3rTBBiKZlEbqaXps430
IqUEFgjXatW60+nW9u/zbdB7r710mKThQJX/MVwWBxQikqS3rTmpQyKWP0X7ugSFKscAVxc5ejqi
LRQ+crC16ZAOg2+y20MmNNjKjswiWIaDhPEscN092cDTI9mOidii6kzAeW79hKGeU4NIU8v9ntrk
86H/XOnWpADGN5ON1tlPHroo9HkSLC2SD4jlbx8SfbvcrvSwxp6GBrmLJIZyUxjmCraAPAD9FG6f
dGNNago6lNGJfnHNJe6Vc/lW2t9qWewvsKWRkXjGeC7Wj5ZYWHkghj0e4On7Q0++JCuhDr7Rglc6
kwneq7L+WMznrCDIJW57kqOhDe3Xvj/LUW2u125A35vq1+JodBDfQ6w991Gu+CgiRXYQDwDWWmII
qY2TZNMAMpe5ES6QIOpDGu/X/S21/MUnNfWLf8XcpcIivWE6t+5NyNu4BH0J8Haat//sFcCrf0Fs
RcYAKh69cFmdUksROVLH2863Ud5MVLiWqF9mixE8JZZ0ZIYEa4BqKs3rbbvuAIetpRYowlsJE1Yz
LitKv+Xaf3u6chDR1zv4G5DZRA74LRPW2kM73qSh4vNiHN/uUjmTgvnDqTv6EHXfYMjf41t5TDsS
P6qBrwJ8rum+I/m7XibqXUFhWn5JO3t1e0GcmFO+CtJcDWNcukisgjZfsS+IE7/soicJ1cqUHDLR
E4v3D5Hs3Ex/hd1ylWNKAc6mUj+nyS++T1xkwscP7YktMFt1XsS2KkU0g20y87haXQ1OyYviU8LW
cuMvp1GNAuENnfWzrKl7IC7hxjpSLQ4g4MGv8seP6nW0vSmmlWOrAUANTsgSnDUAC+Z8rQHtP+RV
qzt21tFaiWmbyjcmc1NDjF7A3+qtyfPXMRfntO5Ta9zs7VNpmWBfl7vugbLmrS7vnpWONUDJjA1G
0tT83X2zWUJ9gVBcDpkoryAE3vlWv3rCRKtCvKeLae7v3JL+uBiwoFYAA5w5a4t1BDDm9DARBBvm
Xc/NInGpCxCbxBsWEKXbldnsUUaR3XsbSSWnnChcsUHvcTNDbzeK41Gb3UTeDF45/bq7lcqWxYmz
2N1ppGH7Slkt7KUVYnjyAWgebe0l6J873umYD6abi4+xvqSxluRB+e+JVqAEGRbZT+MP2VUjjdDT
r/InHaxI581TtMLspJDd4Zv3AaIb1vYl4PQ3O6h+8zn3gn/4CL7zKtNGbX1rmaO3Rk//bM32nJtS
TTW8dcgqQWGFBx25xi3rodaWhXkDuLf1cEt8/yX6aidk27AdK/92yQFw74h47yWUDAamrp16z1QZ
1Pfax3HiSIbXvAOrR36vh58rM5Zaqxt8ZIVLOcsZNAOxU2dWUzKy+I4X8Qh+K1MWDz4491bWOIpB
7SCS6HptnQFvkXWUWOqw86odc/xH2hJLkbv/p1Ev6RWMGywoMY99SLc5llb6HclMbwN/Wa6gQd4O
T32/mV7GaSWFQ8mIKLETbtw0fF6KFba1DBdR5cEvfx9U4L+Uwrez6439ITuFS8I28cbHTmc1ZQKj
3ucLf2XT5pCuzb1peaiI4TNDALZSu8w2/6tKy0+mFlPdLGWb+ydnkSYBgQzGJqD15/0KqaZJuex0
efxYNmVpNf9Ylq77M6qYlQPDZdlOuFzp5icmg0zySW28Yl+8+B25rUW2xcFeKsiHafzGAg3pj+Wi
Io9JOMIXEV3NLO5tZA4ig2UJqRJ5KrbFuYS1dqzCw2LcIDK6pyHCUnHhBe/Xsp9wvFpcRqpni1tl
pyz1J/VE1ERWi6nHeVH/xSncGN/HaPRCOw3NjYFAi8/DjVugbraJpeohFkcqJH/4Lv8ks9Df5xDH
vcTx3zcAQor3Ejr3sC1+8DhLIJ8jlhdd70/SPIINECGVJ9bfK5zjn6Xr9nSTNIwZA6lPAUbZ5gSw
VUI71at7Q9RKQF68PIuedhL5NXu5FmJI0zHznk/FG+A6SYtE+9xHKfXFChQuK2nmHwc47QBLI057
1puLzk1ADh4T+o4j0VEAC6dMW6Ds40bigPXyM2huHrN+gQHQproFSQ+9/dbusQ2oeGYl1cM+Wp1f
rZe7rXOOABDzr3bu1LcR6vW0xG3zhlsLBOgxNEewDIirOJ39N3lTd3NxhQ8TmVrn81jitYIm+san
Y6rwkol0En1R1qLXc/vJN8TOFa0girmuLSntDAoZNO1ltfaU1wzzQK/8ZJgPbCTSFTSA+5xlOwgu
lGsppiMA0K1LLvPVYgDg4r5TpO3GkmLC8SaraGdSbAOGQkAJ1ZwDTZFJrpnheiWoBki9nUQm2MwN
1lAH3IRmj+na11Ouj3TaWdmuomJ7wDkvrZ3duLrmddmqnVpxBUfd2J0Zz0MKU6EP2V0zdz5ununV
KfnbAltMbjVQTCyL5wc0rCASD4JmrRdmfMT/1NXmsMYys7ZTRyrxV6wdkfsHc7RH70tXfxsWktRn
qwrfbdc6eRS/qr4MpQvqGVmwAnUbApWeondYGcRG5l8EGt7rMd0h1hj1rPCa61RxMXkKB+JeI43X
8CShgc/AptGaxorMWDLt1/Z9A0c1QnprjTArtyDUvmWGIVRUgbInFC90Uj8o5sa2/JAz65KTKuxO
WF12WxYTP0oxXl36W3PPIibZq/5kHK8tIoJHZBgHWc23W8LgF0B94sxDwSmMF1WH1x7TVSlVxpqZ
WKCr9j9zI8VaUXKO/xqZXf//gCessVFR0R2BULzBvNKgVWciCR5fUgX+PK3XyfoN/dNUsOtW5a+3
6WCwKmVWokck8/g4rfJBAhhdksYFOrqH8/PNM3xZbYAER69ATm+sVexbj3wMjDVKAh9uKlsptir/
6SZZD7RFyBybhEQDrk4udTBs+G6DUKhIkFWgI6CbnF6NBTTh/NKOiRHwXPGvKl9hYXFWQqdWt8rT
OZL2KG8bUPuISBSc1NlR4SjuBBLKRx9KLGpMCGHLbHDUOugyIviQa6vqcqI2Kanlc6xIskxmIowM
PKJ4pJJp3S5bqluNH2MqhaxORW7x8X/79GPw/UcGiO0o7+P9oAzZvGFVwYoQPsUf92kNfUwyT7wb
02LE+p8y2P+Ta/42ZIpWLraUaIdmoV5n2OXTpueYfNv75ulBUbKNisS28hhwJaKf+04wPQo7+Eic
+rTsDZcaWtdYAMOIi+4aS5nw+Fsvg/MeuTSxVhLzWZxoc2Z6BxnwpedeBzUMBuuoeNPIRoAG6A3v
F1+creH4eyXf1ZSC9F3Goxkw08Tfn6WgvoF2lv9OQ7xOhSSkfAJAuMaYw4nkaBL6+hoR7gw/wgp+
9Jw6dLFo9RaP2xgM2RuxIsjvR9PD7+zFLFpKNPWgiWRQcab6yLADFpjtAsyFp6cEnvN7wIuXNMog
r63wpB8B6wenuBtiUPq8bFMoqj1z6KhwGl5vOdopsxxwa7h9Xyxm5LQD47Q8aVvdLomj3iyfPnTg
jGFXQ8f/xwfJ2xdFSTRIdbHdhTtVwURAbxOJhgRkJw21Lg3QWquRTF6X8SWD08zRb8i1LRH6/UIp
nsguE1HwlvIUmJN2cMXLxrXz1JxmVrPaA62nc1F6eVZbPUmFGTt8kj0DDved9Zch5uJA1P3QHNpt
dYLf651LzTItkuVeJfW4bHeLkGfowMf/wQNRGOcBZlw5dgvV275E6HrCUmGfI3IZJF/bvBbABnKi
AzyIeADaS79BX2nKd23BuaAIcDlGc6dBZD3dC1/7kTtU+T82dTSqOB6v/vfjn0aZEqSGHvBFDl/p
A330nhtS9fJhUCUjiXE9QGW4+Y0icyTu+t+cz0iKF+0e6rE/jruXqcwKrAfPa9ATbWgDXB6B5NVZ
YLgO+KxzBSVv2NDNEWKE6/h+RUBa84L06XjuilXh01BwErCR0OQ8s8KhfErGQI8enToBBSDaR1gR
PDUQAnskLXdi5+TodsdWfKDV49u3csvO+KjWprgQdx7hMwro0sl1XA37AV6ZXDW4DNwaOwkx72DB
TKSiAn6MtxJNodGpBSSVlB+FZUVmAkW2gR9khTBM2/0zVt/mEw+mepyApfJgozaAz2VdWpcyxUes
QN0StHcqfwvyhyAn+HWZeo5akpJ4+uYCVKrXvZffgdW8Ueaf1uYqFV6gjEv8lYApqc1eDFmnJgrQ
8Jd0b17uWrozdkWpUnaUL9kzQ823DsV4pjKhnNEn5QGCBTGCQM2c2uumyxwJoKZnzh119KcmWR+3
4X93qa2j84KhQ3wfnTv6M4JDWWDK5UVNMUWL1tQuP/fAiuoJCCneARBbqTRQZG6S/Nc9VtN/hdLd
/ZUtOHF18XmAAGyMNd3juv2sN9aNV66+9ZC70tTqzRloM+qXG6bI+HmpKo5X3WoE5eKT6/yOPdSt
SCFIuludmQikHg2apW2cp++76pigPzDpFZdWBZvHQULdHOI+BTahxY1GgBBB+akSQsTk7lud3dx7
AcV4nFU+TjarWKxaIxS72yMPCUSL+892RqFiYmpsCyNEkkVvN1bTkrW0pPinBKSvtEZVzcrzvV64
Wp9sCHOb6m1VJXZZV9QDzZ68lcVK15a4Bx3rQlBUXETDG0v/9owdV7jnwtYz2uvfro+HGvpL7OaS
VSk/1LJ5gnJNmgrHsAF65i3gZ6+wMZGpiFCujk4TDcO0E1XTs6W0EZdHs4Q6EuwUkMcXYkLPpaoY
Mcjhqscdp00EN3kUpSxTNyayonZEFt6Hk2N4v39eRSMBkc4mX4nT82ebafeWdpXYEGTEJcDkfkOI
1SY4f6aRO5UzUmGiwXmbNXXwMUQyIsELn0ad/eQhFNXVL3C9yZaZIGH3FDJ22QG6Zmct9cKtEww/
plzf7JcaijNLuD//ms32yw5AuyPQezs0obH/YDr/dqBJ00pzw+uv64SnE/r3iMRli0UBkNTfTGhv
5kAJo1qyVBDDzPYtHm5zq3cQhkbO8z0taiZKQCw+C773QNZ3XmfhotqPZtqn2unBN32jTbvkpLmG
Rbcml9afb8iVqp1To5Q01FJxgNBqlEeksAuBqYgSTbgyZu2QTNwD+zqPZ9lrQr2NAe2g5X826pdE
Mu8V7qCrjL0+sjqXsU66HIQPUjvd8i1/9SuirHi64GGSYs7pO3v9HDEHKLWCDp2z00zQFMeZr/pb
jr4tpQmGRcgLZ35s0eqrhepG9tapVpru5Zs2vggk1ydzbNpRiQCnq0q5nHBGxNM+axVj/6q2hwY3
bIr4vcpCcvklsr5XKp9JKldPEjpOOzeBwvDWtQ2Z3kblKVY7TDm5H1tGLdMA6fJJNhrygNU7W80w
/QME0/n2ExWxmvPmH3bRnqp9qrmYgQR2wfjvNejPRVqu2+UDQ0Ik9QxWysYwHBPIt9dw3J1zgCKA
t8FqPEGUZqy8A1oIXun9zxUWOFAl/Mtv5nzwTPVAAqeVzvDE36EP4OCEq9rRmPWEtynWjev0B6VH
0iIcO60h1Zl9FbDKTgXDeM2kcItFzmKrClCWIqGvE5gum8shcLUVCyqcxhxl+QtMysOWQpAGucv6
gjF/i65O3CKDbSyoHFWHhV1DC2hyqbUyscCTxHZ4M6MO5Vl4dDn4BYDgwn0E9SXcn3roBLqHMaDR
YvcV2dJjLP3k/hauQyJUDO1XXKtUQzQqBMkV3IxdEGRvK3jGstoY+prTvu2I/Rpf58BAY3R7o0XB
uB91eAi7gynEQaaKiHeGJrleMTNSOGzVRLBhyNjbYsC4gr5aB1oIUMOEMZYkhEViaArRKVrG+VVE
Xn0tsXTOeDP9OTeJeDtchwN+OUHct5H4lKggf+jUb3o04M4qxsv/wlO+GpVcDIk1bwKBiE7LjBWO
FB4IqE66+unCN5tuFATXPObHFB9qWeZ0vBouiPyD6d8kI4F3LsNFUeIg9Tdao0fvs6JhsC6zMY/L
MQZ9LztVFVIEiWtK9oL5nd5jgwx4E4UajtBviFnk8ptn9qhsQZhxb6BbAO0F7IqDEUFX6vnvYcpG
C8z1RdlNyRvMOZm+QQwDCP6XYh/g90/jLOXjtvzQ3bPZw5ZpFIX4hPytI91KBFuQZAdp+/oZoFjv
VRNGJ8zo2bgWmIQ9h4Q9bMIAOHiJVqTIzvv72s1kAy+qh9i2LWjO2IM02tuNNM2zGqQ2AteiSxb0
eLd47kk/oc1U+4vW712eEgXpbL7tqs3sZJOepBaLsMM6Xikd4Za8A8l9znelIhOYaOdH0vgUXwjW
U884x7KzXtCqvGXpSV3/H/ZIdm9CKrr3/B2cQVZXl+lPNLZxlA78egx0VAL5bkkpiOyL0XHfVn7T
O8n3EoM5fzA7qaaL9Kr87ue0ZDMt6KP1ZMq3RYSuty2zkY3Ve72y4jNoP26bbOCE5hOg04k2e59w
gbN8iBtglDlEAiNzq6+8yA9LmaSp5RNVtPVbiB4XZCti4Z1NzK9Dn3AFpgfMiIHoPM41Cj1xS5GA
OwR6XKpTGcOpVlxVgV9yMbpk4wSOhArusBWHixGvjqXI1IgyJ3PfBjRpCC7zN/erYM7IEpZNdX+7
RJbkCWd0NXj4YsLPop6dZ75MkjSo9ETXqpKimAibI+2pxhzYVB+suWjE9ht58T6KTJDcVDRXK7x2
omVf2huYBEP79zj3wVYSs2wQKkAV5auQi8tDPIYEYyAZtxDGo4Qp8FgU0gLFhe6v2BKYsZ5pwPM7
tG7JNYMkx7O/G/p7540qLKmVrV7E6wYT7zV5uyVkfaWc/1vBh3/9Ja3bG60lhnrNKEKOpEoYGwlu
AJ7zFrs+oSHhzBee88nZ1V3zc7QxcFrJlz59DSXPcD2xggJ1pZOvKuWLU3SoEcXg7G18wcTWMFZC
4tE7HJV3xl86F6dPS/rP5z1E8Iw2gjWxz25KkWIaD5qZPid6M+rfkonaMAzxg8JQCDbqRAYOJOKH
o+LV64TznDeIBGZZh7FskVw2EImLgv4ox/cxTwz7Q1OkmRtAPNi8S1Ys6hxsdf7jBqsv32Tdvkpv
tue007tz0SCI4aludI7x3Rn1sC0fvFUoHm+1QKu4Sb7qQVg6aBGLGAVn0Ib5Y+OZZu4R5xZH4qBg
1NKDkTH9xWgBxYQXCvGozG6DwKfJA/N9bMWmbhD1Cl7SXpGD2iJURHFpF6sKRK1IAu+cIctsu93E
aHsq2VFZx1PUXcRFfs2eKnxEW5lorjzHWRFVLO2ZHr2kyP6kMGQL+s+cXORXa1U1qnHlxmT9wQoj
eUS9IHgjV8lV8ffdIv5FDl0/aaG9ptTCDNFxOqt3dHXXRYrUoWtPBWL+R1Whj63j4Myk63FLCkT4
IqZLHtNe8n5j5td592XFcZK9MzDTzzNVLSjt12AJK37fw1Agv3wKauao4UzpKBH9Ss8le4/8C4C5
kYdLj8wgKH2a9zj1vimuRCmo8fYeOfwmUxJmnd+9f5IqjfumyTTbULTZ+3DP0lb1HlhCr8We0rBp
LEF8IayaZWfthKPhk6EAol2Uyx7SttH1XXycgYLG5Ee296G0s3ZCtSG37hxrhHqsuI/wvc/SNMoZ
BjWwhRWiiJp9VGuLNw6mt8rmgNzUDk8kdxOcsyzwPoAvl7aES/unjNLyv2BbeGxds8SAkpBjghVI
7+HibrL6UvdzDmYwOsXa3AAziJ5lhW/KVPcKWQRx/qaNqUP1r3HcnvRCvuh6g7MSR0WyK9akcRki
l5WYMB08gFe8PtBjxYkenZyFlEdX/wu4/4MnGoMcphfjF/puYGkaK1w2HpNI9FE6eJTuiMT9ciH8
KI3kz4O6B5cd2+HapVNNCjERIooGcz9ICcQdzq1EptAm9r7GIdeIO0BLO4zHSWTIX0AQrrGiV/jV
UlPBSvIZ/IQoYfN5yOBTnZRkItkuLRRt73evAtPCQfXq+1wMbdzRGiCFR9tCFTRqP18ZHCjvHw7a
fnxRVfC09UbXbIa1Kwo5hIxJ+nqDkDXAYnbSbstOth9WEiGa6tfUhiVk2HxdsH3FBj9KYvqW97eS
I5S0+RYT2ZCeOcl7cWdm8yyryfVyIfYIFsIypd3moat19jw5J+sQVXToU6HaWOw1C2Glc5f0PUTT
zuh8R8jc/YD10mK588mhR3zeWkoKHRU59hJ+Aw2o3bWNBaEnCAfSLc8Ank69vAGBluD5j0WrolQA
NlfvTvH9Qsk7SeSzMXDmcW3w2UDDzbHKE8IXbHSDm/KuXmvJjYRy0FpXXlTcdYHVS16DixdNU0LA
QvPjvwAx+LZppAtMb7mu+LXRdxi0Gqzh8rcr0VtBrgYVdx6SdT1ECT7XIkIaE1yDQ2RpXGdaWMGy
KDRIwqbi8Q72He/if50Vii+F4KeFQ4bQfl8TRDEtsvPagQDxqb9dsKPjQR5M3kZsHCsKsw+68K+y
fxN1sx66vOIQ54GnNOIGGMsOFHgCOEhyfpvUxgn5vc7IA33/jhMB864CxFleR2gQaDUFCu3FDZkm
+JhDrxRlY34pBnAqMO78Uach0Z/zfJR94g2/445Nl2+JhvZg5cSNlw54Agl40VIx1YuA9k7TryMs
C/unFLoL8mSQ17j3cZ1FtPP5EcXl6IRAZ4kFkg1YwV+p6ilrfMSpZLCJkoxLEdYgAPo3B6/S2EEJ
VKLxlC7YYFRNQe4kJHCPCfWzbkK9+keUBLJywAJyIxRQ8AyFj5FEHBma+i2kThpRe43R4Noper3z
v8X2usRvKsC7HBVu4l+nhg/6w5edL+jaLMOLjo1mUFRtpBAyN4JFJETVUplt3ZfXJOUsISsS3XZz
gGgDh3j3gUl0Fq/BFhjUaFRK9CKjNz1zuvVi6g8/DyXmMuS0QNUpd4sQdzTbqe9BqACJiwTfROyg
BHvPSQEU2uRfhobLHMQ/k+uCEZ17JDrt6QzKIMoKOU0Fi5dure3OEoKx1u6KjZuyOlPWtCiw8bo5
TVFP/GQ9LTySi/aZvOU+eHtq796eZRbBHSZ0LkSjzUgKMEkcHu2Fb9cXN3YjsESwTO99TpmUGcS9
FVXGgiTYskZtd0h6Pz10UcAWt6wiaTAKCDfHQZU94vmGyGeJSwyalrzZaMu288m//kP/kmpLn/Kz
yHdzTeow5o9c+G8Lnj9mEEupQvj+kiS6hylZaV0LWL/72VULeTqTa85Xuizx9tjgODi33x52FgNK
XochE/JqE8SaHjoCvkNnTe/1iDVIFuxaEJ978+duVmk91iKaAaICqQRLN9ozstl2Gxy93t4qmCk1
g5FgiThS+9daHAMCmaQXzVrlflz/9Si0q4FVUh/fjHfqJILTUo/NVdJ9XpNEfSG2yZss3BKIqmk6
U+zeO8e0Ugn96K0KimaBjm1dkvAw5VPGAvddw6ccpavtuIAKjpvVlXkUZxMi5DhTcT4esJ7cR/TT
lf0s4bnK9CDIU9KlejeKbYLroVk6aCZRh11MDXp43DyczzKQphQJNI0+0ByaQf28Vbib/jDj2WQ3
Pse6TMa5+lXCOKS6EL7D8mthvojDu0Cxr9RrLgTx8Nhge4tVcqy64eNJUOlqV4+QoIz6oRw2hp0T
LXzsPjY+PGSbUByhmkwP7B6qBTiH3QHTCVwJTP90hu2RX1+UpvomjrEEeZqauEjDFDfxK2Fk8olH
gPIqu9ylLJ854SSRFhOEVNGaIAyIjjXBstmMCtRqeth238oZ+/e/xdB2T319sL0eBOm4p+THxHm1
My9WwSt7lC0F6NkNesKVu6+DXRKGstEFjrF3WJLfEUYY5aOuhcgMc2bVmTKuSXBYI1y2oSjepZZf
ABGh7YOCKjzHu6obd5mZ2F9bS7W2MYVLdW123i+xEsIme5qZwvn81hmtNsBE8ajrD85f3rjOIVrm
lTGWQ+JYYA84iMzUlrNhSu+0YDm33dPL6z2Cns6vHR2DpNlJbUq4ndf+bG/7khfXgBEc1pyi4M3w
vI0XdtRDgm+6MW4d3eSoMeydN9+gy4+nQeR7cgH5WpoBWZLbKlTIc2qiTPHakyH6wLMzsodKgiAP
prsFA27Tba5g5ZVuohPRLZ/OwPDYF4gHeIjXxhFnq6V4mz3UWz+bwv0FDAUmOc7YQJzMQXZ9CgzD
Mzx9Acrr7tZMs1H6G8OwO1jlzuKCDJ8Rf5Vptjhq9LTwcIVW+FFFg10brpAPWPkYmXsCEx3CZlh5
uUO8u//EhyGwMaEJ3zd5gQH4JbGriLApQ9Djq6USOp+cIX4Ph9q0kuE+04X566pnZKya3vj67/MS
nwn6WDlcBuLSdM+hlJOvnpeJBvgrtnk2PzJSyzX7JoCMHwVB9qAFAGzWlvACiKmnN/2pn+JcS1Hb
4bPq5eBk4+rfREgmiwATqvxXsQ+Hy/NWYFQgBAPWx+ktOdD2xI03cw/Lghytz4DN4Ef51EJkw8MC
ezR3v7O0KXESFprEn1RKXmklZ3Notrc6Q/0IAblSRPpVx2ZveTC2B85H09gLHoM6UU/gWekzfGGL
EaSg41ROqzPUK8b7SMeDWAuFxKdQ6FLoivCjNZUqRQjSt1lBQw9bN8kX2nply4lYnQh5CqFduCE6
3cdV6GZIh6JNx0d5+WQMgyfHUx7TapX9QuFFiCU2rqAoBgzcQ9Tw05K2QpfsO9LnjWq0N6WkH2b4
NSFtpAtRA0APu9jKHPaXRfEwmsyiR19v+Mqz6tcR2Gw+xBe8Zjz66LCueh92NIjFrZFTcJ6+Z9i0
OyKdEwrOVNg2i+yIIrxyPFUcDr+jW/7N2M0MCZBtJt8uG681N3HgFCO5YU14saS1OkE4zTMZDC1N
Ug6/tvh7wa27aDsfUgB3eeD4Oq117QNivMrIvDlE2lNWBV3QV5ircDIAJb1V+XtfOdySCsmQGJ5W
GNURMjC37NVTeOpjE2+ZEH7n4zc2XouzFu7imVtnzRBeL+EZ9Ri2wcbO8oLYhDVvntTFZRwGvTBW
ukV7cY0vjG4zs4Nha4qOL2bhlYkzvHs9pCjZKpXm3S4+zLgpYRhlfWEBgB7ugRmkOt66w7SJTjh0
5YFPXFB9/lM/KR4H0Nax0nRlPVg8d7WqaSCC8HY9S2o+0wIB4qcpVlRSgLmstsMxy9mDbQO/gQW5
LBShX/X6KH88mPW7UgbbirVJ+QBMnfbGHGnnJu0pUVYKEg83gEnviBVzGtW9GN/mj34+MxxCpyBU
cw4g4Ndcg6GXI92ZYoati1hJU0wxNuxUsO33kuMK+yheU5UkBEE/e6VT1lPmn9qrjUuxNg+F36M9
eTYgIL2hGaPsJ2H5Qq4U0mf+xg+zSlq16yE0rTLmyWqyZSWd5Ts9QuahlRbd5liyBfNLvuapkkbS
O/5hbcM9lkNSN8MYmEvoqjEtQtMk8HbQTkfuIxxdeMnZUgUBizletvIQHonX7ljVrQA4qqI9CeAH
kJdSwGEAAh191rCsuMpuU4JoV8n8+wMNEtm5/q2FOXr6VqmUZTXaWfc4KDDx+jONjQov57teANGA
Kon/UvZX8Vdcq5tIv9DUByiD6cx051QYs7wOq5u2nynjKAEKFLVesvBfAYFoPxybu0zPH5iaenzV
LCViJE8hmjA3JJNgDN8WCkDthArpcif3ZMwurHEaUWvYr6OdmHI8KwnBVxPMManGHPX1DFF4VQIn
B2ZwyD7dukoceFpYzk25XsSS5KjBK8gxvv+6eWWzGa069yerS6QAZaFx8KtcEEgVR8vkjvmX8Dt7
M1lrhT5EioTgvo/qxPcwe30hjgc+2p14exbLkOFdUNItdW5hHZDXK0m+PVqbyXMRjracfE5tq+b0
cQKiB8p5JHjlnydjxICr8A811BrSOQaYv5vC3vEh2EZu6jRbBPakUr2hsFgyPTZvDIgMKdlsjZoX
0c92rau0go+fgFH60p7jnnZRtsdxfH0WfNFZjFt7b+YcQTufF8XE/pHea9wcy3ml4NEvaxdYfKPr
ma4fkptzUMrxf5jOgdPomDoG2lNJFjQmygYM92XZ6sxFlv75mUPZge7EJxbxr72HPHdnJRslO2Jg
SGRa0qbihKoFkNKFo7HN4akBaHi0c/yGJiHHoryasG77vjzRERW5DXLVyeMJBWtde8hRE3QS+rbv
G7VxMlbukE6x1rOntzK3ppn+7X++7j1FVEuZbM0aSKjLPw912FGVc5WOg8PD1VN7U73+T3Uwqmga
9EeZm87tqErPt+dqVMEEiAOxvDpGdMF3CWe62u1T/Qy0RmMz8Ev52Z9dMb2OSU6ghGLTtfX1DOwN
thfdLNt9hZNzSJlCPPo7QJhdeo44Mto3V4IAABhybH/CQ9bbmxsEELG/0DHh8hyGBZAeqGiYC6Ua
Y+ab9Nl68w/Oj039ouEPcb9tR6msH5yn6m/8YjEmcv5AAcUfNsvsaPw6bT8gqDZnfh0FiWQnUN4X
eyCanBUasPMq34eWyFnDqjjDGZWmsDBX6rokiwHzDXtTLNI8F5yJ684ozOHApQlNOnvr4JsFg3Va
um92YJXOAbtuf0BZDR7H61CZ4GOU3y9G6p95gCU7klYdz6cY2/ASbEBT/kBH1qcsamVT8XExMK44
9eO4GpOE3GCDIPnkE37MqQNBIyGoSw31GFVtvzQIrhIB4zTdXZ9K0dx8AHKLzwfMANKk/s38k7uB
5hM83kKIIw0+szCVp5qQNsx0p9hyEdP9BR+h+4tczlO/hxQ7Kmn7MvAtYrCmJ5pG7OyhzNvjKabO
3s/4FCd9Hu5zcL8PYtvvci1fB1EZiHyyElfNxOb6hcVtyM08Zc9m4ngEbq+d9I1RJukd/o9Hu1Om
tC22UpfvmlG6KLEPemcJKuW87W9mMBkFIodk6Fb4+79Igl9jFgA0FpDIaegF2mcqh8W/oobFJd0E
Byuq778eoZA5Bg2fM9eHdCqLSBs/Q54CEvbc6rfhKkvwy4mx9Yjvu6/Yzty55S5EaNYbNcZDADOK
equywTikdbo6FA5QOc2yN5RDa5MZkGVxk5bbi/pD54pFrc1szdW9IDPa+yoKYZqdRHn8Y8SsOse7
pUeDdYW7EWgX4U8UPgLsLt99ouQXCJlXouOiNr33xGXsjCb1LjBBu0wnxKsecu14OzwXKsbg5kpT
PC9PlA4GSOU1KjjlxJhsOtLJcoVNb0O4ebGnaWbBxKzIqlOOGy2i72fOGL1MQtZqGnNAujPfQbJ4
X2fjbVz2yfWiC45ZFMu8qdLF1yc+NMgcgcInmfF6evIUCYY9YF3yz+3JpfYCokMEjlNW1OXPzNeH
2WGKOXTHp9UqGZMasfNkNLVQlNSBDEzq4Mc07DP8BGFOOVCB3qelqW+ZwDxKXTY6gDQM/0C/6CFp
CfCRax61foDL+pb/A+RZz/QqyUIySbH++QWYIz1FIFhq064u9W0F/8uyAJDwUI9RPeTQV99mm4va
t4limB9srzw61fXQA+aZDpLxtM1vhHjCnrli14SoBUNuIqFuWZKXmu9WpFLFAt9FyfvRMOL6UHMg
TLWIF96CSxJdmRr7X53wESAa147JCULqPFMCC5O6m7F1yKFpYNsi6O8tnaT29ohPOGluOcncjkWO
0HnmFNHZg7JxCwr++A6jS2pzf1mA9lOEPa1FLtUzGNDxbrrY2GA3JpPj9VI82DXPxitE99HwGqU7
gSXNUDPiSZUy6hDQRymAiaFXR283XI4/VGv94zsW3wpX/0DcH6HRToVt56Np6Q7xVX3FwBi6d5hz
e6egy3KRmiWaMXwlFFZHfxP0rcPDw5aB2/NH9/pB+QAH3+RTA6+zGt7Y5PZyzvu6I5/p8xNv6MKB
T3UqHmfqJJHuLybV1kluNmq0hd5sbWwdRoqDOXb1ZTaoL8sPQ51ucMbJqoExs+b8iCU80TbaWqH+
GVduZJJyXiJdfcSm5RaclZUfN/scVPBW4WDmnquvIOWk9oAMtVOXmw4mwHrN0t9OSsVSjMrOjmB3
86dd2wOfAkPNBl11WxBWxFGBnzVoRW2S+EGflK/1MoKzTOrJd4laehjiAZcoiel733GiLgyxv9A4
ptcMupHPIUTvtZ1UxQnHp0DC3Hkn/PY+R4X/maE5G/Gf79y2Gaeau23KQnu5Lx6AxNkz3GA3ZErA
KNv6z3XNWJ7uP0UfD50PWTkqRfQHLd2uHakgRkUOUAYxO+MX+PEKTls2KofknFYYxkEDBr41MVoD
FZq2xnaTgmVz1tP2B5eTGGJNQFORiNesd2jttTAvgfu06rFsMxdo+sPMZPl0X/gqamtg//LlrTAl
iX1hf4wex0No9PYsBCW38S1kFHLl4J4aG08te1baXG5zb6eoGNIVMIMVZrd+ikuXfiQOTJeiJ880
zukC0fFO1zw8jSxUJsb0DYnww5ZnLkMSlMygTjRwE9vfJX5jH31p8D6I/bISGYduNUqA6tWzzCh0
xnKyHAz6XSK6nl2WsjQ4+K1v9ClYo1Vapxp1X4tzE5wBvnl273HoaUmakg95WKAAWv1Gs/Sgbt6q
KXzQGPiz5Lv1rWXAIrk84EdOetOLeqH/aN1bzQDYh5iEIlV7lLOCY+CxbCJOf62BNz86grjbo+d/
E2y1W8nkp3ygvpWiM3mGRDmvfK/RKM4KuBcTbNuFeqv2PGJKRV0SY4U+KX5nOEwihZGhEtuOsgmy
km/VGlbvmRWyHRipq8w/cg5/432GDQq/e5kmV7vYY9266boLTE44jvey2Vr5YJY57BXW8fb9DQwc
xj7NLh5feca0JEr/niFE/BikeS0ZKKlLVwgspdZfe6GE6ldwKDcFlwsDAY5tYABO9MbIZfDaRckO
5jpqPChRfqaQS/+mhX5ulzPmmgwTk237lwweHk7dmQTv8Cuv3r9WmsxaYzZpffjT08iM6qTEHRC9
3PfEycDN2Y08DbI2fTak6zSVm/PbzwClQcEIw01nGb1evx2T/EpAMSP9rwG7E5WsLPJwbZi+fyfA
8fO12ouxrnrOTs5Kbzj/Tam3FQ27OeYdlda/W9lfO3xblkr5hn6GB/6S10VjOWOnXNBYXmAu7Pip
pI7lWOBHYWpPXZdLFzpXwYEp+zDJaTROU1Dff966zpvSrcYNl90O/PGbAjPuMMxDVp6W/YJ+hT8r
HBe7Fve/6DQWI2wA5aFqwbP+9aKQsOWCUQiKjs29FP/pWStoYk94qtmUeipdiciaeqTyEoh+gqUp
U8QkCRG7FPOyL0sMUYdwx3/JJTt+I0aCIbGMhxSzCr4x9Ms/l+Jpk9k4DGzcmIvpYJwRgIDec/Yi
fxbhO8jS1dLtlmw4oLjcbCuGY+qxvJvP/Fs0+iozzSRGF1VwnJ97T2TfaoArPMmh2IdwLXmvvkFf
gpsmdI9g507nJ628EcEBckwiHW7ghiW+acpvGr792jw86RMZtE7lBOUkc4eoUIfGsUnaTrVcBrkX
RYSVwZaWl96rQYlHsreydKZhkDaxjQnexjzvR2KDJmoz9exYFFAVKKeQRYCB4wUCAZbo7qbj1Lqx
0pPqkGwm6PQeeyM/vBIv+22L/73RuMTun50gKYETPGrAjZYGT5lxclioEb0rWpSXATDv4UPgUU9J
IkQTNUbdpysVs/7iuXirL+Ml48A1F0BADmJHrg1lA945ISSHcBkAmtb3BW6Hvuy9LhxAaunEY781
HLcKem1OgbMZ1gtTXRHDUfzQgMjGBEIudAp5BajZv0Hsdmj7qTLB9xsG7YlsOLnm04CH5isy9iHn
rHSOFrpuov0kJetRDU8+4958LKHqHAQNcEW0o+j4q9SniG4CxdtdC3tfX/Or1kaUMte7Myb02lLq
ucHdv8yEW8Ox4njQd/c9jQrQb9pcVnafDFmFHObWYPP/g3C5QmBPFCtmLxJmzxY1k/Jvrpe2SDkx
lfd95ceKiDCI2HJTVRX2CpXrzaX/4a8oR5cXxm7PkjV/TPloAxaNjKXbM138X1R1vYdK2OIkwvqo
et5OSeXuTafcHYX/O9G3AQDNYuee+aOLoxdF6zk65CHAjv1mUNkjvjdgu1QM6mAo1gdk1cW2e2PZ
KugjecGD6NBqWxQZ1Z89Hy18QXg5h4w9S7pKJ3KJeTinJC6v89NsJNP0NhzS7B7HtDaKX3/tQG4R
mKwcklfhI6BrmsZLe0j24Sz5kScsQT3rsdhk6rI3JmEjCbL3MdJEwJDIOp42sp7wfNzzBUTqaNg4
cVMuHqaqXrGl62DATTMn+LMqjaeRH4r+Dzz8gyG4pDSB8ijAXdpfc3mhLHzksLV2c3JA+BsaCssS
jmyYoF7G5nGbZXJw423VhA0H4qKYidrKKkDKufCf6gxBeWffXMMVSsU8LP/ZlFEBpYNItLhAzbf9
/jaYnInrQno3BxeoI9znGGZWdxSpvFScpOEvYaO+coMGwcHReuwtoTHktrLKr0ISTB+TC1Hj48xL
rkv6gvTDa4DBjpivSyn6SpzxpoRZXx4RP3SVmWYIcOAaOL+syEZ9ZIqdnqPVXMXR/ZBbU6kyrC0W
5CfIN0eLzRCEGGgXYMPt95CLQ5YSySvKMwgLjEq/R+GECvOkvvZ/0bpvrDzJP6Zbdd/LjycEyuYM
NCALK5Eiqze4ITOnhP/disFaWddVxkHPqXbot3A2B4uGblfvxateQ0pIzlQqkyoLN6yYD8pSdyr+
C7EJk6/bTWperU1qIEckibYANp3tO0kAegjynLmsbyo0Ix4dFyxOUwt5lp0zuYrIkeThpofcwi3i
SOUiLKFPkpSTmbZW64BMZZXSdXNrK2QL6nH8zJnj3JeZprBdzVWk1pLIBqVbPxMlLiCp/aCpb4hZ
V9d0N5tTDi2JvAFqN0l5PHquHI7xLSDsORAu2YA3w8WMfMKJ6FahSNT2pWYKLPRzl56TUfX1zpUG
N8/ZcFDHP0dBdE8qpWOTM6B69Yg6bkLaxcXAgAwHj4tXenFDTYtdCsAWmYlZYokvOMrBZ4vJpcIw
PW1XCVlQCU7edS9GVqijuZWLq55Eb+3+QQnxFWwjhiC2JB59gq1W+OZZwJYbkHTs1tMBy2db+4jV
NpSOm1MGTSGJhfDKyKVlvbdWAUOMNyaDNtui7GvouqBZ1cPftFCZIsubkHTijhvpdq36ZgUAbukx
oDXTyz5WMeVJDCQr+RjJ28Oofix03rETGIQedDX9YdyOYATTZqIVVL4ErKIu2/fRQgBteOg/FT+R
YfhCA/k3609L/CPkW0NusHvlsuUl+BC0Z7LvyTPuC2ScmsJqADwiIygoEf9DpbwNzqiiKKKV0iyM
LpPLJZtfUaPPVkGVq7GK06DLIrTzBK2Vs/HPVQaoneDmOFExFWICFW1GAWr39d8RG0dnY31p+5X8
/L2d1EcfQRvXJYh7SO+UCN+OCuu5PiujEU0JOWg+8UduGC4KbTAFeUwVJ3b0H2T8yqtL6BqouBxI
OShvYu2l1dCfnoog8zEfFIT8A2U9YZ834XYRY50Ip12vVet00w+c3U2m2eBz6XgGXyTATNf25f9/
J/UdB18fMqD9Pr5S8emYsKR7SDAaN5N6wY8uJJdiiY7J/ZUKoaVqXKOp4FP3eSLWmr0YPNv9MABT
J21dzNSXbBI94OawsJ+pBC9JhYHg4E/q04w5bNk/TXUeSQpD/akLRCIoCIlbVl57QjqwlTwahV+S
iQduDaGa8XYH6SFAnIhUDa9FkoHlgp6Ff+4zWmTLeSxgNvkQeGJN4RkH+Nedog23Zm0FJn7aI8PC
BuFzSjZ5qdHB6kKZTxZtE3K7pJhMI8Hud5iKpngZT2J22vfwNk1goP2ecRphmXp3r6ue0NPGR8KM
7DeRxvsGQI7Mjz9NbldSoqmmnlfIBzfp7gjKaCS5Le70vNg1cwv5BMY3WH0j4cBBYdVlrOQqCXX3
Xx9IWI8Jg32itcrxZ9eYxfQc550q26I4D1uzv/0yVNfh38BJ65agCfYnDK792+aW6tiHgAE3SRG2
dddcKozOC+aj3q/4nEeCylk21B4q4XOpzoK/yr9HZDrpWqDkJLZDmVZ6tUoNSkRbUpN71Ha/tWCZ
/fGhDJFCaE6oAdjotEOy22/0u1C+d8MoRFSYJCfcTzskM+jS2g4H5W6nilQj9n0bPw4qKvmbsnou
hvYPwhi0a0UnKgQI9atPWBp0uVCK1DF60EN2AhuIC22JIutGU5An1d7dhwenGVw5tKh/jk86o4UN
iNvkxgvST5k3ly8f418A4rRRJtihmSp9m30yBjT/vATdPL+4E04852sqKThvZ13Kv91nhL1vyQ4T
g0wJid2qpkVN+m4Du0YJpjf7zbV7ApALmz0TaJujqvT84i/8pkXdcjCYGxj+CwXJCD9fM63ytzFd
N1i300tcmiECmrPjGXyDibEG7UVe+wwy44vThpPShMyFsdcqO4fqqyi6xlt+HLlR6A8n9A93p8+7
lGlB5fs6Bsfq804YHvptJ4iSKDizKKCeKtLTus5qe9l7ynG9MIBLUCjQTyFWCzE2H6QR02uGXeyl
49POAxmZHo1TN7Yef6tuz62BpCO68Yc6WkptUZes/1woYMgAJht6zy0IEARXLIgxld5K47+ooXGH
/EwjDo3ZVlcE4fVUWA0Bpu9j0qyXRf8XKIBNkH3sS6JWL/o3DSivThXVwp60x7qkGi05o5TZOK7M
HP1PlrBVVOdkFn0AgyaRUjrMhmLZsw/im0ry0JvDeLWMpVKix3pjp8aIo4f68z9eP2BkzoQYE0vz
1G1jmwLXFvm4uNNVoMOvmgqDCFCtHk22wGvJXVUoPTshBzLjzHX7WNfdOLXc3miz6yDb7bg4w2Zg
XyeF3le40PZjMID90PaNVvQMFdnk7S5buJ23+Z7dAtzbWZe1O/5TWvCl8FPr0aqVn3byIMxAjUSq
L017QRc0WiaIYwsjAcOZqe/eDM+YxK41FbU5gVxYIzK75wqceCLkBtHyMGs9liJansKu9HW+Cxi9
GIybwpKB9OfKPq1l91d2KXVG6CEoj2436Rw/aAkvKBGeuOyooffAMitM0eWsX3z4uOEjk/WYBIio
AssgHMVtdi3jCc2Ym64SXK0DBCOHynTIvsjgZ4cnBS5EJ2sglo32yWKZPwdml1usPctZS9uf6lGq
j+AzdUpeNmVbrA6fqTHge/sItNosp6yecbF1tgt4sm8ClNmXslf+uqlY5LBFH44mpmnsOr3SMhu9
MeJjni4ggrwg67sdqEeJkTF4nMfpu+630i1ZEZzBoApPvbKZP9wHQIN9FJF2l0/Be0d3Q7bWxE5H
nTM4H3iIE5jTnJu6LxPzf1W41PtoCJWEHpOhaQm/gBucVWdiQKq4k1AQmdkqBCSAcdCaN/3S2oIJ
Oj3lC2M0g5SskDnjpGW99h4afuCvkQK5RDtQeFddtU04Wz9au+eXEziOXpz3f436G2intaoaI19X
Har7uVoEMCQMJPLVQTptsrdTyyNu0j0rsE1oulKaL9KyOiCdN6mkIafifKkU7CS9ijGr0CfZUYS1
6t+XowGhnZOiAL0Fhs1H9O2n3v8+l/a+kBNhBhuMSFt+2inIYp5FOoK/SDffYymRk/RFRuRBNLwo
BayYBniDUxNGQ/zPwXbexMv6zv7254jai5Jkvb98n1kejqJ2LVFtmCfmDgYKOj/t7V7EiHI9+1l3
rTtcR6oMhJjgVMzoLmHOPij4I+cDAvKrja+1Sjxpsv7Vl/+yyh/oXYq9duPp8n84kCFhvNQDaH/W
f0cQoQNzn6j7Lm1wDlmapJQSFQZKfnM0GXGfwh+If83rAT7uNzMEpSROAqnZZoz7XYtuq3/dTZas
OqRpe7Qs5KrlM9YryeFLNkakVmBktNJHqQAijoydsAqzsuHpbIsTkUSpf0Tql4YeuUl9e/ltud5R
UhndaTJB9Mit6ba015JU7l+aQyaFBjrYg3k1/8HS+wwnqXtJcuWPgJCv0Jc6hV6jDJSnsWVNnV2B
TnuGFp0J3otMlnFCatWanYNKDBW5TBcp2r1ZypKuk51HapaEA0X8LWA3CccwEToZHk8tO1OGNrEi
gP0bAZk+FzhI6xUB5ofPn4kTFi1IBBS9yI1S2bRealZZM0HBt7K5eQ1aS9H+dtbaaOBb+s5IYt2k
E7i8lpNstDNsqFx3wIu6gfWTuMu7crkqCkfJF96nIpCy/a70UpZEX7PuT8u03MbDaHB206IGDu8p
6HoqeR/Lu7uG5b6ePxjOzTrnhdJw6vQkT7g4ujBQknjVn0dLiz1VtwB3y0R9c+aOdhTCPWjbmPLg
GzSdrKluUW2G5+uPiLrO6uTH738922nFA2lN8psh3hdYD4GkuIcifxsxPuYe86YlQ8jdAuBkNXsZ
wYzKLF+N7SLKVda8B5JITinoiSv1gjNIqy6uetRm//ELdoAqWzQMapHhpYU7AWtAhZiy+v7PB0h1
bU6gUReGq2XsLL0lfaw/yq0wY/TtAy8kgLH+1LLPBlcxGLskfNE8OzqyIxUggemi9jruqrrhnewl
tAHTrpdz3Vf9R+Qgmj/0Ug8yyT0tYRpyCNBR4HAwlEE6wMxuYnFinDYkxWxUltzJ8vgSfkim43XS
rgIsq+4rKtT0cPXQg+2yUxT3DInonvOzZt/3KvQHZrY1Bh6/SCg4uv/fl9DLNm0xlLIHuUM+BPv1
muJKLRLJfdT1fchBIDYk+n0bkCHPzgjfcULS5JJ5N81Q0SrOt1LNCCWL2qp1i2Oa4DW00qsmU7rN
h2oj/UmSpeUy/x5p0rH/Y0mNEzako3rySlSdC/L0wmsO3i6j9uZo3xtMPj0Nl4ABcj7coSnPJ300
u/4EcwcHVuP2YVgFbvjTcsDs3coZJnXrIDLFQuzn3BVavtoDJfiZ1Xjaejh8TNLQOLXHBsclB3Qe
Usmdr73MAsGzbUN/SqLlu5ymfUvJ7xwtCUqEWvkeaGBosfCbdX89pAfGy/O1T1xwfOWm+0H/gg2b
DTXlWCuIpvaBBonkT9Rbru+G2/GHwWQOMhgi0z19+x7sOXTCGUh20DnLp0hJiMxgVw76MD0cworu
Qx56zNw6OJI3tEaOi9LlQMzXxMHNFdWoJpgpS6NDZCNiWZ3oiLCVPR8AUeyE6GNm9IWPSaN9Mx73
gdPHCVmOrwK7vk1CpJKhHCXbzALdojonGlNj56C1DtBmNccNuuVUIk8JlBO0a75xk+jvXTVQUSLU
lAvkZPwVdtouflprb1Be6GwjYLyz3osfCO5xmHZmQVoCxayCKqWM4Gq33CwFd7UivYkSRw2Yfnu/
7PvOAvTDnjuIkcbdelSL4EYmsxJNtIRcyOhbethJk5JDaLmclOkof+E0NbO69dKBT3GAQhNOwRGn
f+ic+49/ZLf+k68bhQ+PgXsPZ+IIG4myQD/tgFP35P70+wvELNTdwMyPL1UaSch1fVHONDbNrxZO
mkaBlEd3hNgiS3Y5hF2orXQIAs3T0faCpqy1P6guOfj7DkmN2kqUKIvuYdYIDW5Vq/65I60pCLHW
85KDm9lcSTEAF4K8Zor0kCftjMKzhdcrnUedcOlVqnU0OQ/4sEt/YSm6X8JkLY4YZtjobI8JClnA
0JhBVMxatzLKIdLKo4Xxp9DZXet2/3xxZmVLanAIQZ5+uTBybOA5kXGog/wCHQWMVWdez3T06Zsp
bTBoF4E3T4ACgUHtdcFCatb/BF7eYJXTwCS/qeeL9OQbRGeq6zxx08+4EnjQqPErUA2RaAIaN8ih
7i+QllFNzCJ+qWsqQzVvcTPPlzyZ+oXjNwovm9Ujgwx+orjO8a1yhOllzCYP4ypO9PF864fzxzL6
sxMHVcwsyV4j0nccQLL/CbEL7xMt4kuHxjFrq8fd8ZxEKuwIUUHSfDqNT3kHmnsW84Kd3zKOBQ+m
lc9NlkbSa5wxY7PU9JhgNXlWnTXTGShke/tUoNhPQG2y5zjjQgIl4D1L5N5Og5kBlvJL7gBYtNfV
ayt1173XRRNM+5pxMKSAchUi36wu8/v7oJJCjbiNNLEhqNrebNUZOwanydJbn0flvgTTzao137qN
e0g0DKsvUKGEHVX1UavCXvmScvw9tR+DiUMaQm6CchwDl4R/JtR8sxVdr5FQOXTnXst45Tx4yEFC
KJSG8fFWXETfOgCmZ2adaGt2MNGDF5auNRYMAqbCVFzNoeDwI9QFFserMvwfskm8cd0IN/lKs3aB
QAx413AIu9sTcwmkJvWk7NobGmoaJsCOZlI7ua7QfFHDL+mRJ2RqxKraCSL+i9qNCH7myPLA+O37
5S5R77jHdjo9c5l0MSI3D/F2oOAP8+kg5QNmRrv8+UeBfSsrlqGsVtz//CP2MXdDWIPNkXrV8r4L
I6iyza725bYoakyXfYPsqCxyWTwoVAvRvJLo9aMIfvBDfJKoAgVKjtwcsmRv74XD223PR/5kgEmX
3bkB0F41RWH/cD/o/0ldhQ18Reckp7TSKMhgrnz0d5UCrGIeOp6DcFbZSYr4+RTULbcS8SrystQV
r0PBukfSrxnuw1XFO2fIXk2DtU0lWnxHyGkUkYFQow6+EIq+R+nhsph8ZYzfoBYy7j8qjoSwN0pD
UYi9giyCMR1UtsIu/yU+jWyVY3DYqv1H/wgaDV5eyhA8HT/7rkMJV+muxkBx4lJI82iChcDwclJq
+YqLv6i1PcpYZNTDZAYXnc+IHRZpFyvU4uyqt666dbx9+EUcnHoHGfGBm63vxCfrCo2xjOETrfc5
5heqnU4f/l+SDYxAm5fP7qFQti1b2NCn5Tgpg21uXrgrC2+nysboL+Tgb2mBrxCunR3BwtXd1obV
jWJh1o5GKiLXXWZcUkfxE4EtFRhGLZMTmq/sTOIC36X4Gk8kwBAIw97Zkgx8FgyCOTLBWiBuuKPY
xSX9/y6hHfZnMIhLg1fa77VoRZrGQdOh0nUCDNZ1+fLp/ZsaeSLe4Wrtjhi42l3ASXZFUNh/MZXx
BjEC6S4Y/xhPAEJsaPmRTeIDLmwNrontKeaspnMYzk/q07tIlGCLy6StQL9ipIFYud+BLiJN500O
Ua85I9DhgTuLIIJuMWUeagG6apNc9gSISPKIthL9QJBnftaHgCAsQE8g+URsu+BxHcgH7wgxvKpO
uQOAD7U2nUFt7a1nTpVQY9dEbhUL9MbN6CESkU53J7LFwUK6Tr9gPcZFDe3Enm7niifye0bJqW3c
4ndKcqm/A6cNXKhRCZvcLFsi9v4nJKJmI0eCyel6VwBDw/8eeEGWRCPIAoJ9NmOd5LMiFMUAQGIq
puTqr8ZqaJgCWuJtmuOJfgg5d3bf/UijT26R5Fw4ykvmVs3RGnLv7qGXnkLf16dEeFJ1IYfX3dhP
LljSfgQxR9g//OxFgs5U1SYDblBD5UeTYxfeWuXPIczxDZThTWvo3dzsbyASjOtbTRUx5SFDuW+y
NkqZ19syb011kMQLBxxjFROOwOco3gFdTXkgk2VRln4xBFsPF1jg8l0Xvh3I4Wy99S8W2ks3Y8n2
92/gyrU1kjX7uSGF1ZFHl9+iot2Y7kG6wMDgWnDHyT3ME+qoLu8CMsFYtfglTkvYqQlM82StR6qA
jLCU0u5VZhlc3t02L5RjEmBG+mZrKPdC8L3j/o4TEH75vGzZwO0/8OSAtppwxKDaFxw/bO/laHD0
+kZPH2NLonK1WGaWuFI7n7hH8nPeY1jh54Vgm8BH4Pr/JzqYiLkHnsZW5wT7JoRVgHQZFffo6gOl
4E0z9yI6aBxUNXxdCzwfK1EdPR1zJ6ArwQa4rTTRy8Btnfsmn7TONJ+VOgI2x2P5G7XRMTHrActi
MSq6r5+fUSbjmjw/Gv/ReylLDogYuQG7QLFvsaKrta+LXcN/NR52yR5SYIyv+nr3cZJv9bTE2KEC
I1K8DQDCc0A/+ry6BgQ4PeWYGm2+2Tqgdw0XfDqcF4pIC5giO3xRxsNKRjuSxoSVqRMhQRUAN7pZ
Jrn7JcHAUTsdpbNbmEHhkciP9UQMMHc5U3KTwpiKg9L4SE9eJcT8EwZCDzjOJ418tQOlCLHrteDe
ZWYN0hIrHt1T5+FF7rHGCOiWYMWv1FzEQDrdCvZ7XucT42VW4Y4+Dl+DqVkRBXt3c0MQxqg8zTIO
3Nm8xifx5n+SA8CgAnEKJg7vRnrQqOY8NbDzZ/pHrjdZHU3fHK2PGf+BpDy1TGEAaCQYWnzCDGv5
LIOp1estNLOkekeP+QMR4H3EkrwjY8GgEyX0aGAzpFLRXGUt9CHhKRwWvLa6Y/jgQ8fjb7ItpJOI
68EJT6qC1MCAorWaFcHpzq5siurBLsyjLeTUWzNcBNpGYubl6d/1FIZKlJ6C6j44s6mLxxZ9C+J8
5GDcwho3erzZaeJi9I5YTP9Lb+t0H3yDGZrntEoiE7yWDC6EQmkppbENLReIejQ633oXrCf7wIDM
A1hAyCYBKCmYlh5PmSuchNebr09n64CW79APLoHFlRWGdKOFu6sIGRN0N5HXl/hiq/5zL2iUT61l
+LpvFw8kYGiMQKag46tfSojOiZkkVBNDp+JYTFnynrqG2kgvWOJfSNUHeuzFKbKe7Fmqgd76Bu4R
d50IQj8lvEez/OOY60vo+l5P+8O5Dg7RmOak04GBP5iisJrMj8R3zq44JK68ULv+pSmvamDsER17
TYRadXxv5oyEN+LBgt2yR2ywBZxA3U4AwzJZNJPeVLhBhmt2wYWor5f0Zj9pz+IWJbfoz0biIIHn
i2YUc4iHUOZnUkCJojWWlFM5meBpis1iJQTBI8mSvuZmOBbhpeVZIgVomcf8aKpejNvhX11x4Mw+
N0IFX3vh98juGHJpf9mU9YFxEc04Q1GxA5fl8exVbk/Jcdx0vbz8hmSRcRCbnnfDsB/k0QoB3nps
DVXaCn8qWKX0tah5akMOSVnE8n8IPRnKUD+y4STJGydfIi0Cu+Spk4AmX69rT/zWlcMm7or7/i+d
jOsFBHCJ07WishniLrgAa0FSeyU9gDYbjfNatG3znVE2GLquND/eJPtIKsXVY8U7+yWpIExIXsIX
aKk3DuRoHGyQAi9u1D0HmoJOzqR+nrDEsvhUlv7ipGBLoKTxTYtHRhkAgCFF+qFej18RsqkCrTmn
dC7LDVEAWoh+W1j3iM/i8Aa26wSBfy7ruaw2qyT4spZmQewGrFvic6tzFVpJQvSpvaN1f8bKu3fK
XEa5bONrHVfSUjuFQDDcZ5N9KaN6hJu9uyG5UXlAeNwkFqma0/dziiQ3VFCnQsQB9NGZ3HiOdehp
FaqQGMKZg2OTA2rI/AE/1BbB8AEHbww3geIaBaId8r2w0v+VUtVpn4uFhEWDoOE46znGtr0rgyEP
g7eFYETPRqBjRNUyBDHJ9UhvyeXfBIv1RsNOioFnf+eI09aDr0YEFevnl/wO8TrjjioRqkN2Miy6
/p8YyEy2miDzMAKmqbaQOHOWwN87tt6s93IflXFUjdc6MDSxenJupQ+Y84PUHhpD7KHLkvYs0FVi
E/GbKb9Hiunyv1V0Wa83sD/D1G3lYOzzJhSoJ7JecIoDGWRbGK9pQnSmbT+uOSPH4HcYqROnKATI
S6ahWpeleahUBO3u4jz0eA0QZPlOkmxxeWEwfYjWfOsay2HHE/cjN1a8XNRNpshRxZf3uZ8XmfbT
zU7YBtdn/+pkTNDsA0tExUOKTkvKj0LqweQQte91JjcQO6/mY/1VdI6IlI3nOxmM3P203Tcc7MlT
eD9sDClhx/PP9LMJsf+ffkiBv9vplkyPIbQdFpxMnBU+xScgOXyC1RuI3pMo5Gk295xrwK74tdvs
SA/a+itkeJYI+6IfXpaFdCtwxVqq5l5PBjJ+SMdMiX/eltpsWTOpChrJf3FX4Z7QM5/o2Q/dqbXX
zLbvEAlAjPh/gugrAwnha4CXz+OvWkHux9oFIaXh0RlcAiZkMAIOlNCQpQ2bkPA5zqC6zEXKNTdj
bN04iunqrN3+Gq0Mb/5tSrmjv8n4ipsHc3OIqgtedFzPvdxI/gsKOwBWK5PEq5cV/wxou2gOVVgx
8jVLNyPm5qD7OzJi7AHnQ6MB6mVz5P1ZwyPXFp7v6K73qLsTlui/M/rVDSpr4DlvJsChi706sHg9
yZy8BudxshJeCdilWAXaN6pD4eJd0ecqImnuBB5UMtgW+HOdeFUn98SV08Wg220DwdapGqQQwLny
r89f454txIirnlSdIrt4PjUJG23VRXcvZDKEZlEWsKGX+kXtjjf0eMvdUL8Vbt9K+wUQCFlo24Xm
UzQ/I3yNEyI54pgTTrKVM0/jDqxjrQNiS0syHxWbEqUJHg5vjQwFv+h5zon/c9PIAYobB9YaQX3y
FBvg5/JNBG5IbzLcDPm2S8uaJlANLw45dLWmlrwuixZYfNoyiUGNTCVRiL3ziBHUH64XK1hN+amM
TAyuXyzGEw7NaGxvRZHRmPfWQZJEx0AytOn/BMCTPYnLyalsGvyngAc9PXQb8+X/3K5APwiJPS4T
d78pnfut2h8FVxBnw74lF9U7iODRslfiJmK8xvWSUX54D8uOeZMDcqz6vWmEPX7iruDMQoL43EXl
tmPBcSexsl43t7pTm/a8aMaJY2asL+ir03QIP0xzGx6xubzi0OAVjsUe+L4wT5qZKIrOgDS2dxVQ
23cEW+nkbBKZp0CJSZUoErsBXbBVheH2MrKEB1a+G/jn46juAZvG10CdUuanJg/szhCMf3AuQEsH
wxfexiWdq8GhuGdapcSZIMRqVq6HN+gyjpNi81SkkPU58uKBiUHd9aooM5BWysyCNrdUb36fwdNn
EC7hgb9o6hppp9dG8wfCQBGAflJj+xLfakrZAqvab34kFzyKIhg3GDoi3VGbTD8ppW9qYy8YvR3/
X8FWKxZ2UiSjOyCxEtCe5GTnTT6VaVuc2KDPqZGc8g51U2nvHen38TFeaes97mbs/IMKIjEfqqr2
2Hp7OjctPmDlMfgi3YwaLbuYzAfQ3gFjgrZc6EzUIbRfEC4liqFITXj+As7PF1e2JPyDEDib0Crb
CY1b0E/g/NQp5SwUGiGnByZ2Fs6xQ1KSoPJ2y3n7OCDocAn9JHnvoHaskBqou9OFCbLmhjhR+MNR
D7CsX/+X4LLOhuRseSOaIOeCUlZtZzCaZi6Yq97Av1iaaf3WMV9WWQI8QMJiObSfdixage75IflF
IjxlehFz6KTAgWichb8XBYt9Dq/mB7orWYrKzxN6WykjaVNiK7cMbZidU1ln5YNPPMV3OdTk9rOW
jszxOLvigT0iRaLKnpKb59O5hJXvf5PA4qy++NM0z/snz/tcnyUNM4dRTvUhqqa23tg8BZ4dKvuz
DzdQLSS4E9uqJ1CvHyuXxjWTeX1hMCRzpBg0ie/hJ4yuqhxIqrwyojNeVpdjMWglksI/0Ym/n+pn
IgtZeqP7t484ydZAeUjAA+KsvVGZtSxCA0qE3AaILvSvbVDyi49cakuRYkyphbYr3s/v/tZ4q6z9
6/OCxrmoK8KRy7JXsNvTFwpK6wnJRkPeMwWEDvMboqnh4nrCKjEsz/AeNpnbkzmSmWkqAoWdIx8M
0CH7+scvAMRDGYCJH9sir+4ToW4LqRAk5xgBNYFqkBKh7IHMp9zQXWO8/E+9uiftDAZtYajKneSC
YVtE7MfNsMA7aer5vbe0Jgp64JnBn3gKflRiXGI22zSsCYgnM3eQGCepKDiuBKtAVjRWTCw+p4GQ
s5Kyqv+1mmqy0FOO9cr6vecqLgp5+Y0fWGi2i+EQwHlEaQ4KhTrdgeGDaJJvmuZAFXGHzBCbNAtJ
KVtbIGjByZozAOjfm0ZaXZzqvizVE1DDpTZ73I0tVmiCHXhQmGm2qDOoX+gSbhN+Vxa+opJsmZ+E
t0PnZ9chUVJrbPHQTvk1n8qTXGWDE99sC11Q01SpAhl2bifKZEcp7EBtN32TQshzC/ydreLk+C1r
+fqJO++m8AMXxlx/QqtNFK6TJhk7bJGmTxDXEpQeNOut/PZrNHMVpqPWfs26LY8U6Z2roORw0pY9
PX0a7sRyFB8jYcCGw+n+wc/EFRWPBluq6/Kp+7uPALxuK7ciCLABwpL1S5ykL8JPrrbyCNULbWpE
Ob6ArwW4PpnlM4etzb/MFdtEsxYC16Nle8M8z001jX87X2rjfMDkzVNaWzWDymDhrjzP4Aqr+d4C
8pMSV+gFZq1rPURlHALG7pBX7rdShBF8UZwGxiHdQbx3NzLl1EBhKQtVrN7fRGxcreM8BJwOlCPM
0SmGkE/VtuVcPaHbME8kRjrSxzTIl4knCtRGjtnPJZWOMynNVB1fFKd3XQ1a1kWiNWeqUCJsovJw
WtjeqcNj/wq/6Tj9E971JQKIDai4nqasRVrQo9gSTpFnV/pC4tIltT2v/rBYBMHkrxS00/VVbfhu
vF8PPTh1unnwwJSDeSoiQtIBv9YCMQUlVIBy9U9zUUIko4fG9y7Q1QZsdPe4xMmDudu6irBERQhq
UyhiaymMa8slLs/LHg6hGLDGMV0sYbqT9ehGN9PyjHi0yDsk8g4LG/040gsRaxzfy0a5GgTj2P6X
uF7xJ4vGpj8qtViC3T1+FJP0trxfM+Ua6YlG1x+o9G0KCOJwB8HWobAyh0XMyf/U3kmFlHuu2yaP
Shym3gUOvb5sJ6OL8WiIzV056LL+ehA1K2ggC8Dk3fGUVF1idl7QIN+Uk9qi+aD4xUyZ0X0XjXqv
mFn4MPs9l+vUC9k1S2YVNf+c5enbZMY6xNU7WQZN4v6R3AFoZulZ4YQvbMEr3mBfv3eeeQjqcAGS
2+dKLPqPmbFvafRQGYsj/ycJGLh7vHJzxbxpXPnR6YN0l0Tr5qJjQWRaTg/qZ1kL+GdFSGh4Gel8
HvhmGl0mwyFRr/2hKlPKK8/LcMteNU3cQ0K8+ZtndCPtfNgReq3+4Un7j88tfQwhOA4tHNFUMZJh
U2YDwW4MrY5poZUvKYoioGrkLDH+Q+TdffrceUcpHsPbmNFyhAxG6K7Ew018p3ZkcjmjITvxicpd
uE0VT0MG9u/MufZBnRepBaQJg/zjJSJotJa/h0jNj1C8f9gxGncvzdzNYQWUQC0OKhG5LXWvG6xN
sNAphxV0emGRwlKltTsAEioN/ayuSmZqH4OoN0qxeFOmrtYqlCVi3yU+Z1reEdY7L9L0teseZIR/
04D2job3zdtQcgTLPoD/zMT0rkFDphFLhxFBT10SxmxY1OjE7jCY/5mmPNfnKh0f2+Ky3JVFUlqI
AIADLIqHtZbUdSb2YtCt0PqH455k7+bku5ly7rgav1a37dcQN7ojR74oFJCW2awz9WTX6mI+gpeV
YHfXaonDGFZt9XTbZ/JTXRrDzk7ZTdgBYzFvbsP92t9qhN2rNZfxi+eGI34fC0CBvxdgBJ8tGE5w
Iw5SlJZVHjAPN9RBI6R4rL12+REoqJetIzRWJsvUThDa0T03QklgnHejnixiKRPKjbbeFEOUhsUT
CA2v8hwA0T3gIoNVAhHR+Qv34I6rTmZ05aO0dhUJf4SJ6bFZGuYhaDg12jf0dIor/E2U7HwI1b61
pUqZpRsV7wXl8EL6XrMGnmHAzb3U34jeZPL/bBPY33/7Gj5aeDhwd4GQimHVmNRDYhlf1HOEmqZI
bpfBVsQ5OVwMmnpcJeRTWV62vCfTHmceJkQWYrJ3HU6d1Bx7008O/kudrB7jnQGEYaCNiH0Jgq9+
8FdjvdLQWFJiT3jCkCs9yxGNlGwkwB10dRVG6+5jiLUGrBwVjD+WKWmvzmoNqx9zTRfLUtRnhQT0
UgYRWYyWDDflSazJXMfzrfHBTjh9ip/mJIUbBEjXy1sPXlhH4GgINx8CARjuyWYtNX73nSEP8MIo
hX2VwMtoMrnf85naEflnBcTRvWdsenBfMc+dtPWisJXVrDyZkeABFYfL4lQMQcGjZ8X4G+XuTAqn
tis8FTbNjOku0B3IYwMOqvk23f8kpv/y+zATlZXzUERv2d4pxGG/VJpUvoUrhpXFXzydg0KDFqtQ
3WeOE95B4WkwyCY3gnA+uVV+ttjjiOUL6uhy2rufSnDhclOWCao7MInMRMvqaYl5Bxmrx8Zl/mpJ
kGLfTABXOoyfwnyjPZFhABuuliCOCZ/l2ekR9ItEvWqi7+iuCbkfLCieOx1icBr/ehm0JbLGdsbJ
YerTriFu0BrkUVi8Gb1Il6ks/R4HHpUf9DZ4Caa+VZvSsHGGkWOfh2GibyEWIDrcHQFzrP7DDG8j
VhfI+vvMYisTsNWKNtoJz2NlAtXSGru6bInyaNlgC3q0QMkNDHJ3Y1COLRW6quF6avfTcFB6xMfm
ZYBqJ7PCJ0KqklUyWleaTjddmuPMOU2NKfNF7dLXoBYhD0XYm3PWZLR/cJCNzZcYz8iNtrg2OMeO
o8EcVeCTyUi9u8p8l3gtZsjk6xo8k4C+RnP//1uR8o6fzkRuAEKV2Q7MpqB5WPQtce1RnJSDJhoQ
ZFxOzVIpIk9VyJu/vWNOoV4wKEGiqGTIdGvsjU5HPULDQcIfWpxGlujpeFJDfeO7aHqCv9gW5idn
OZSotqUDfZTTxqfO5Ddt/zmtdEiEmdfCg1+bayCwDFNfpSiu4qk1xkO/AwXhtKsLZ0yjnABYYiEQ
iZ5k04DakuifCgMIPdY6IhtpZhQE8y/ev9uGtUyXkFierct/bsUkhCb812DUG9RtiyF5r+1CEIWO
jCfW0uNvzWuVFkziNQIYUEgun8W3Lz9SQgzw2k1AXOWfB/IdBDOlwaNZtATxMquKvqQLTDqGMRgw
mi6AxYqfVbQ505jeHartTKgvc/boawWIRclFSCJ0ZdJI9LRxsEPulEBtqiVJwf/zWqi0WcwYFm8y
mYcjL9nr5awwcFX1J4JjlnD5ZIeODL1asjwzN7Dys7cPJoHqU9FwgwOG3FNj66CUAxF/6T0EQowf
1E7ISS3sh+YiO/C5tOAcz4LCrJK5dNMYaYm3f7KZGlqid7Pn1Y/9oYvcBG6R29/IfG4sVvIcd9m8
GIz/28eZ0fMpXLf1zJfyKyYQWRmRPnwdJSyRKHFVxRlh+vdAdEyF03YFFUvFdQFifO2J2H/VeiGR
6bgm3bK0iVyA3BH/5GvNMWv7je84nfQUvxGwFKeuiO7iZm6OLboqSt1D/C7keXXZgdQtpr7ZYg/M
g17WV7/F1362gnlnqVLPNeAxr2UiAdGpp3t225C7Vy7bxsEsYqLdq7JbWMEiojcUD2VysMn2+wXH
gc30Y1egNcdoKUfyuEActefgjnpWelz615pwPY44CJNFsgerx2soE3nUS9FtVG72Ab7z8v6jolYu
HSePGqa8iBz0/27+LvHx4o61Et6ESBscyvT222qs/M6oVO6ANn10PNTiYHtHyOhg2mGMOn69Xu6D
fJl+TBR3okJCHcJqAtLVbyti6VL06OW5zkTznEBoQYqwkLUFOD6KhmsHbnCvj5rTyGUxF+S8slup
cES8mifxdMILNjqxGWJnVyQ6IniOUKAU7LBJp+OtZ5s/SRxAYGLv22pMYW2Ub/sGEE6qrSJPgvBc
w8zIhcIhZIPhkoUEVEWkD4UUCIp3+tMi4Mol8fmk86uaCIxyvrv5YJAbq+AEZ/luhXWVDY3HLMMX
14Rzk/PxYu2Q8J3Gn6qIXb8fFklNh0hNngkGQlEiyck49h+PxLtSK1LqK3lZ1A2z7EbJyUTG+xWr
bB0swFh6HAoPxYJSmxIoMSuL6+wYTYwHsQ0K72Z56iCkUCV7w4a9H9Xx+IUXtPqfrVxtvWnXMwbi
FrgtF1y/ldQ/6wBWoAGkP75P9oPbYZnAfa4+/Y/eQTI2ngHd8/UICNDnRXv9N+fsQcwVwJKyV+7l
ytNvWFrot7gzkw4tzSS5x6UAjXcTmEcK03o/fBjD3BFS2bw8uJmQibUBTuZ0izivkdBulBSokOiT
325KYEj+Zj8psQn4ER1eGAeQB7rC+fuW/SXeNf/IkCg8Kr9YxcfPJY6worotFbR8+2QL3SDZhYpy
p94ApJ3g53YVnoa7SWlV23IDqN9kfdrFce0LD3KMgRNzI39RT0qrs+1Ze5zWgIw0iOHU11gzDGB8
+HvkH4uUeY7qBJUAQoTU4Ii8jB+Pdx6qMg0hRy9UaF+PDcGbfnxuBLba2IlJ+5fnrRgPSK4gH1zc
UuEsacP3e1MBmAF6bYBNVwA7h3lCgyJqQUxW8rJwKeqPU4lboAr9QWUp6WT4WMkpifxWs1A2/nOK
9HVpfWxIv56TbuXNOVgJxEsU0/exrQ1GLXE70EabkEO9vo8/UUequkPtkvyBmHn+cvcDVh/6mCC/
i64QUq9Q8fpG/jW7ZGwVXBX4z2Sz2c++mvA0iZVviTO8iNgh+yW+ms+zq3rKChpmNUZ0b45AU3rh
AMijLX6/cwLHOzoV3xM14lcI8b2xUU5pml2TphFAkQ6ScIZuvChDTOft5hUQxrQ1+rBRSbrUNUEc
7ktj8s6kvyswR6KjV4UFrCr8YYWE+fGW+RgVVPw7kkWMBKTX8RQxVR5P3MnRSBqY4z/tKCYjcYFT
i1jTOxlGUDYYcP9y4JnXqoN08XFnqFcxisyjR376kYCnj1JfF7ZdpMzRn7eGgYOKuzI7Jw0nh5OS
ImqWaJSlvPxT/6H1pDBVCy0ShDLxr8EjLtDP/A8weR4ZqyielwlX+E0O3lsTaJ1Nf2fKZk8cLTgE
FMwc6boay+pL2nPTMGyXoPz/SBW6U8O+68fN6Ik00ZVbKEj1m5yDKeQitG3661KzY4HzTZ+g0gnI
7J0OSKar28yLkuD0qkcgBgx36aAXa9y0wtl5DLThqY8v99MhrnkkAjGextjO5xRnx7aSJSTMQVwa
wiNQuzD65hd0o+90A4ai9oVfriQyejHyE/tBCofQ8I4pP449afQy0V16Lkq6gmSaC1wF02gZ33xL
h0THZk70q7yXjFjAkgl20HKtFxIJekOJywAq+hpnqt3falcEKGFit9syCeSHq16FwCGe6wl3IGez
LF1Py1Hs71bTXh9YJNrxprdRcvCS6/vxY5FIv+RhqAcEkezuP+KvRbbp+xUbE5kzy4CuIEd8Wvnj
gEljhzR5w946dgfn/uPcWLNxWFvll5UuPdTKGv62XVngbwcn1oLAClcvX/eX9yaLP4+qnppJ+6+B
cZHBeWr0n8VRe2ciO3an7mM9dBXI+kedAajGCnTwZXM8XtWjNvwyxf2+BZTVPKWE4ve92st5kmDt
oR34u4OEDe7GezXi1Lxy/1Jt9G0bLodBTV73iBy5E2zd7xQmrTLwQ1kNaAjPdRUuUpoA1rbc7ASq
eU7g8LgteSmuExidBKY2iPVTgc/+pABRUseVzSUu0BLQkmEtntnB5kfaemanQ2v5YVABjIlJQnyx
1QvvnPM7Uuq6cdXx1xTCjqQM+pwF1CjgNJ5z6p+V+SKDbS0NdOGJVGX2FZGSp2kJRx+6SbwwlbXc
aL0fImL23GkWaX5mq+m/oDCpxU/HfyVkI9KTylGEKmgNBk1cOWwhHPgSExsjkFEbERxYQLRxOLog
d31Mt4QFyuacTiPOvZL2xlcvhC/r03OKeTMKmdHmZlSfhgCyTZPr0OmkRjvWhcRaEXppeHob2tg1
YKIXN6jFCgsw9KQadutvj4UaOtCfg1BCLExIWVN/HRIgqZNGnG/m+w9tj2UuK3wnfnMFgsOUiQHT
gXkdRBThhXaArLDkbA1mwE66BV2rus7n3R05p81SNJNkUftLcuIT6bnc6fEvJM/pkPhJhx7lxa9A
4wEvpIoR+cIAtKlio7SCxzfa8c7IpFNQzPTn0MpdQyR9koBHHO6Z1Vl4kK2h+YgDPa0XcATHiI/3
HIvb4nmWBojYokxjMuZwLVwDpC8YUeN2EfeShFzdIW3ySqx4Py6v/EjkmhmDlvxaMrAOQPW0fVud
X8nwGYGyNDiCvjYX5C93anU9lWOQKElA1H22UMkXZcrDLWxo08nHiOmtG3OCg3OgrxliHze0lnCG
hT6xEiUxaagoJRox6YQwsV6Bm7qtv68I3VIxn1nVnJllb0gAuH3fXV9A0fql0WmHx4gwEY732tzp
1QfNtrbAUC4Wp+6MfbGmARzpgxY8y3ee3dOvnkvX0PLQVyQ3EDSari4I/C+s+iCDPtpx8TnIDSHH
mA9K5ly8kuJbYbVprJFExY+mQ6fNaPVMP7NWrs/upydZ8lKt14UQIc4nt1ePOY430iGkyassvRr4
aJLqqY5g0z05/k7CPeprtNCPtsTxkglT32t4PHrz9YYw2G7ctWqLnWWcuJ4kLI+z2GB3ukV8hzOe
QlGjhBHK2dKwOG9KeUO0uvOloPZJWS10yCMHrtz6j0TdGjfe7YPQIoVHmKrDIEHOZXUVwUqrTCC6
HtOwMQsYI4tsOzclKXRTFCLstFEvqd9XfYrI8189Y49sYLNo61j/ogG0vi6iXGsPjFQZD0bI8iNM
7ESgV0YUz7J0Hm9kyaOSjmNWRDxTRzGscKu/7xysDv6Xk4p0u7MUVX6Rt6aGaT2uyH9GZzu0XS0A
nluFYAdsHztL81MTZ7SysE+wgjd7qadaItjFs7uTQb1ztTcck8k7LwPrI+Z95Tq9SWRsNJ68FPV+
GBf0BM6zDHs/Wzw8d9brgR1He2GPg0DtxFeX0kLaC70a33uyeFLinRWZj3MouwRdXSuXfziARqkY
IThasb9+yJ7o4laFBNu4ui37SknkrbzvP5S4maS+xnGcg9EscksFqO6cDFK41rO7Z/3SATPMTgeo
pWsq8tPgil2c4cj8r/k4X/nwzAS8hH11UHDECp8xRNCOvRCeHaZdx4k3OkuegPytKNYM2VuZRZ7U
30d9hlt87il+C65nzDuizflL0L9aR5FmqzwZsEyNN5thLejRdWeWw0UxrwqfrNre32IPm7oDK9Zx
lg6+XvSLW37DZL0/4ubioVZC7PV88a3hFe6nobL2RPfWdhoK3hR2le5ET/J5CU/UELSI+YPbBg8e
BUIueesyJC0dx52jP79xfF4l7W3qCNCpBJkfL1KMhycr768cUBQ5twlYEallLdfqP0UJ+1GouRQH
CEnD8sAgAbPhU+NJeU24lhXmxVfTs7q9gOrVn945QDn8BPRAgZDYt5UTVaY9ZmPt/hcQQxOg0PI/
/s/G9RdXF4PSa+Xjd2jHztRVB2qT4wbOfR78x3UNUW2VXnTlDflfO8Ml1QtPrDVbXDNSnZjHzIuK
AnZd6Kt92cCAbxFIKJmnkehMeLxMFGOPDdiQE1LOIXkwTvGO1TaVAdzup1VJphbcZPjKFsXNEQRe
Pk7SDmsvtkrsk1YaDlBsti3XWUhKo8Lx7MSFPBs50ac4LUPp6LPXXqi7LHwH/8J6VJLZnn//8Xzy
8yH+qZv03gnYFbHwzGoD5j8f3zb1lEb2PbZHW7m8O+B2k8aI3Vn0eDRjF4+gcQOSv9uYzMrkCsUN
yQnZjz6oLFRA94uPCbXI9uBdkd9hIeX/KnzfzEEVUt3SAFUJedbPq1Fk0yxQLf99jpRMAgwSsgRW
KYsNLiYD74vE5vID8zsnslD1JTdQ5mUUdyEpTu8pWHjiSIIcwJnHx1PqPMeoE+q2stwcDHXsAhaT
3AzBKdG/o+i7ZM3VNH7AW22EqkoTJHD2b1jxXOXhtC8zAtrH8UqmHs96UzXYRzhbYWe3a7GZetvO
kF6hRzcUCG2j+1Hp+HDNbeJrEU2B+862xUly+fndCz3C2ECgATZNQ231NTZq6amozjN4v2ZSji2b
bR8UAiJB5NqI+8AhALwfgSq2Vn3Tl0hq4SM+9VErjchvkbDIf/MRMI+U8UGYZsN+gb1vAG3SKh5c
gm+ZZzIS2UQuPO5ZoUYFxlyi+a7POMDMK9bqFoNyEMZshiuH3uB4b4g87wGnv8trKTz5pADMqZNi
rs8aSkINaNWpaS0fzTDQTV2wHSgIMFo1BLfyeuhi3LV/CWM7UzD0fjyg5fQv+baJQVY4Hgscxn+l
ks5RLoguISHLz/Lq68UmEwVvfQVq0BYoyELkjC77/esD6AJKbCWClOhpU4IxEGouU8Wr8mSNFwZx
IXI+uHcekH+3SjyEZMv/YVWB7CD7qxjL48w4VpzFIYcYsau4JW5VeaHIW/XlodWhVc4Y+t5brsh2
3JNuyqMUsajFDHg2X6mr7ZmmL0cs9hAcVw416Csd2V2DzWf/a410H+A/JZjmbttWv+LUajLwogpx
Xf201B8fzD3kVdrW0QIYe+QmkDo96OdQ78OF/ohGikXem+x/r136izm9X8e2aa34zujcPnOKA52U
O8G146jzRYhdGT8FJ+C6L29x8uCKzCmfSf5TKz4JubdbnRFKcWVyYgK/1OCi172VjUhtxmXVrZaA
ULIHV85s3qCBe0YGZLFs0/ccju6OafEtm3pK+5V/Byb3v6CJMi7u9x/qT9eMFMqCWb1dKNIC4hjw
uOCZv8ZerryYqSyVHTnqifSVSwQ9NjMC8o8dA329aDLaor7tz5rzqRzM7PPaviZRkKql2FKoh0WT
buoiZ0FHLXLK/NJjz2Af0yW6umqOJdWJ6PqIaknwhPn83deyMI03LxZgkvJQDX8Tz6n147VB8RuO
Gg+hut7ZYawbLF7hB698DInb9VQDOJzS6HIhaytop1CWaSZDH8lILKMPkY17k8GUvEvAR3UcdjAk
dsWhDBP/Usu5NPnHtxcTCFUOLYV2wVSk4GpQ0AM1nVtvE6ud0aX2sc1ZszhpNp6edxHtZLrydxKc
udP7+ptzCYq4BbYzcKVjPFHRZU7ecQtSpXtK29cSt0I2ablruSdKCmDo7ThJBYMFRWsM5R7qi4IY
s4P9M1QoktrhEVHKkrAezeWLiNdDUT7qzFYRxj4F9t862lju9QaSKhwMnIDp7zSZjIDnoaOzPYPS
8Bk5Z07ZxzKtQ6RQ/SqXUQnQQ3E/gRgWJiuof0xJXDrx1tvk2BI2LrrKDSgYcNBDCm1s5mWxFvS+
5lkbNRZoO0kD2UX1Ll416vxF4hn30Z9I3JPEfpLpVFL5V0GbINtlEPu+PWSwmCqNPYtsNCdpAA9w
TyhTEunI3ReaM8rwNV7hBJpYe2kYJkwUShvMGRWUD/Bw+Jd3mDXvvSHmvdO3DulfZABiVeK8qBNM
db7SNS6i+H/E+MhAxxmBBXzMmEOTGeT8IQcOxXo6y+ggiTZZrBzS11YzAY9RzOIzncnBDzLK7xY1
i6tBoIY41awxzGGv0ygahvhtN/yTQcgRN5uTPeNYlWrFPnSo8I041+rJJOlMDXIhCUeyoYVhRspx
b3NEReQ4j4pa68n5K2r7UD+MXIn0QpooPb2QoneEwhSLjJVOzYMDi5UAkfGnEAvuGFK5pGD1Mt/I
DhgW1E07wLOzPK8Xlrcr396RERda57Ekx6xloDL6FlYsQC6FV1Xv6ThUm6PLujozR2L6tkN3PEwH
usQMSEjc32KBKjDFO7uNtw2tUZwNa8xaIZ/mP45PPRnUvB2f1YMrKh3DtD+vkD/eQYpQP9I1vYcA
pxVJV9k/9EWNm9+0/Wf8mWZWGBtonLv/ZLbjKAp7iEN5fCRbb+HgcZLlmd/DxJV5YGUBWjrG+oMa
xWgQduzU5YPbhYdp4Ejt3WXykySDKs8zToFQSdwM9xALIpI1zApTLwaxSo0HvVgpLcuJLGdP4VL8
Zj5KBnJ5e/Dl/rV5IEOLfFEZJRxnWdsDOpmmbijZMumV1/P418kcvDCGBGDlYXboQsJKjUJGLB+Q
g25RwdBPk8+gWXF8J4ThNH4on+tApDICrs1anSvwiXdfn7KAHNDoIZ+i3zZn1qsYHkFwrNiJtQWd
PiP+xmjuyy0Efp8y5+0tUDAQVjSral+iQrPj1NeQzLM9ufU1U/3eTh+Njv1zllM1T/BvaOsbLWZk
3oG/k8w8Z9AqCuyULLaCv9llZYAlRpshbtS/Y6T7KnVjXR8QUE745o7YNYqLCTE9WLlJZzyHSYqz
458ynxHl8tTNa2eut07SmckIH6ki89rPL3WbQ67cAXS2v6LkaYOm2Rlz6TuTRZKOULutZy4tsGf5
ByHwbAPMKPBeyPHV9aOE51yiecHTsdtuxJhwVxjZcfj9Y38NM4F9ac4j3EkoNlMTR9XMjlxHEfBw
85JbARZyK2xFvT9eeeAZKl6T9DqiruB15yP65+Jnv0aBgt4spo+i6w2/w1mXua53Xn6KU/50nPTu
o24mEBvZuGC/fRFrNCgOrfxvzsXaypcIMoK7lXmya3CQQfmEGJH5qm32kbWpYfShoGmhietwJE7r
QeJTPz6aQndONDfdDRjrGohI9oi/k14qaw733oNlkkrowiBKXxMhusq+9xTF+i14mMLNbDBVZdIc
5El/1QOQACPEGwLblb9rL7jv6Mh4LJJv7XVFmss+/jN23Xio46cnva5njqGrGPHM2anfbc8ceRT/
cgt8iHZqQvYFAJN44TbMfEQ1UAlXbwZu8HA0H0wGabNAjyqCqkL3nKAT4zKFdnpmkOmmPwJZ3pze
2a+muEjLXmTkLlgsG+MOXSzpDuIBeGXiuWIjfuXhylQIL0IZDPHDNz7qhX8IErksSTJY3+xN9vhn
JoevLYsBW9sb3b7pwnwu5aQc2Dgw3v8RO3NgxIP8ckciQZg6Uu6DpsilfxXihpDzQ5qrRetLZe9B
Dei38Od9AIJGcuFG+HAOn/2NiCIXJ2p2M+W43ZKBDaxVromK360vJDGh/Ii4d/mvx7UQL08461/n
JOotMshSV0/hLSxvs73YL9aXmCYTzONaRWqGy6YlAPCiXRILmQRX+K5HELGXEl0rRviusPvt7TR2
Ci9ewJmRjYmLURRFu6abu5tc2bFFJP02sKrS6vzYb42SEOZm0t2jx76iIZqvnYMLLOx6YhD+etWe
tDDSRwmtR4GkI0dw0F4hw2RjF/xOV5AIEw2a7M8hMfZN2mcxWc7Kp4g7XRYZfPP5/HM28fvwRlya
gXuzPcPYPRJqQZDWy8XOJPaMNa7JrKHCaDdhOiXlqFHvPjkhjDK6Jc5Ve/RMUouyYeSCVBOTUfz8
tai/TjJRSthInwEQImKzkXiR7G6JJZg9HyxcyW8j4HgSeLaHp2HGBZUQjC6hNMlAC5UOZA5RXEqr
c9B3sVBasPbr9WJzQyuI9g6eCTtd2MrnxBWKEQ6reI39vf9w95INa0ck62rca2V3rJWMu3FluniD
qicSyhNLHEli2D3SxsthAW8Mn1BucKKisbexKBwEtRqVzOLVWNLF/mlhQzHpTp5mq/hePCYvCpj+
AaUmcwx7d2nrrOgXzmPr+tDt+qlMDeGL4PUgcBZ9u7lwV0c4orNOBMBLpAmet9SytMJWNi0d3SP2
CeLJJ3TnXTRsQvMx9Pp8YjoZ4ioWDU3jy62Pr26GIztRh3buB8zVI7ignoSRv+hnfk4rv0dFPcvO
9Ve5vgdrMWqDAu0i3sSl8eAe9EfGMBDL7hvaNozb6TzNr0WKodIXdEklemXS/tcg/EUiv6Gm1yn9
N40EY0JVhcQ9D33bTu3cfqNb0c0g7NkhyJ9omO+N5MdO1y2Op1i1MvLShK0CxEk63BCtBZXjPQZl
lQ8ebnC1N9lPP60bDiYvdyhxrJp6DqLctzanyi+IEJ3DUTivrhGnd1iqlUehAMQDBqkylpRoJDiE
HH0LxzXjJ4YUBSCQXyFyx/PT+BptAlhTmnQqMUz08504av1uKnVsF6hsTn08tWy/Pnq312W7YMd7
RvmqRYGmT4FhiNhP2cjYqaCj0iy58npQMHD48qa2Rw/nW5V1a3c2Fis4HaYW1Jx7ES+XC2RUpBZ0
F7iCKC52/kh42+MpTbb9nQ98K+vcepFJ0D6q67w+ZR8+EFCj9Wzup0gBZCG6uT07Ba0vTVwX/SLo
r3uqUnX2VJGJ/QTCZljkSk00b0gfbOPeufC9Q8A9oGS3TdeEsub1nqfU4x3n+FRa/B3mhFz+a8GP
kQaYSTBcafnbd+RV2njZWKtz59Nq5/pGWN9EgF4OQA+FRN4xgQnnz8O64oLmD5hFWCGZpJDFHYBP
sa3GKZx/4TQwjK0IH7M58RGgxB9DCGz7XLKCsvMw0MvkLk7yBWXbwy4j3e85w6RouF1c8pAb0ZCG
Z1WB2cdjisEMI4syl17uX9wR2oMKJZ0IkvsgXy+ljGN0oErdi1pchNJsEbOYV+5P8grQI1ecHYFD
Wb1uYDkyrc0dibFA0N3Ql28ySWx8tlucdbOnQ+ddSBUHwMh3IDRJifPSBQj/LW7IDE872vGoLd+T
vV45U1KrjcFSCM9aVnJi7eqklTucpJGZdb9VXZEeEjgr2TXLnJ+kGUHPavxizQgX1xTAmdzqKWGe
RL/GkXpVSlJ45Vah8xE9AUF0+52/06pkH1FCkMyJY5qX34y9P3Ldy/l1JTvVIDdycAgo3MRUSb9/
OPrNO8Inhy72B3wTFDcXGS+st7KH7DSRoCeDtJH8Xy7wAQChsTgEF05rwZMv7eJYDQHONn5aUGcb
2WudpBsegtGWOgPKHbZNIasZvJZMz0PPgI8Gl6UWsH/Hi/YyjXcUSX4Jo7VmfgvxUf3BCmOxFbBO
+2Vda8CP4Y0vcq0vXsRRBrviG56t40mGz+8pjtI+d5qGPQAgnN7U/dTG/qiumXc7/WWPuh+bjJtE
PfYOseLYjg6a/fy4QpxwbRgwO8tE28R8AhQzgybdz1p39leE630VevK2jASRcrlHJ71wKOw810A9
g72t9qkShi+E91+uQYcFVE9S4z8RcQ9SNJFwbTnFIhDtm6f0rpv/0W2pcON20LhTHy4+SRSFxa6s
wjFsY9bLAmhwqVt8LT5x4pAllHl2sLXDdizuOzBokz8u6wvNziwzMEVgk6ChZrEPKYrMR9dTVhcR
VslykYSl8qKBdj5f3zQD7B4Lg0nR3LwBYZ33NHMdfZ4K+4OE5uNT5UvDkO+x/rguAtFR+ZmrRchJ
tV29gciqO4q8uYewvhgzCJ6ADvoGgctWxsMgJQOuSTYqEgeXTR5j2jixHnBcLDnritWDxuLBwZw3
dtJTTCcDr3h22ud9NCRvNza56kDBVmkhDvfrJNqyQyrRuJf2yFeInFhi07izzCkSuNLB5jspbL2A
EyQasuPM2+Xl9lozAmilKe4SvoiU2b1kP4QBwDSGuw9dwgREOFzqBZM67XHrc6Q9PpKfq84ehzgV
DZmBoPFeTMdvv6emmN7yXCs1BKuQBVn2XqgGii+KP4rRkE+33TmSNlCb8HCh1qn6ZWZyeqS6vK4L
I30Q4xv4AjbRlGHQe9XDj4+IRRF2s5ooOhjotic6UTmQUR6zebE0y50GMrhExFj9j3ELutC+LoDk
8XvvzrET5ZbVwm8WXwGGMihdDNeh04zC6cYnFGFM4MAAPJEQ0KS9EQvv25HtoYnEOkYvzNyrFzD6
mwrwBLBRopqc7xYoYQHIInqz/gORcDdfuCTbe0abP4tEydkYdX/F0WbD+u24+uU0/1Y4S+olcOK2
PyMocVPiKod/npMRVA4QHfCFibhxLYoOYoUe/zSDUcEcOydJfS+d8aWhHS+IIE/MxPAND9NC5Q9v
blLHvm8clEUDotORreqV/aQ5i6OiOpcKmR3lXS6VntPXfyI4/zCt14MLnK6RPgyyzeb9CVmXzRPz
yJan3FekherniUmjTUSoKB+oh/aw8buzOtwEtLpBcPP9+1oZfRVedMrGIRf0k0TRYOlMxyMZSjam
6lFLPYX5KlgnwLjzcI7LN4ZoAb+4nRRJVCnUnbszbAFcklnKS1TT9nPIpSMwvebR5aP+vhSdDoh5
2peY3n1RrJs53tfTlud2QFVaQf3oSj8K+3b2CTdZobivnx+DfcvQJmRVRv2IDsFLG6fGPHzMqKoA
z4v3mlv9A4jQIcKKbCewJSnSNIh6/4NbGcb68OzVCqX8HU3n2g6x+JQSPEr85i01hoKcXtGbXDh8
CC8OYfBt90PDRztuqOUMDpVj08tXJDhm0ejgsLl42U0gAy62T7D/WhP8WRZZWq2vUte2RIPiIQGh
IuqWWrzYu0gHyod4dGQ+JNG1OaXrqABmhH0E9yM4kcxJs5Pl6gqtz7kLUpjYhxh8RMZXt5Rpbsni
bHMWnnZRaUZR/olHEb8xxAfmoe1pEO+Cip5JlioKsbPeTnIit3eg2A1ei0hLHwPLmaip76FSgvhT
7OeSPfdcuie17z/MiX2ZdaPxCpQqwcPtwpKMvvGT5DbiJQsct26TQaSgljAURCjpeTT4EwGKPjcx
vJfBkT2OLJwZh/zvGdlLnLjlxe+C19rRzNlagPPa3yJm56tYTDYU5clz8qQO02Dxqp1RZ+jMFl1j
RPyUPLIEjbr3kIyhUkX3Q5igQY5EXsALVxKH3E8zp8H3pxvset4qm55xp22MbhjStOI4JKxKCgp9
UWNyZlEjCpjga5tzLQFHzsnTpEttbTXOS/53z79Zp3DL0JWeTbgdCRdoMo7UI5u33VfA22vocaEk
nDMzaTt2ebb86Zsc8Mfys8hgibjjFpI4yP31/w3Zytjw3lyhNrMmzv1L1wt8mGodqOK7qF7MosMd
4WWyoS05QHdR1+kJ2c8fnLNQYdyUmsbWJOH9GdsqkmTwsLSCeTjgITUrp2/f0rnWGPZl1JhdB0FK
OFhebKwJj7umAPfzwq5gyS9/oeCi5RZ9N9ioHXCskV1yqHLiNjI2jy9Ue44hVFxLcEkPUq99u+N3
SshC562Uz07lBZn+WAOq39zBYjf7OT2UuDBRN5oIHK45FyhHIqBPi3SFNS20rePNdk9/EE2F8lKk
vo425wI0QbPz6KsrKQgag+VdBaUiKoHs7XZBstj5Uo8U5vgisKB3Lmq0cSYhJODvU7vJxLaBDwLJ
AItEcAQBcjzxAczQ/ESDeIHH0GfVh0HcgDlb4nrpLminrbhdVGWz6nwsLwV95L4KD20frS+iPWF1
8mo4voiHv4k7KVVndnlgTjS1pjzSHnnsOq4PjEOYYSJPDLYQuhM6sB5ryffG1M/ZcIo6xSsOHugZ
REh00U58Qe54p8p5aGC4hRmapvJVXY70aJ4jTPeVc0vs3afvqxAKZyAU6V/z/TGo2EfOyVmam4vx
6bFx2U/Dt0QoKBTtAOxAbM46XBIMR4ePn2Mq9NC01Kiqg7FEnq51rDuB2CZWphjjNhkEaU0MuLIk
le63TwxQxm401/xjlumLGmwkY5yO/QBJFX3RrvWd9Gta9BjIUwxWHfF18yWxoWvqcFhP/Bkh5WZr
DlZIBj5JxZZUmW238PJmHxjTno48f5/sqIymACrFL/GCG66yBJfm7+X5wCppqE4qWljWI+xtJM8A
lu5perKGGCvChGxIQi50VC5BIeLqiFVeh/dramK+osdcaMZ0FNQEZAb5IQJT4VEr8S84kRa7fuVY
UHSJ+hlCQvNQQNFz6060j6+//HAG+MDUTzclvRLPV4/N5A/nyyz0S/RhKae+UaWkimYHoj4AL/q0
BCm9Seib3dOG24CtmmC2sAqHU3tMq6KAbGnAH9DJErxHOWWmOENkOSU89mG8TB2MpsJvja3BhH4W
8oYhLHp7M8KfSO+fjiL8fAENSZXSdn93NuXPejHnhDppjgeAwA6gafCjyCX/htNeYHwGTdbg2DUt
oWPWu1slMTKHta3y5yAw/z0FThqj9jMTyBjAfjTd8ym6p4FFqs2ZdlKG9SaWBlImbGPzsnvkDOsj
bjZ32AaT9AIlBPzPFquSpqrsNaWpN0HnkImB/s/kQEBJXUUXTLoGSUvcRNYYMJ8tnr5l9z5NHR6J
SMIxBuSkUZbknCJsk2onHVfVv7nmNIwFsOmpbhTUxE3IXTSaVWMCLnrAvUhBaxW5zKIfkYXxS2wd
UQyGxjSVyclEFF5ukWs65eiiA6uZssCVkL7dOPTEjgjv5HeBqcdWd1vXTZWB3azjNXGpRr+itnpc
J/qU4N6aJ5I2BbNJPD1hXy2ejmaBQOD4KhtiVLhETyMz7jcGfaJMgmWH5ol8cZqVz26tpMu9R9hl
H1IVcQ9Czdh4wHGQTOOMmVOiLXwqUN6mpQ6gLUH6Q/MgCNGchhI/KVtCHJPJsE++1VZWz1Yj1K1D
kIzvPU078KfXQiiHoPXoBrt7Emvl6wHjqr/iUX04IAYiRkgXmsAZc3lbzib3YXxk+peH7lXRPgsI
7upd4nju+rYIeK8Swwftxl7FF0ujq1ZMcTeDt0Ey6puJFAoCWsH66GZkuscEKYa7hbrieq1P4QOZ
dmLYrL/TeSpXA3fej2J/geOzoDhjIvhqrTDSLhh6qJPachN6Oaw835m9pjMC3RUZaq08o0jMSAul
0nrM2Qp0kPBwXcZ/bzFvQDPkqiIcK7H+ZrnoECU3AHFIY2vERUgRE/guFUJoT2SGvx1S9jsskiwu
vSx6baZPMRkX96nWrq+X1yFS+Yp0rZ/+X9ylmU37amt+zGYaaD6kdafn7Vz5MhV6mRnmDPI2YHMH
ezUmG/V92USYcSHHCZ7Yt6uMg5sfdFTkrGXArlf2vquR3P4KNZ6F+LPveWIvsPK9aqgHPK8gAFYE
JQ+z46tYBFyuAxSH3k5zKwNfVc97sPjKYW3Yr4FmzUxrkHFcC0jk1W+jRZTebpKqKCn/JrprU/IQ
94zkRv61zpnkWu9vURorZM0ouPNqg3DE46smBV0auFUIaxrseh146vCluaKDWw5PAvuIfWG909wn
yZzfDhxWfqHMKzmAPNQrAf33Rmi/s83PKsDvwYaUIu+UMjEhdZzzxW8U+kn+a1A9z4nxM5WJ5rd/
8KK7avzRAuYl9YcHUAVrcuUAO2vKSXoLxAe3DgVeqp5a1MA7Y989P6TRMMFZI1+ZE2D7MeeTT7XA
Tc5kcaeRuFETzut5NX+yTU7LG625DbR6l3ldB394fFzRYndgTdp/8omO94liUU/wExWgb8jUN/UO
SQNcqWyVhBifYhhGf1ktgLNI+xegpxQMGJO+tyGJ+mZVWk29tult5VvwgdVedJFdVJv2n9g8LgMf
SNIxzAmviYvMzzU5jpao+BrSKILkjkc+AskVQ2REBQJnyM5TcCPpU8sI9u6lqaq+4kqp+Li5/gme
3PhmB+xidkn+F0gbMvkLrZvu7KGCUyB8aounnrvA0qVd3kjHIbisJ5q1PU7zy8/aJkNu8ByJQnYt
mBazizseZpjRpD2eT0iS40Scn63dIGd7nq5QZoKyy18OiOmLhh9XsQKl5J6oZreVaqLJ9MAyhNlT
vBDdlL342mAb92YLQvDbVxXkS8YMAU7SPhmkb/mRxpqJMaAAJtIx5ADFxLbhO2Dt/iSLU29XR+I5
jucCCr60Xzgt/9KnLq5ZWC074GVOJRSPPeXyl66nwHaYnSy2vOXeMI2lmdmomKajYwf+6anZoFFS
yj1sRSlqU3AQ5BYUhVZWolXZ0EN9C9VMDZe5iUdetL2QF+sQ3l9vKiNHrzhptK8HflKfeMwrtoff
vUxzc5b+qWcRZ4EJtGWj/uu9IjNPI9r0X9bvYFuYGDOOyqcOEiTjVd7Qqdc/K+iFrjkJCpIbZneT
upPsoLfrQV0/nezzP4j2xe/BTHhf4lU+FFo9IxeIS95A6szmDIMcWNrKrmc6Oanmu0zmQc/0K0f0
/CoP9dsJoOeL7m8+W3H3zeLE4t2VG6yc9xaEyMEL82BZ2mvjpSQcWZR/jEFRLm84D8uWdIBuYq7V
ArWY5PUBe0vY9fSZ8GC3oUCSzXnhQ9iNu2ivEVHWivmU7znu4xgoP2wQVPSTNAYKrA+TYuNF324q
Z0XwAXwk3vY5ml8Ctq2UzlqsR2ptAlz0A80zBE86peAJug/edKXHBv1YvBtiL6DYyFbgijWy9IXe
HqVjELRK3JmElLUe9ltD1lIRWCLiyB6/Ghr8sykPK2bahr5e9N5cDkuU4P/VxCXMOA0vTOfq+svf
jUiOIm+ZQnStnt6QT6izA/M19WIJaBuLaKI/vHzlko4oYNySUJFqxGqLPWJNzS9Xj4RNzaQvq9hP
5lmiAJr+5cFtuiRoZCfMvUU1tfSfRW6MqZxdVybt1jRfq4aZB1ZBdh8mkhbbN+okl9YF2d09roh5
U5ujfgpfChiBBdNq27FpK1OLDqsNh1XXAn0LV/60YbNH7pKVCHEkNdhDbn/XLYczrMSauJa0Opdg
LLGr0IbC6KZ2hNk1eH3Y4VQo7/FRsMukDqbkxTf+Zc1Fd+LgMyKaecYHt0l4ffvQBtFDPtT6jlN6
PSWxABBHqNJN/AU8c/PICITTHiBv0/jD7JPZhk0YfYq6UeZoksgHvKAfH8Md8S4UhS/Lb3Wy6vNw
gIzwVklgO1EKICWq/SxuO/iVDJT2mXeBiCiRuuNeRf6/IdZjjtJYK7aMv7kbefu4ne9et87FkIwQ
j9hdyYpv3Gu4wpDdXX7ASFsroVOBl0DEP3L0gkxCr8EYXlw1FgxNJQHp516fxBUSyLlQcuPO4bnJ
OSHYdYAdELYRVoS8tJePvM9Fid0AQbQeGrx0S3UVow3zNBGeAfUH9J9chILikeK/AvxaMPeSoLEb
8+Fpq2Kk019sg/khNwnEoN5zl53fHuaPAhqiVc3kMKcs15VrPZTX/MGzNjoGQAslfEFsbRJmFrwd
k8+Wmimua5JBkzp3AXpw1/+4QSo1+LIRkv5QOVEMhPcEM44l4gYiFJP+QpdtQyNy+uSs/zY4HfpB
uz2qaBXA7EQce7AGtFuwtCYgZ9EsQM2uHIDz9ii9mWaaH7GAXzajTeT2XC/sGs8DsNs/6A8JpU3x
FL2rrpNE2qzOmFxzBggRcHBECjcnXdNiqN63OedQ9aJCilh/aSG9YvnHNoAeyGuJT2v8lfSWSnYt
PUkZe9cmLhVlKeKxWgnOn2sC20P2svzHc5D3cYV1XksvwO0rbpPw7RUIy9HTa/X5FsVRCZNYQW6K
WOk6jK5/xA4keOU84u8BM8qrliLgE9nN254/AGtvHwXmsjJm8WYqCLgaQBcqrH5piRfrLsSPa19F
9OP+8D7TRzGZ/ndzvFfVA/EeAQQUrLHWN7zaeveVKJHP4i22lkLruETp/7EZ138o6q2jUPC1i3M0
Xjo3e/FrSs9xuiTuUcZ/BR18L8RNS1spbj+uHG/z9ino2PWK1oSbYH+pdlmm49TYgQiDQiieGlBY
3hhapWPTwV9/ECbigMghJFq4yUwFnyZcsaWAzRVxbRjfRzMAi/qwX6d07zMfKwlC59yWMmIxnAL7
Iu7KAW6fYuwoL4ixSDLVmJ/bZ5CMHFljEg8x7QNcvMDX8ktw40mtWmjdL4jkTVb1I6omrvDci3hQ
CPMW2+mFlnYTHNFQ9its1Hq9YvsUuK6VEtanEaoDzF+iJMGHPSVBpmOnAo8MHRwn0owhzMkFUEI7
JOSg28ht0QvJ9+QHNmFSRehQG5ZYHunULdY5RmYUf7HNRQYLph+F5Q8uYLo9Ir4yzsAw54bnXuFr
Mf8Eg80q/WDloeugtD8i3FWoJezMOV1tuM7tYjgrkQfMatZfhx4j/LTjCEWjkPXC8MSEUqJ9o178
cmQ6hPT0JtF9AISfXwd8qKLfHmvctzug7RKR75ABME03Ci2GWOJcv8YLoJoDAIv053b3vk1Pv10o
PN8C8AU9bwsgjfIrLku4Ej41QihskeSqFVVdMm9/m9GB9wZyWAFwfyozGHSMiwuRuxo2foEYJoYt
bHG9EmDSxbIXSKoIkYW6k6qB5j6JX5b0mK2ogwf0N/Kit9+l1y8Uxy0soRj4HzdHLK+VsErKSdjv
kvIH0cCsKwbTXSqqh308DIxGMIpcHjyC+Sa0VNwuyXb76hnILlc3IyZAmicJduldOw6rTgkNkggJ
muGwC9wrbB2lMRYLrFrCxM3ykw7jCkzB69dy+p9arPnuYyWX3wsLKqjbwSZ6JgZ0LY5bYVzLAEOB
Rlc1I+D/F3dLQea87HqYtsTiLnxdVmPlQiX24vFb/DoumrxeNm1VWZGu8PsP8UFb2MrkRKEpRaeL
hxWMg6c6NS7LztgngiHmye+/cNfKvY5mlGLK69TSogku4lxOvVaTLT4604sI0WCa0mp3t9EmspY2
gCLPdWTcAEI+UhlLXFxG0B042N33E8i062WHMPSNKcwQkETJOxM0jaK7NA9bnBDhLQrOrdJvW/x1
IIMZsJ/v1gLo89/6y4CmKfVGnyYTg/EO9d5SjmXzW+Sk8LW0FvGAbeFyiv5GSZjx6V3OW4ptXX24
H3KuwG8tROJT0RJ9K+wO3crrGPKXXxts7+8X+4UFn65Ryqvkqf+/7KHOIHaKiRV2+coZQATUUbyM
8SaGqydDelRpdwoDn8K/s3R3TBe7E/QCB2+cnwqA2+BdA4R6p6T+emqXE2GwD1NLnLNySoMjb4nZ
aF9RkVUXVUQ4SFcyCq8om2PsGBHYrLpDCGYEX3AEgfcbh5rW0Jx1TxVNUvxtqzXEftJpWr/D/Y12
lPZqK/e3235gKzpSVNZggi2RiHO6q0o4e8HUEkgOFOvj3bItLmf3oiuS3MnrguGgM6DbkVflJa+Q
EsUV+sjL8EwjcYsAB1Go2HoTvG8na1GwPkvNFe31MsP12X8RO/AIKYCE9uLxv6cpFwwDHnIlzfTy
yPy+qeP92GSMsLKregH1Q/OMR+SIIU6d6tiVPJhdBYJ8ueRIeP4BtWa6yb0r5LZThCQLB0/HiLPc
fCaZXLy3jzQbVTcLngNtMZEk+H2DuXFcCaKQj8+y1g4X6ShtKYrG1b32Bku92GjR0/wC5ql7lQgT
GWxFYQ77zZQNYXBZV8sVkZOf6O/uSWMQL9fn8gNs3e+C5Q8jILy8qOug7F3AJyRGjlLA5BaeX5i8
dQ5FvtQKi3uf6C/SU5QBRNH/rLmmbdfFpoLsYE55iHzx1B5SKVNPZrFhASuyxpCYaJ41r6fmDteM
cxQ8MSW1xVd5LTsRq0tJv9sHCBn8a3S0iCLGaLSTIOwKIxp+g9V6CBlNfKOcOoLbz9XABmXpTGOh
vES4s9pdIq6rK92trX2QKpVfYsgtwnxgWkCnB5+D4u31pHTaImCuCSqurhZO9wWDLWk90jwCA4zh
IrTGUcB7zSNIHygYFMzEQ47yKUo8Dz0u0K4AcJbPBqXRx3LR7I8/A4hh8uAk1QnriO7W2dtrfZo8
fqEeWMzdFAYlylMzOh6H9ZW1VxoAyWxexPPy6P2SH3liMG2Xc9DEhILE4rBwtz/WzclsszpytS3X
Bv0zCl0AFjLRc9NnigEBwmWKWmsTVsyMVGAybzEe0/+j7208l0gNHWvGyhlicIL2jf+/hOZYYLsG
UOpYwMcjNGcdwX81qWUStJJc5Tzs9ofgrqBnVFdKPWl1PLcZdiFj8B4Y4npzRbPLrKiAkrixLNsL
Xf/9EfVMK2KNt7XhxI7jIIUFaQDwq8kboQ9nCbUeppgg2i7dtAHIWHau9mbfHmLXKLOfn2pwcX3q
/AM4wmQMfehh3UkmEBUbpnGGwmkXEFY5IHH/VdDv9sHW1efEiOSfhaeIii3ZKtSLB+dfOktugxeZ
PiXGEFJ3izU03UXo9aLgBF8cPZH6lMWSzJ9LW2Q1BQhegKLorK8+FOlVOEVFZHHLAudD73qIgOlM
JDt9oPtjtTgYGg8t+KtESmJPMELeh+2tUrjwauSOPnukdi3Oe4JLerqafV99yzydRzxCrf0x8n+d
5VxUrBhHDG2Fgbp0Mfo3O41I5DO9rO+OcZ7J6YnSqrlcXkA03Wv4TQZmQlejtYsTHljtpwfDOFsc
WTevw/hn1HrniG/RAaSrFNsclQLacW3QiPqlUC7taVtSaTOhTIdhqkdCrX5ggBGYK/ahBuzwD6L2
Nulbvdq1Dn9iXO8Y7rgeWKhNEUcGGrUtDrIxvWxUtcNJ8hNc9I0y76ooMPLzxXy+s4DPyM1T3LcL
yLSFgCwAQDxeGlKCBPQpneTQSotOHLiEqurXP1139Fp6ZUXgRfTl0zghdV/eW9VRLIRXeEEELy2Z
vyC+4fvbRCAK1v0DM0TfZwP0eyKNrrC3LA/ES+GnMbTnJ0xaeW2Z+sZypnUIGsNM7z2iUDBLQiwQ
+hmMxB2NrlVYAIgma6yBq3r2f4bzaW/YxDb2/dvJYQ6rix0qEyXGCGLsQQdF4KGZ5Nb90W1D+dG/
y7eG8X4le7L8ZgBAq7xelY8mb/b3dzAz0LjCNqjkj7k51mU5S9Hg3cRk9PzOnafjrl5r54BPJguz
iJO7j+Me/E3nct0avon7xfAiWft1OuhdQ66zd7zmbqqFciSsYlDZorwxK2yk7zPJI8w/5AqdnpJP
I/ZBi242AZ/pdj+0pk4Ht7mFCPMJA2l6FUYVep/8H0rVQcCXQQY6ThDsdMzIenQDW/p7JA6ZHcwT
MdlF1GtS6IGFq9QViS86aqqwTmJE5nooAmsrtvzARPcIrvpkyrpwyINcJDzqQjfUXNOZCbN4VvFS
8stCxat/o+UE67goF/mjINd4eX3LDFk+A8xw8QtZOp6m7qrf4bGv3/LSZ5bVQVrxBGFDJevRwDoH
rdK46PTLsGm7qUvHrfqIZ503PPjQj8rIL5h0iyzLGHiOBPb/IGMzM6hgOZljEAUNpMVHHVkMST/v
4aERFpyUEoEqwptj0yCDLY3Wfk8v/aczxo3yKMehkkYGvf/OgmN86Lw7vOwCDjLNXHqdQhUH2Wwb
4OlxltS/OxcpnGcybJc27lTCXxdZOhI0gT/CpNSxitk9xlhwiJFAFOWCQbpFQKAuo1MEmv4RPAHK
+HlCe+DDPQHoVddstXHh8xDS4exG8B8mTR2Hv6UlDoHocaIFSFvAPlYGZZejcvDMXHbzoGDhWqNr
MuUTPjq0GCsLYNCNz+66E/r+JCk9ltJgrzbrFVs7WXcE5n8+w5OkslZC9xX8xH5iWrXxbqA+B8Wz
7xZKuHkrfwPKK8Sw3+QX3dzDi0boVOzmiOMVduhqxZTNSj9UDITHKgzlT4+BRMMBESFOHrW3dFU2
ij7jceK4ouGKoqeYjkJIn2AoSd4KVYfzzZBq+yTg37EO8At0UAGxnLn6luBTslOCXoitvZHB1HX1
GaijCKCzlEsDsc09VuuBZH46NIMb5FNI6DOjKEX+owbJ9oke6U6OQqsONcTsdIje4iC3lDzak2Ny
NxrL29q3QbvRs5QE+raxIer1Uf7uDOs7H6qtKDHhjwM4GgbXT1q976qweUO+DjO+eA8X47O+SX/U
k5+nGSxbRaTFInM2h9TmTjgUOFjT7DvjrCb1Q8iW87h3PD7Feq7eznfkcqaKSXSPmctzZ2kd+frQ
EEFVrEpmwut95tNRza+t0pKzy6vTM046EF7/uJlFTszSZ5w9ij4t9+nPxg79G3D+/IR+aM46CaG2
CPHntNe4RVsGdHovxfz2N89g9s0zj1xYDXPgOcNzNL04zLRAuB+qIYi+h2VaGe6m46/th50npYyW
LDhUYLtk2JsBcra0vILNO5Th8C/HAjdjeJoiBp11a6vH1vBtqrmUZ2iz5z4H25EAkn7JjE1uBm26
lGglY0D40Q6FHtDeafSwA1olj5qktGTGHle4iuTjUfl6O899En6XjZmzYA7UM226bXywhmzc+4q1
8BbCXJLFLwDSErsMKNptDadcJBGrmCrTCKbTBhuLx2TqbvrwTYPRT6g2bTF4HMbGO5hVI7dG25yf
65JGrzYYxxlP0JQ93CIZkokt+horMCPBvMvb9Niu8T/uNNh4vW+5Fe//gV9RYgjZ/su8PwqcRJ1n
fKPfyq9wf4DANhJS9u8TqlMWiZWcZ+1FvBz9cQwUsO7AdL/HbUPx1OnpzaYl0xVMzstBR4HVHKuP
MiHzRemaFPXfGigjNcloeR43XjRW71PSXs0oZZVpyo38tCerXPl4dwcMfFkkvcW8Sq1AKL2J5FBe
FG13WXHGpvGtqq1Rt6/W0Mrz0uOJStg1WPxlbh8CbwixySAsjhZFvOMhkBBxJWwqMmDgoClOYYSS
Uqgw9cx70E7zxgKeJNlqNDS9CCEXw2Se4o3Bz5iffOV2BZf2NPUByL/u28Zu4Me9g32M5LO05gKh
Ln51T9GjFAdPvPqCtbMO8h6i3HEw3xVxUdEigz2zGEmNPHr7w87UH1OtfMRqvosF+Q7E3QR9KzNx
pt8ufffbOGajpV0yXIjnN95eE4MtA3kfEXwZiGaeAWbwapt8UML6nZ30v78FPdxIvrcj34w40RYo
yTUNnn6n6TAf3g/gtCzxpkaza4ts/AkemMRibgzqYsD3wjrdCQ/wKQxm1I5kEBU9sAHBQia9Xnre
pum0+4vDHyJm/xM6zb/vwMatO/QpOZakO+wlg7G+68UKj5hIHdtipbmvP1tYflN5Jo05DMQH6aJ3
HvHry7yxfaUNueTy5MzQ1UYJL2jRpwGj7tfg7rR8Tm8vB5ZUbsRSmLZlLxmW7gqbB96SI1D4CNvg
eh0enQhjTksahPX0aBhlGemhEl5mKZoOl5b85S4Cv/tby8femvf2+P5UanZ78Qsx2rKUprZpOHM2
XjMrIb6aW5qVsP06YiR2xyNbi3NSUX6zmXRt1fnm9udJi37BigGx3OP0s7roSGWWMKjcNjn68KlR
vZeJhz31uDoI8R8d4L/6tbR00a0jnaPOBEAeMb5m0sDY818FVamLpWT9cWhtWAYmI+tUMy3kVOVg
LHK37OY1fcMWjMnxTWHUGseHkPQX00JY1/RTN++6YDaKcpn5W8DhzO6o8TMhDKX4fEhFg9vAKkf5
E6f/gBZZ9pzEtrOgtR1fbxTCO2BuRyqFLmK6sdho+XmGZPjYprqR9T112X/vzkaFED0RTXmTRCLz
SEoulAk060l5lZoOHTGdkr0Hb6V+Ti+nf/Z8Gv7iHKRL1snHALScbJMpE6N5E4WMg+U8aFFEyR+e
TFLu9zfJzQFm7tUKDk19ci8Gv6f1jInKimORVJOWyVo8OSeZX39hIh+BHNu0kI+o1ektQ4suu/pP
CRxJtVTrpUBKXjph4xkPK9DVzzV9jlavpF8HJB4f0D0Dl7EbbvdMVLI5ir+fGv03SqVvJR+dh32d
EJ4HV38B50yPPViUe3YYYWnQmA/TJrUUNpHZ3iSeZXHeJSRxHIi4ciwdZDy8HXt8+QBasO5eIV5+
VTZkQqNUZDiOpTjYHAri8F5G3jscHnjnFSpNSJjw0jXSHL7Mo/t5GM0FNMzHxVF4rTNmluBtsQx3
ybqyYQjk8vOJ2EYp2Pci/700OtuHkIMrA6b0DycElo2VFXGRFmiPh4184ZXwhr+/6Lazl/wmOY1e
Pom2pBhWp0dFwsF6KXcIaefzDRy1xZ8eLULjPrWSAp7FrgcY2XabVnu1qEBzUqm3LejoZmkblQ8H
8DCwipl0R9Kon2CjS35x8+U/uvgB5NSVcHfcgII0CF73GQPFf00JpIm6EOE4n80W6Cn5m4CbakEs
WTFQS3KFkzd96PLyvxiI/6aHzNIhbe0HGeh1HtnlMSt8asyPNbZkg8kYThGylyYQq4x+0T1cuPCT
wiIWt0TUqgoUXbzLY7IqZG1NznoreKSrjWIGaGoNjuGCwtTLd8SvPd9n2VK18ml+GAt/e0+zdadR
a8a1//OSJrPIyoeg4SbBb5yDcee1jZY5nG3zYs2g5jRBqp0CPCNa8vU4+sgpXLLaUgW0soC8JLz1
f9MKj8PopFmUo46OGCD/dhyp+iOTDKv/8HaaYfaH/9ITImbYA2pqOQpqXDR2ux51Ikowg4MYhdCN
VdGQtisM0n+7z5VLavlUEHg/JDq7u2YPs/qmmXrE0Krg63S8d8PvHbRmP1IwYnK06UTf83dgciFN
p15C3bqcaHd3q+GxKYSqT9h2wE5+e10BIitzu6DXMDhpKbysQlqvebF2RK9CZATm7aix1zogsvKs
P9nXu1Cq2arPsOgOJz4hZaBCXjovY/iTagqS8agD0YfEA+qcvNdPvB3Rj0xFJP+miM5NcnbZegBD
KzgPRXIKW3CKieSEyXaECBwVoTdtdpj3LstOntWNXyaqK3jr7catpG1X5ny/Q5dGDTvbZu6gNJ8i
1alRh/k3DsEyBGGZlQj33OTCCeF39gG/ZxMyw8pz3Boy3L+6lPPKoQbaRjanA5poZ4f1ETk2iyMN
neyIeP1pFySC2Pc+AgBRLLHaBQyM09WXch/x5nBlqRfdM68RITree27i1TxI/aL1dYWLdPgeTUWq
BFQXVr4ayKWMpUBgAS4IDU8ufhuU2DZfIKmYoMgh/rX9WvVO/KlkPHyyNqlvhKk0huTmUZhly1qK
3SHQKTA9sFZAooRs931F+Of6eBSHF04Sb0D15pjcrJp1APf3tyl4EBvsXHWgqrAK9KSnWIIM8zmX
VBtf8swGunux6Gr+9nkqoX2qIXtiIkGGYbYJrcw2Qh//Cp32Oo1qZLTn32xVGzYmCZ/4jh9xR2rX
XQFHaSzAlD6SquPOIhneXeuzftdxjjq3JeM+Wg7H4KkLxrS3p1LfTSsEPnDabpNBeAxX5ETL5Yr9
KPJBqG/nyIOIoqmSRgaINFiFluDKHQulGfP/3P8vZqCG4JDsI4xUAvtz4CNq2R1wmpbEr5xmKEK6
I6RRXWP+xfz1v29QfvHGhb6FaLW2z5f0GGbBPj3hDxiECx2s85hh0GYBly73YH6sYyUXJeK56BFT
jz9NyjCiqxNA9MufY7eDoBVBaatjcg9oVEUHIaGnL32aDSZGB7zDobm2lIY1qyDsYCA1GjrVU7aN
ZvhHnlBguAbQ2m4Yw08Z8lZwVVOoeHl1u/s3eodUdIHkJZxLu/whcOnUmXF4yboLW8ChWsonUhci
YmJ03ZL6eqODGwzHxSAj/WAmsdSag5b6Nvt07qrXLYSiRhFrBfWGsdFbXWun6IsO5YOrz/JMBSbF
/gv+4yW7Rws9/NLkn+24Y1obKwnaO85re3wBlamblrKDx/KYx7oSz7fko7KVbzvXKRWfmpXPifEa
JYJtnAJpq7PScku97NGwgt6ImdxNi8Ec9g7Xg0iqfewk7ldxB4p6QmcFbmUjTqWymv2lkrWbARyB
Hq02RhpcpSyi2PmhXbqDtiZmosVS8aeqGZ3a4sS/wjpPy8g18UzWEwZYS3vxqSYU4ksIV42U3Vro
x0QFzBthJqTLJUX4ytNWzmSSf1a+qGW7DWxM7cdvha+umqOpXrufvtS3xBcDqgwWQ37cnOWeFKwb
Oe/SG6q9XAKPRQ2TO/NrWBUo/tzFkCzMQ+YKQweDR4eTS2y/P084OwOZ12G3eg4yKUYH9YV2fWGC
Q3vtyuQX1qGx9ghbOy7MGCfCAuIfBfDDSPBp1m6Fu26Q99poi/PsBjWiIA09STstHNw/5gI4Gw0E
i4NwbyqNn6zE3W1tJiJRHyUsJNPpWScmvVEUrp3rNvz1UTHNEeNy0VPufV3fpw/BTWvKiP7uq7Mm
O0UotFF6m28eGh0jvWtn8rb/HGdSFTXc+eGi6VRXXKc4DPnqBRJHkFJAXEP1c7hurTupVftWJoWd
R/Zy36dx6sVL65qRBvITJfz0BjoZC7J7kXObWwdXrs+5yuE/ohmst+BgzprgZRoYjiOpwM8XruJX
76CHY+qJ4PR6x+VjDnw++IKrsfihELLklT93kCkpcBQzs0qNSBJeINa228Axnn67KdmVl4h2/5NT
sFNTYURqprvpEiG3Si2e6jzvGh9q4pB7Z+f9e0a7g+4VcBq6ggRYObPCgHNM4GMz2kECqS8fx5H4
NDFu3eDyyLyolOU01UhBaNb8egqtiFNXFJtSPk7FckDpbHAJ5Oehsv79ays3RpPihfgz7Al9dp45
3VgCZPFa7IqIWSbC70wmjedusjFfVJ7WDzJV0FENOfmtJPFmg/OHCrmDNNpe8jffU9I8dSsrGl01
febBhJx8CO8aDcHxmL85YbE9/Td5bQoUH1NVB8TVP/84Cgft9hyEHl5ASn7Upad1lbEzaI2/fYIf
om1ToOWFH3DIciaUCA1tuMY0VmgNBa6qPDD3T30x/NuUgvDOgHt41FqhTNHUFRM4a3L3sa+uaQ/t
xNq0E8uJUty1URDW/Vc0/8OenGhaonTUtDNDUKcegWACiGXGRQNhspQ6+kTNewnDh2Irrb8Zsawh
UtSfY9uYoekwYncEY62BA5UlHMiXvc+6wjP9TI1YYE9NwPTyQAHlZB4bGfvARxyhbxrMWQ137YP7
mC0q8vsozPsO1n0ra1SYySxNuLrR0ly957pDBYSTIiVl9lqfNLV6MaEDYR28Qf9xPkMqCR0DgDDM
sZgwTH4FYV5MxTaskqdOgmh5AvcqOM8nXM4PMrUCiK3LuzcgGf0g0hDS37HE3LtjRRcc+kJ7pnin
CXl4cjBBIm/sAy95H2VKKCHdansijpzodFads6Tn8cmv5KxbIrmfaMQFHfZfJfQFRdIJN9KqZlPP
n+laZhjTW1CaKHQMXiMAbZRbjyse7LiiktF+2ptHGDBPhbJ4tKBqkFMmH/5d1ZsKKvIZkiOBmCPV
UdGie3Rl2wfbBYOdAAmhJZBccFDk55VJMXQtBoe8pivKbVKXaMTi4lHFyOEFAUuOYLb4NR/HcZ2s
Z8AKTOvDUsp+3Iyf4VDGRbQoo/xSANtJRYbWZrinlo9O7ktxOqztHUksynG4/l22m9P+hrbYdHUs
s9duZlx9oi2GMJKrwrMAKV5CRrkyAT+Uj5mrIK+WhH89KmkOAj9GPRoxnr/Rz0b4I0St+OTDrCx5
MGaRa1S2rC6J9MS/02stCKa0tZqMj3DGs3nRnIDK4kR/RCIbt7M3QUeSCt03vX6Goi3GNrwK5q0I
XG9IQcjAnY6l9ng36vONL5qUVrs3S9NSxdyv59aZ75FN/kJsXuhVkCMguTEjbCkdwOP6anMcTGUW
kXmm8GoszSyj4q7TCK+TdDJEABgzVvm6bzEkONTkI2mHxSbmb2wZwIknLXEW0w4gU9zZNaKT9Aiu
gXkWmtszQRWPj4BsnGXpichklvzJzyBUe1QJ2J+O2KARvzwgOXbreeS8gdA6RXvTeISebKM3faZ6
2JfhPXwyAaVeObMhaTTa13DRQNyLCTyvlMnwPOM1GMsf6sJ/tLex649ZO/4jhj6N6QnwpNYYm1Az
pkL1qIJlu88bxSWsgjYp7kot4oogRoYSd5oqqPS0hgwYHdPXO1hLJxApiZ7RQKFI2gU0quJ7oO/L
wdHdeqc2g50+PF3nbMwxdkzNK/aolcnpIs7MFfgx5VJ6ZT/li8wtk0dms1iM1JYyLD2KQwgAVmyN
6omOQhMDJbC+gMwjQLtkfWmyT+ATjjc+wgdj3t34PleeG1lvWs13YHrO9mVcIuTs8dMx+LSjIKXk
Lz2f21Mp9c2xMmQPsQujrUvanbSwOR9ySWE02s2bJQ0Lr0KJ4fmWMqpW7loKmq9IsXLIutDLmvgw
4dOcT2oPcVASp4iH4DgaLaO50W2KN+0CPJMSC7OLrTmtUNahJTrN9QaW9M4F7owHOdYifQk/X9Ib
3xXr+TQQe514zoBSYAcEDfiUJVmS2pPzzJ1kXYMh8Nq1CmzSjUW3UGxVWOhgQvAE6ciPE9qnmdFN
3Zi7VYdHmX3rZrLugYnsIncCytyHJpLCPkAXVXCn0TXjG4GQOU+MWmwbEeAqziDN6e0pMlFIVi2n
RSzkEQWU+56NENBB2QHZu0zFOncrhz8Hi02BxJUSmycslQUAvPAPCilDLRuF+/R9kwU1GImsH1M4
FZ8rQZPqK61GiFqCJ2XSKgX1h9GOY+o4ictUPVcpdCQcs2KX162lulXArUfrpJ7OFpZ9d6VACgtb
UdpBiP6mrDiz6XmmKzVx4dbirizWkdHibzWuDdeXnJxdRFiYT9qB8xuzoyPLPNG8CVvQO7/JZJle
Vr9jnp/KtOgSyqdBJ4zPEMu6QWfQYuCTolmvlDx35XtuVJ2ZR1Kp46B3eWek13BdGW9tlZk8wUOW
P9SmIJKQNSdoudp7jJY7Q/t+B4FdYL/s44U3vMA64T0u/HD29coMZbDSNCoBa+pr+CHqCemqAV34
jknEPBHoeKwktAjQ7J5B7+bHGJrqklkT/ljr2dxQlbIWZ9J7WSzL500I8nHFE/soR8g+X/ozZy0V
8vJF97bi4EaHBieloDRNL0fWku5ghT2zRn73QTj3gauHjVgp5x4tc79TMQzKtC5W5b54Wcu+eqec
FGdXVz2SlkvLVxYdcRb2rLXk1ztsJELlqp8jq9A0Aw0qrDH3PBbgNIhG+6K6bNxFUVIdLvJm8Z2e
ARxKFo2HkMBx10fttxO8eo2l/7UA7/Qho3MHbG4muZetiH1pIChsWt+IV/APOSTLwc8qTRKMXXMo
GOoG/xWMo+AaTm6p7jUYdpAcJRW2tsPKaTZvQeM+LMLH5GBVICPzm/znWN9ObuqtSA/vUCGY1A89
7uJXgONhTNzQOYScA4PcG3/mxI/xMmjvl1vmg+wJeMV4LkfzMhdt4xwZdyKtVTrcSNSMyC4xNL9D
60NQdTb/KZYAz1X+L0Bt2sbP8Lv/UmdOMnet8uZTTXjDv3mpKtWq6wDpGbIcSzkB/R5js/nZyvRW
4OCSNZHz9XhJE8E88TQxAOBmyP83mFB5sd9N1ZasOw/trXlgvQi4lyM/Q6lA7zlk+gpi1hFf7u8s
RThrtrm1BvBRyLOxEPuF0ETBzL5Ra0emTXs+xeCya4jJjD6FfTaDdvo3Ug3gZjPRsW/LmEZKciCm
z8mluiLiQvwpu5dphv5VpU+7OehtmFsZrBmwLqbyWVtrgKeZ9OJ58vCLqtT8Qcizano4Ok2pi77n
ySuE/xztRw2fEhaOTSvGlSXS890xqURhG7OBG+blCxmyPChcZFH/sa6IboEDFCnCD0ZTaZXlVQmP
aUOQhb+/anIbxse8M4t0V79oez4V9EcI8opCSB6OmXc91//WFsAQkqjw4c0mwK0qzrKlR/EpvqYK
pnb3DsFj0d3fB/5Cc0clYRv1tFKHqElIo3RKchhCy92or9wSUMk6H1g44Fgyy5ueNNK90XdPloXC
qs0hRwrz1sKOkJeM8buV+OQr9mX0cTCAL1ZJalOh3MMmPG2l6w2NisIMZzM3RS2LfYzpEr6Dc/lq
HshgqNSfpzCSWZaktEWJ526PL6beN+bppXKEjiKkcyUjejoEWWAyT3JIBi36GKwiBYCK30BNZjL6
mVz6AFRi1MXdAT2YL8komyfDW4JCB1x9hVbg1rHD7YV53/H8kDyplC+Yfn/clxs/O/qIvyAGLnFu
WXUrkpjEpsfUDg9AKDOGRi49zTHPOfQK4Q4Le8Puu/a29QdCjd8nzL85lHJ6OXPBzbBJRhAU9Rka
s2tYSGpvI2AV4eBgzURgoSTu0FeaQc6Yfh0dpDqYNAkeaTU35uTJ2Uso/C8FSDwv7iYXsNTjY9Zb
0GUvUAxwhe4jUrMATue1J21TYGIPsTEoajpUJQk6D63ezklQ41+kLOoP2+17cd8Km6XY0V8OOtS1
m+HTDfO01UHMsUws7jOAMvSfcj8823v2dMz/nZ+5mUXjpRHFn/AzJz0qaeheFYXNfXi22jyrwjIZ
7IBliPdoIyOWqO/gPL2le/Z+xROyYzKlKw+2Exadgx7sBdVn8zTqilX/7J0Ol0YKSA84bBDQuAVw
v6Xr0uK1HmWli6AMoIz2AHPNVdXJEIG/8WmI9sJRQPBpd5HKfP65QLQ0cNUa+4xQaKwQjI36p4CZ
iGnTgYAtBRFmkyBISF7L4+jJBGItVn4Z1g9kk6AVUSLNdbKjCsdcSnt795Paw8ZHtRhKsIbMi6bj
PT2g0al43GKJe/a4ETRpicI6xjWFfTLJQM+NFj7SUL9iqzCDNS12F8tLb/6F0XT/Czxml5IKBFe6
O7nTvBzkpdjzIJ8uLdWIpRBiBvy8slZI+D8KUMx9pIN0cOa6/LOsMsUAU69niAZCNNW3oY2hDR7x
9tY7Vw+jn/Vd2aCQJy+X4e1jDKd11psm09lQqflcI6fnBiC7Ki/xc14M9q7Yn7sNu+mHRv9vNohB
yPFT8r/ZnMAYMatDLoUqQ6X99RTd2+cQfwOmw6IaVWuMmPWWkKZ8GIps3cQEZ/EpqvyqbM52VAa+
RaS5/MyHlrmD6FpalVB50SDpjihh2RWtVKjRQi7KlGQYbqGRacdALQutCcrSicOI5mcuyxT+jg1t
SCllKmQ9wtiQfWWHiCZIxIWMcnGRUAhscQezXBG3+tgtKTsGhUZQPZ8d5v/z/vrsoMPkoD1m4B7U
cIimyFChYI/CL0oIdjsg6Wf/z2XaUwaHbCU333dip8h2Ke35KXQG7TsSiAQ2aPTz8mskTSHynyxl
Yq63NyAo/c4NE75HEOD82yfeXd+2J5L9AsT1kg7YZcqWlPrcEmCVGeGg5GauTAzH/WeURT3vzB9s
1u+F+0v6MRVUOOj1reRGRg5Cjx3ZR2IYk+dJhDt4vm6ecMuAlClI5WjEkHhQJFj04DehIANp0gpx
pq3NCR9qtTBskYXGxeyakEWazZvaaRJZfNVQLkyln+K5t4u3bii+nsKMKhdONyTU9aPTkq54DITY
VOZHALlXbh2PiCxszSzcbvyM4evWub4qJxFH3MGHcYJGFXVzQHf3XPGExCAS02hWnVSv8ptlBXrQ
Wv8ZzYRH4bLWgRLiieCjDA5+aNdc3TBzEi7BCNG6g0bN9INzxAFZhH9b1lCAcROfUKtBY0yk7EMW
lT7ng25FaiphKB4BQhl9bSd5XrRy4aKJRTuxXJugqYML6zEw1woCNoYM1ouIyympKpvi5ony9FA2
q5YU07uOQAW0uS1HuTiQzZwCbPfsv5PGNxFJKiNfSuVcTNP5UH50TCd+9DSvLde4UnvJAnhznoeE
1g+GfvSKq9n9Mn23EhD6UPf0USgC3ZDwnUb4BHCAAL1iUoomS14PI5YQ1r9XVIJ3XTTOTM317P6C
LnOufmrmG6SIbUfoWwGRRqTYefewK7Ej1xBJZpM+tlN6bKqCHX2oKXLIJYhdJ0PfzUyEViawKaNz
Ek8ccaihrBQr7O6EEHAaEAPKE2F7Y84swemEuqC2320KqIQajx14wKmXMGjwvT3OeUhDCECNx021
r/icltM3GTsLYVE8Js1425O+g+D9hQJW5cRcaEo0pb/cJCkitf4JoZdWKOtBme4mz3n29/6SNysA
4BgcBESPT7UbVIyHpB9Q5i0DJU+SpKkonfcVGdt8TDSs77bTJDtOfAuJVrCGAvuMYSdXR3JqUJFJ
k45uaX9i35IXsx0LmpeI8N/9SFbDOpN7DzLEU5Ee9i4Rgbc8u7sKAzoQzDNG6H+z7I5wLEgwHkj0
xMdyMubNLBwd/TPXwYwgIilTpqBEw8DZj3N8p6VVqFdehoOKWuOS4BytLNNIGlYBRzw8ufy34QI0
Ebt6SBRM07Kmadtsb2EyTPwSlRft40HPma9TIwT/9huyOpk7qvPMKmKjifUnjMzvfOzTKNwnhtII
8GrhGgf+1qR2/ApB/IjjSO2/xm296ZpFHghlu7ZddyNs1es075EvlD8b5sEipPm6ClRArmASyBUc
cMmvnoyVcQvwc3nnITafUPIdVjeYRKOJGWpFMtJ4hNIQ1JZkEusJ0FtFWjXvMjXtil8wixUaG7Um
dwkK1jf8IitmAk9XKS1g/YTBzi2mvkHmD5a2QfisH0Kqy1k0Jyvba7l1kzDlTZ/lRz8/2R8UMpkb
mNYo1DnRiSk7rk7dSkzmRPfPvWQUbuljSR49EinDupGXQhfysUCn/fivXehAg9xo7uINaexKERAZ
Z9VwNtgBsWztfjEUqMVLwAVYzvgnnSFly6pT7mAR+mQOa+Gfg1cZQ2Gf8j6gJ+HV05cARTPs0ahH
EwwJKuvV4TpV17jhQ/NDicw6jXlf3U9LiqffMNYdTWk0VCKQuDqGOMxyS8QbZfPw25onu8SWH6Xf
mcf+kfyh4kTCmr601Iy5Ku4HjXEsaqsUwH/qDm52f2+Q8Qe2+TyVEGN0+/Igw5glt7gRU4En1OmT
jErQ2rhlzb/nXPkZKJzp45OkbeqH/JZfQfWoUfYwWd1CqqKcYl0J3SLrHwfiV746EU6ZpRgWrso/
+UXvQcBPgadJ5KeQRcNkf/iJPN4QdWALtrdAs+WL006C8/ELNHx3ku8n4CbCCLVhx5cmuG1PWInM
Tf6DQCADK1wrD0mFdTeGfqrYQH31tz1MdXQ4oXfS3YMKtDjK6a1GAgS1jtQy+1pz9Gk/Kgcl5MU4
B3XIibqqqJ5fo5bxfQtoeY+3ZUx/gYWTEkonXDvCmryeXApHLg0Fe7rV7Pzfx669/LCBtcPT1nKa
SDRhJI1TuvM3Ex475muGYAeBJaSsEMbyTIzEVkdQhuEZu8wG/d2Jx6xjsEv9tZXT8BGDyeEv6GoL
1pZDM/iAHWG1b9Q3NX8MO9LZNpE6SnVyhEBuBPqVCuvE2/zsvL3AzBVSirxvbn5DB75CGeipj+fi
cJP2mWJbdLMUBo/gdDSu0rZHtC4H1QsYmtiXMBxQq/C146D7Sc0x97Ego1C2MlUIb0+ev0MYQ1pE
HLg+gXxayMHX/CS31cqvtDsKoylMxOQ8Km/4w+VlqZVTrPNejaBRScoraal3HxPtvXUQ32ScjaH2
PmEWNggotr6+a0TxzP8bma3jlNl66BnDK0Xk5FR/FOXAHnCNuuj3eOwhRLzXIos+0hkp0nkICCjf
AXBwGMNDLBO25Eyr0DNde8WBP9IO/QAe3Ziq9r9/eP91SF59VR7eFRs4mmIVJcuJJZZzDukFNod8
kyl58GM6fdTOzfhypov1nisW5ZAs1v+xlHvLlyPM0d3HWMD/Lzlc4A1fz30VZXuJ3nUiiDrBiQQN
xaUKslzQmFxqaphGdnMl7mCdTvNUHm9PJTrkG6P6YSMlfOkRVKa7OzKX3C/evUSsEmxyc9x0qLHk
/8U629kdFHOfRwbMPRM1sl15kAELRMEr82h7U38h9YuzAZDOpDkHaQrUgVUaNDio8nxqMX6AtMLb
ao9Lu4RQj3zA9HO6TOoVSfQWrb5X1e8fmBP+yVEGgp5T0a4Kem2n5fX4DuJc6mB1vxqL6BHUbk6B
RbZ/zSRav26MYWZjfVAnJrJPgZSp+dvBieKUv/3/+5+ORwmKVzuBTwKVdT5EjuwhGDxs/uQiHA9T
adyyFD5zjhVo3SK+JvKfpYPpkOmuG8kH8BUp14dZXoMlEtIddM2MLnUSySCp2pvdRUXyVgAb5yZL
VABQbjS7Nd2L/oSB6vmTZx/tE6MH6k7AT/XbIvowLVG1vXBlG6CUpWsrnZBtr2ahbBQ6qZyxY0Yd
Q4xpO/L9KrOuLUSxy54aIse1sUbSmWBVMXSrsWyfS0BG5QR1qsUzWbWh8oXpeFDINhY42QWwVUy1
zsl14d5nWRAit6hn68NHlwgPekGHXnc6q9AA4H+p/iW1goMTSk1HYnF1J/nSffh/eSmw/NOBMNMM
amMV5m3eR4REZ/Z9H4Ex2EcqA4Kfj0qk/CELfAYfzAHroufAkI+WOFJYKfSBIi8SLgnoSbUV1FiV
0sHfOv1i4iIZW3WM4BuME2CcH+KswxkqrjMtR7fbHVC1uy4/ZsS9Z48KgsAdUvmQyaeEM2EU9urz
K+AnkKADPNzUwV3NF7KJPU9rt8WYTx72jTniU7Iwyv5nkmcHtcX2ROHH3z3NOop7kbKiy+fNZY7b
/h43ovJWepvNpJpB3GRoKmMOtBx1ZhWtQZxdaIHDyGmDDqWvq4fJYKil7WyqtLPfnyvjN3Aqlxy+
tIOWZQP4l+QHK3Kvmn4a/lzabcU/Hf248me5X4MZM87J/IY31lefK7vvq7aT22Gpfw+adWPcOZ0v
YgNdgu4h+NzbD/ieg/lo6wyjwsDPbSnWAhAJfkBu6g5Dexd/uayqRi/5ldD7i3Aum8c70naiFMXb
u6LC2uVilRtpKQBwJcv9QdG6SgiExiry27xTS/uPIbJ69YOrAeLCooou0NbUiP6NYpZj/YHq11wu
VU7FL9HYtro1yBLSpBlo5KCN+0moYUr/1LsH24EsIK1RT05ZPxXhkXz/2qXexmiwEz3/uYqYQzZv
Nbm0mvLBSGH6cLs646Yu3BzIEoUdPXykcge4GAOilLEMhfYkH/lqd/XzJLYr7+JqLfQq8C+mp5k7
rTacIAB4o+MGcXTLI4uiqKrmQbKN10VBo/PfC78zEHCqsWW9sDvmyjZBkbp5c1ULMFs5J2d4vPN+
0D5uIvEkQuNJqisf6sJPFz3xlHJeuOvETAI3ny2u0OmT7904m4nKiWHRwTKN+FL/HMak0rElvIdU
humERCYq5qWPUIMEepQNmgZe/p3gC1xCYVjuyiO/gUFgPtupPSh39Kf+kELHdF402ZUBzalRJ3WD
gbuX+/U1LZcKucicgKKgGlaQ7yDSFyCetJ9Q1JIKfLDwV8HbnAZ7k8KE4mh1/VWRnMbQTDY7/TTl
5k+uB3tcqYl6IrLM2ImX2R0SwMZb6hHG8cOMHREWKVSDSLIeFj0Smj4C9ndv41k21TZlKHJh0VlN
cdVe8JAgW6Cu/BG39YxK4MA9+4obJxca25XOmKyYnd+kd2bjtMiNkkcKMtJftIkrqN4DQpfqQl6Y
1Ql+cayRrs6rll28TScKKlv7Ck/3SDmggGI8/re+zIZcrlzkVd1YfFEN+95gb2inuQI4NntJQa1J
5BaYtk/vxE+Y+JXFF6xDoumKlt5mkwJTOnK2HQXuMDwJ595K3EiWFl9NpnQ2aFSU/Ke4XmDqGJv6
KiK04Iks9bO1FVCYSm0YXCDjtI/sgit3AocIOfMOaAKzrNjuA+zSwXCRbPHnl2tA5/65oXp2dQl5
0HYYthMPOrgFB0nIk2WW82MWrjI+J3vbXgzsAg7IXV20bDWJnYDMHVX8luILpmn98zjYGhJWj0H1
JaBzBKvch90P5JkHruBbMBs2MBGfhAbbdwLWSkPVbcHHcFGTxNt/ARKI+luUQYel5suRvAHI2ed7
7H53/pb6ozCRgW9vy1kYSo7m0ieWMI1ywyB4z2Jdmv0OZnU7bJN2CUpBtZ/Jx7xDQ5Qjai2KHGUH
zmZ7Xph/o1K5oEE91KZcvKlhmCk1+NpbYmW53TqMaYDvNsV21yUpf9D2e6pbj6U5SUqUTAGM6Omp
6UX7rrzlScwvs0wLBsFt9lIfiCjdVqF4rVTm9WgUc8w2dq6PdCKLbqcG1suAGuBiXAwfL13pM7Lh
Syo23aBKqvIcqpNeMVNGKJOiboYzn59dl76c/lr1Ax1RfRE3c8xTEMQImzvnizI7R0yLp84cVlUl
U6vEoaU2o4s/3cHo5wXhk2tjmO9LiuXpYkma+etuYX8tqHNbeOjJ2ekwXC+xZy5nVkeQ72sHsA3j
T+7lCGh7zj9/uyDX88Q0qdloDmHbrfcBd8F2fx5YKOUvtuFiSPSYy8AdeG7al++/f23hHy7jqpJB
4+J4rbgqb1OnkCs7KB7YIx5ETQz1KnefWICpfh6njONQI+G6MBXt9PHL7ADJUM4xG6n5SJzQp0/N
a3CNae2W/Q5cMXRc5Ti0m7bNkqwDLgFohmQg6BrZgZ8AxkbcBaJjhUsWjD9giBcIr6IqLV29qWeZ
ft8mPFbAPnT7TZaAH5KgHAwLsqKdMdo7HVC14Pqt+FSFXj52xPMbu/Rs9lrf+kU4ooy59rs2wEcV
kvVKxtnJYZ7F0sHO4aHxEpDg80o9JUXkp2H2lGRH1AKMVyHxiEvH7nKdrXgfSh1iNtt16Xw2J0LK
MwJfxFV0WGzBvFHqPHBf6BZBEG2y9TNahU6PkUy0DxGHQtb7/+ygoS/DeUltX8N64cKzkMmY1hmd
BlQPEwJLj+lGy7zJVAQmXLLKozKt3htwWCYfk1ng6jbVSqsLceqJRoR1j0yMUW0tZoYcs+7AAUMM
jfB5B1/4b/91g+M3iMi+G1rLdyX3yh3UHsc6M3oN5UzD7lY0bnBrONe+Sel1L32uppV+JztPFykV
OnQlLlSJc9w7FmTmj6xsioJs6kU9n1f2cDH8332Ir6tk6Y7/R28p5B7PnouCWE4gdyv0Q4Bqbrq1
pN09UeA1x09RCpa03bUfE2JdYOKJpJCVpGA4WIx6bf0mOoG2vlcdttC9edFVrM6fG3Ai7154Gp2O
Il4FtfwRrDkJKc+2i9dq7YsXNx/OIZE7AwPqpCTL1hEzKPzxohEJXH78M4CDUrXIsRkyKycuVDbJ
2654C3JTNo5DAycDFs/QLK/e1HjkpXaTuQBnltS5aLBIWUteL41Qft31sQeDI4lKzU5PcNnm2UQp
2yejUFkckhRwEWLfIZ9dqL2VBcC5mz+FumSdaiEHP6sB2V4OoOoHekjT8BEtFXZH7TtMq3m7thgF
3reNKCnGCWnNjMnm5iln1mSh70rSlgblwyhiU4e2wfVfSL0TBEqvgXvV6NdgbAYwAw2ttT/z0eFc
5dvrKl54a5aQb57vsofl91v3GEiK2bOxTmg6hpinb23reTfUy+JMxYs91bEWPvAl6SzK4fumhPDw
YWMX/scDXJ+6a+YksTK4UDZE/wAaAcj0XMIHXjAQlIZm+uS/I4YsgQGrU1Zv9ZLMPlmG9q9oYohv
fHjBDvZRcNzDmzi6l6uMFAguCfv4JsrUKxI0vLm1OB2WabqgoVXmKSWyU96ntk6kW59A+8nnscrS
PhRm7V50XSbmJnidhTqw6vy653r14RTrZcWN0wd5jb86NGqO+nWMbwOz6t+P0PMlVqD/q1mNg0WE
4RfrLK7duAT7Q9V3AaD3jyDaV5TGF1vOehY8S9SZFHwBCESKhqjd2BxOZMELxK/ykc+bztFJLbbd
mon9QM7eABNL11uFe6Ohj+IBZ7gILFk+bQvbdGcsEx8XxQ9NoSilJaC1/xpXApe1RkFfGo61sn6h
P/GbsjTDOG+nOHsL+dPzbXH9PKoUg0Bby7GG3FdGmgdrZlZULB+jGs+ie6rB5qaJ0soCp0qaNCI9
jIR+x7tgj1C8xvsy1UnW14ZZnLoKLSicjbyXz2dyeooynxNFnJ3SkjHYVISFCdCw6AAMddFFoyln
3Co4+4lwGj4mzCDo5/LCKZSe2ab65jKbn5EFT+K+6lrrgDsL9yUrgR7/o/tE41F/Jp2fRhxbyoSf
0PP2oQHKy5c+9bGVP8Am81gFiCcMkTNKJwZFXK+z9utjsE7e/4WSrCqYwZlIuQw+fpISImV4qvrW
jfTBxTCXxBQjJ+yxEi3szew5Fr649BS8JfmWVYcy7EbltJbt7sUG5rsRxs5ADp6ChRLdg841MoUZ
qBHxf2wXP5vJ81yQa/N47Ag8J+t8T1sZk2J+0YqHkESrhQtaXAtAscwQfx/xiYWGtP0h99PLFS7+
Pi9tyXLR05I1iXe96kkgjYyJN4MCOs4RyO90EJ5wEkho8eLmRoytRr6xUOsqtMlpCrsq+WD2kp7f
SmGhF1J3cNtF4Mu5Uhd3becFdUzHRrE7U8pLp7EfOO78m5yz1flhRbHwn5GRHW/eH//RBkercDl/
dnsJFBkLjo9cob0F4j5rqpWQunqNFZnoxDjNQ+0BClDGXC6CjrAlUHp4Q+oi+3Qa3gug42YMhwIv
NxNvsTFgh+hvvSw0lbhyjnsT8FBvYUz6ylzEVAa4jgUpTcdJuTH1DLDcymowml6bwb5UvPAS1InE
QkjB1Lh1KImyw2F6QlENcJsSHQLvr/K2mUUqJJ43/SDRimCkY4wpqIMX/llDA4uibc7JHEpAIWbu
SqB6XA/PusJTwAtt+3PdtziqkDOhvpVeZzAj//OREbgZ3i0aR3LDp8M4/kTnZh3lWsiVM7GZM0fy
qrXbT17vPQIpTUiY7wsbDRXOqZlFbAavolsMOqlOb+M+DROjhfWr+4Hmjlmifqpk5TbqNQ7mY8Vk
BQsUnu1uDxzIxrcHSvIl+GYzGNA+wuTKzSUqIaFPW3FX3htEzWzIujEmkVjZxMv4MuKiLVjJKvQW
GV7jiEEMtqSzB8CejalT+5yfAk72eSak53ekL+V/ldpLcSFtSz9D6ASJPy+djd1/y75I6zd2Kcud
JtcJT9n99gFqE0ORf5mzoFbhHixm02zlALe3jZzkUaP+1wpEgR05hm2zG/KJnVfn8DXk7ARFUpv6
8YaYMwinc5wV2AAkmnLSEQSRKOlJYvDRSurnQSeXGURKgbatQOZTHBBeI22rSKmsbXxm6wapypgr
h2mazXlDyXLeXF5me18j/3qGXpxX1wpWmdPZxlKPTWt+IzzOD2SVuUhMa8cQ2wcAY+4yv+WC7DyD
SgX8Bq325o/1ZiZ8ZiyyECPrgcgYfyeEbHN3ALSH9MIG51Tdr6YoI2WYD1ctCNMFRjRgIqruzfbO
X8aNs2DhdI3/7PLsv0JbMNNHD3nRlpYaot8aLZdUYwdffhjs+aBrJ9K0SlarCvcHaeIYTpMeCcOg
zAesqMF65fMR7tAXJh3kRd20vbmHVqUqA5wfQswHF7CmP0Uvamp1X6aLOA4+7nex+NqKE9y7On4Q
6/Hc0VA7a0iIZqGU+UOCO2td2kVEH/Cifc8HVA+FtYpLpG41VYDKgKcuR/aAluTHYTmCuhKx0+aW
yHhcEcU0lQTY0Dq+UWJAcLXnJcx/I+4Rulyr3R0HDbc5udU7AmYwzAquqd9/J35YKcrKaN7UGjP1
XF8/DVY3d+Rtol1w9wtkD9ecds1GUYrHS9Kd4wGC9LWhUg4/xStSoMGuEpz0KeDg9fonrBZ54H5Y
roNKl6lczaYKg6NeT0aimcFpL3Ji5Y+5/c/OVvRMz7xSkpP66BIUAoYXhKIP3xqNjaPzstB96Bag
TpKWAyEZeep5Hv7QhNuXAKNxDgze1so7gR/U8ZTP1XhFMqCAxjSw+rHw8z9PgLDs7rqobd2kQklv
v8E+hwCwgQ6r0vXpUgkGXAudhYwRirJ3JFR0LvolEYuWUBwWzs9h6T9ar+dIfvnur+djYQVu0af9
AUAjXulFY8DKIgbVEPS5lGp8rK+CvJJuwkB1Vb+lRVcYS9xyg24fCW58kAIdtR9lQ/dfZRgQxz+k
dmqeaeePJM/m6k5GndpasaJrD8dIsCoKs3ZEYhTB+X01OJsU3P7IXUuvGXyT0xT8922B7w0p2y5T
SWR+cU1IpAEAvCwNe5wR9GxOmgtxuZZTqyWw/Z748lVd59FD1+lrTVp4YdMPMU69dIk35x6Nz73P
ikWuCdjA53G74gJ4BY9Lh1rqca75CgnmYGLYKCn2ACJKCD7Dn0UGJxK5FXJdIEJN9Lj3PemOfkho
8RCCAtQL9JCzTBTrCKRQmfzKxsRuCpddz0zt/jwDclt1Yl8WaUx846zmDTNyHqTnfUS+Bwrjy7US
LMdwvfyqENEiklvKfg78wu7kwYYf30gzWUePC2ntC8gYx8ysMWEdrUGRDIzGUH/i3hnlK0PHVPwR
L+ym6C6pYC3p0EsokxAt163FKLiCdi52eip6PheMNHM1HHPEjrA3UQ+tresMniTjJYy3ZkMV1yFg
GewLh2AMAWHs8LKLzDgTw648bPjQIoAaQPnXJoh2UnQTqhpYNN0/PfB3mTIEsbgeoyemXAeb/tlH
RuNL43N5h2ytom4Ae0iOz/nCwQDo8rwokpEKxUxyAMl2CM+B1zi7P5lrh0PdZdV5TI5cVJCwTE6B
GDk3v5T73y0zyCxTwVXL5sNLdk8T8vT0V1RhA3jk96xaUkOGkLthX3ffmFyE56nSE15jhJnc7pXF
Sfvqv0vYZ0wyPMdi3cQP6A1Wwav1HysRU8kWKVIYnjjV0Dxic+vxzZ6WC9OEXoG9KEPSV+uKMzhH
rsQsNjXXH/7fQu88BiR2ub2RCRa/VrSkRqaz6b0CNBMhzU6+Clqb20LAVvYVtfZfpHPqpem2EV+J
DGePqdRtHwiw8sMhC/9XfP0LgPXVFe0mgmCRBDm9uXxybBDt5pbu2TT50SWDZ4D1hK8Rr2unlwBG
nLc8+iiYK8q5mW3E5z8HFJ3mCY9lk/zecSSjafSb+tTEwfm+296FoRYV1AS7CgvInPlKenoa3Pft
7qNGGfV1+m17rfNSvbXzp3eqK6yYtlZsyzIRvWwg+z1sURxSFsR0D7mF7mRq6+habhCfYxuk8Zhr
j4opUKjfbilix1pCPiNMpljWgEbcl4X/vU2pwzx0BNlFc17nfSKOVvDGNKu4Oq12noPl17vZfe8q
5eqIJDRH+P5B6uA1T6wx4w/2GRya48LwND8IdQ5B/LgpcKJjUh6JrUnfkIPBvCIYgFoaKk+xNFk/
9mQmEDoIrFzyo8kegy4B2P4bVq6XR7cwuIYxdWjICi0OFtQfr61phcB56Q6eYQbpARxXVOCY5DEs
LZk38pl9q8HYzHUYNusyZN23pG5U3Z+OeXSQfXcdKy90Zimtnq+BiNpNeKX0JyD/qL+Bjpn/YL7/
5hb2+cQMa0ii+IWYzZR/TTT4PP44L2attyFDs7c2XpMnKMvkWMBDyty3fyvutuD0+EQ65cP1gec+
G4QsJe7rfDtM6gnqSsbGFlnTunOuccPO6gm4cUazZQphfIkVpGATJDR6NFDIaiXC/vRfbApcHUPY
G+/qX5j1oamBLZRiC9LGP92bwi1tAH7SrxuvSeeRSbfgCGDqAr8WXAjmlI++I1aD3T+nxYFytBbs
jzsk8eUkn9B1snAd7UCr+2b9RcDTJZX5zDpZAC6s9F1jSixHo4v6SIrytpENq+RJNqdR+4dDCaag
FpDFn4ybrY7hp2Cj9X0LEf7Rt1P33RWJI0z9oMhNtCv4FZ8ZIg2S/Q5CFw0VuSOUwNsgmZeRARy8
/yk2vOixRm/NJPluf6gLt2mycVLwVlA1x79t5uxankhKE4I6Whvy8EkQid09mIJ3deaNK7DkJMvU
7NWem6rBEJVBtf/n+hO0BQZKskHDFnteIk0X0gT029fLAYK3vH2kXqF/e20CH1bNckv0yZw9KND2
acQzKl5tVGhC8Br9oGLzQUJ5GaUA6xqvSota5xleEXWYrcmpplGDaDXsYGa8voOaLf2BDhUmOC0k
2dQdgDE0h/1NBGr9I/SWWeKwVJyeHCbQTN921hoqPIC4Dx9M/B5L7ZNZ9F+vveM32UPYAG4LuGxx
HlvP50Wbrt6qnlpmKFype5JsGP83WaLCFLISdSQKfyLRmKhYTTY9J91EkqtK9N9GA3We+nW7E/os
DZ1oRD4sgfkXoJKcGKPA+ZsM8QqwY86WkldVpnGfkQYHdBzNqsuZM7rl5/dQhH6jigPG5NoIWo+e
rcO3I0/y52dNlCsmHa6FWIz8TsIBYlc2yyeBIrNiJwuvT6wHjJVVBUY5Cne6kyxId5Li/jDfXiaK
VlEeKdGf0PUx+fUy63g1rUSw5pgRVpfN2Xy+FGogmLHTARigWEmPIu5P+TG/3W9SzheZy6VWthoc
hkEC5ydKiqFKNNz7uBfmoQ4oL/d/CZwUflWHF1h5OUXwBtbpZiUyX5+NR+da+OduUUbTKEfGJTe6
o31GJu0pZrmNAHyeg3TEAJF1kGqjw5q1D/t8xFAb60AtKT5V7MbHkaBN0TV3IFuv2obW4MfQQ3Qy
7qpfqsrGRO+v0DFyBqDWLyZxftNgkuLB8SanGtvBmRDBtHfXr57Y4jg9wxFJ9ahALwyTiCH8/GJ1
Wey2ipzQuAi++g7FobmTBy0b8sy9yp0V9oVXJ7V8CiYV0FS+UJ2AeC8i5SVwhyEk+oEAntI74zW4
7NR+bGDyhDJnFx0TJJ1jbDjiMJoYzTUiW4srC7GFvtoVovcbG2oBB9h5yBwU+zx7vKEvNlBsgM4W
U1Q9oBbeG75OzvPZi5t4ORCePERLN6cVPXFcn0+Y/Q8eFH4Gl+nQSCdHM90+d/2yyYrXL/pAW6tb
ccrT6RVXn6RbSiYSJ7XlCAsUTvr4wNkKWn6R0Z7Zfk40N4wB5roFn6KxWqzC+TjM2/SkBZu+K+7O
YRa9kA3Jfm7/RafAnapDR+NgiTK7967k3ejy7gUnJIOZ+GIn5MaZTzpVNe4gv26QRZQU3UwnUhzh
5JY5csWqT3BaxGQ7us4fg0dFBnU9PG/kTcddDECm9HWqwIZcOzRv7OyH99PPmYJYREkJDUuxTfnt
mRcm2DsiWWBqL3vb7CQC/lvTRfHKlrV5naiRa6EckTiaxgV/wlZCRClzDoWN7/2bB/01c5v6GLY4
FkqZqzMhT06ASuTHGMCttk3EUCo1JKW5Qbv7e2qvqN1Rtq4NXqf24sL60RJqTmqIDXpVaGH63gQN
2pr9fdW2qfOycLKOgFexjHJu9VPvzdKnKvYO8WPYWnXDKT3HIm2NkU6ld0KP7T35biCyGmg/KVe6
lfHSgemlUtqW09Fl91QfjdjIMrpH3DlJr8rzFRy2voi83B27wI7Pldc7j2/6tOYtaBdkTeFA1Xxf
wh8cmeVt1W2MS5u/ClPbBV+1RFxRXlRZnpJXckpahFZa2LWIklWr4MPDi5f2Q2+PuGwaQuAE8NmQ
YufVPD1TNsRhrsUoOOynm6iIm8gkSNdRYusAduTWdoifVfU7VX5xcB70ICvktwRJybDWShwivK4p
UM79jhw6HRucWO4+ytZ5fjvakqwXbwZ3HvU5/Fr2VAehliAhjfVxyUDo2n8+jfpooNVFiK9vKq/i
W8x3zWzDZ/f7fMLcYIkdHfyhVFAZGWYuJeOuf/DG/YVIsaUYqO268AdANdLussm1OboLqwZys7aV
p9gRK1MBJoWecDsaikzty3/Xv8VbGnoBl569qNE4zT64vRKf5mBZrgft9FHox3ZvUXcYB31cFvJB
CI1ODdPW5yilEzs1SeVvyLe1uAzB1szh6mUE1pvUX6PCCQULiIPCcxMGHqnXMGUwELxlHOvg3iAz
JLruQDvKkjU+WYIAvVtjAgtpQLUAnSzpsK0HZpfdYTL65npDYBkEuceh1WQvZma2VFXjRVs/MAE3
+jX4LIZVPTJVhNXDX/629y1sFSjrT1iJ5FjuoiY7N55KBHRVdLkYw+mWWA34s1i3eS2COlm1GI5/
wDDwuH0dl2UDQX2lc33eLZH1JuGGjNx4YJTvo/Vo4b78bBjuWCfXTD1QIS/fVm/gp4wSCsbk4e9/
+SVL63rTyAbSImL9b8u2mH1IjGiCdqji35Wf050y9ViMcwA+xHuUAD9+XwLJMgeZyOKTLWI8uz2z
yMGJYkAWIq5ybVlSFjlDFypnECeTytYlvbaW4VoqIrjOdWbvZOBomCb9r1PS0jN7YW7J8Oj2diuk
Y1SOpc+kGJ7QTgvHnr8Omh/KPr2hSWnWI5YTHJz6k1A9BZSkyRlV5pmI430ysZN4skfdXpDFUnUQ
aJXDC92Li64I34JlhxlwKHhD2FdnVxSpTSBwACw19N1uhFON8Jmc4DeMds7lNDhnYtkJpleDeOh7
OHbarkJZ53CPjt38KiF6D7ps7VOmM/R2PkuGrxR9C52aU7WbdcS2hp0naSvcUo1bCpfVUDgGJZ78
wczUv6x9NLsN4uynh7kapi566F93WlYUBz5rIwiPhJ2HPPrncnyDyDfqCg6RU5U8Dmcaity0Pq5n
cIe0ehd0yDdtvZymcX9gNXYJ/lof9tvNf+0WKynqEusESUSff3VFF8TuZIg1Js74WrcLbzB3UPS5
h+tpwTM1oHzUM5EMbZ218PUGnHbTSSCLaubOpp+wXTUrnUhRzicvSYcoPTlT3VNHRuu6EN4Qw7uS
M/NGBsGM6wiCouncZ5dTgwoCqeMWtNql1bqzKhyKNbS5nLvruYmexGctTDSNMXWt8vbKbuJalRn+
44ubWCOiovVY0TVGD/eUS0hdiYBPnv5kbQmaZ1dOolbamaf/qa4BsIgnEG0zm+7DxOOV44ssh5ZV
xTla10/BHo94ysNsq61kNsIvA+gO3eiRBI9Fj/N6qjlKrCVj84kuxGA6FRSTRfKSeWoIJFVWDADE
LdzR16nu3xpSDiZ+GSQN0rXSuWjFDlwgOSZCAllu6A6pixrIl32xA3bnlSEPSP5Nsw128K/yFKhi
74sK0Cl13rkf/9J8h+84YGfSRyqI7NqcaxY1Y/ZA/L6Fv9nvZTLH95qS/gseS7j+U0VKXeBVfJOB
fU78yZwnhh2R0mN9Nj8d7l1bNlPlxbSwg2nXaOLc8Mtlch9ppJKs4vE2uqC5G4FnvGJg6sXtJFPW
T9kF+eacd4MMALRqiuDvIuKiEBu2XqgD2itTeCXsDko0KqZAcwhj24VMUPpB3WpjKrgc0/I35I72
QevSUbt2aotlKzaW6G0CCKIsVo2ONc0pgjeqCkDoU6FFcCVeYgbHxZVr0YIy6rX5zygQ+fqTfI86
l8v7rA1Wmi9zUD/7h5WaDuLy4NELjsVsfQGXhueY9V7NgYSdj+qLTUn4vkx8F3n/54MyO5gq7Ax2
DrOaJ+ECTkhESX0weXf3cDPHOXFWYfdedQDZGenMSAgJF9OAYuwv2sFTPF5BDNPUDroMFQ5seoK1
Mn24M0NyHaTp8GCTfRtuH2IZoLMpNAYNZB9r45JasD5w4jMjHMlgJQoIiKXkkVBcI6ceFHLlXMqU
Y0I/qlmfVVmYhfpJXfno8czjhfLKDWXT3ZCjOJBMk32YujxF2Ivd/qL4n8h7jxIXjtLZ79/wsL/R
J7L2gtrlo/chbZgPeRGVGvKXmWCT1uglxuk93v8MJq5r+lOVn4Io3DN1zM3VcuTp+o1APIG068oZ
/uDSjIViNyUjcLQ+nIDJJef/6I9a6OJFlJNQeG6LuwxhdQN/WwbDeQviC6rTXjdgq8gXpqZkEGsX
CoggwN9ZZoUq5NAA4pGH2NW7DEE5VsFiTzZofwP0siJs2tNvR6habp/OUtgTubWZlD5B8BJCmPNJ
xehSrFvtOXboZNZOnafTqfUyHgYm5epT1quQDdxo5u9fPcu40uf4xU89c8DHpv/eLQHnXm3rj/tt
2El2MNWkc88mwqtpWA8aFKMR0Yde0QAjP/5r+OYWnVcAl3PehvVvt/UGt9PDqZvsXVtzdEjTGIpX
WbHksl7HeS4bQz6pU9NzbIqV+s5oTNsNambssY8LBW6cu4G0Q71i16kwg2QPQVg2nrnxIwBrd/MN
5TqOG0altRMvspxFZH3Gc68DTmG56zqlSGwS3x1wf+THhJcqRRcib2qPd7yj5BByrcHHBWDT2UyR
Q0V6Da8CTOYgSIO3pzDDztUxSvfWoefi8MAogGpCT9RcROaoqXnPIthuVaVKE8Uv72/joKVD84XZ
7bKcCEfDfoaKkNXZHxd+NSRLNG0FoGSa6Fdne4bXM54T0PoKx3F8HM1A2SVYHhGvYjNUXmQFR78D
YX0bXvEVDeslrQOa7TrqHpavCBLFdXRQH3iOEyIurUIeKbKa1bDp0Nnvq4UFdd/7xp+O5YTmGH4Q
vR9h2f83CTiU4W7tYJWslQSFINAxrGIG0K0O50QzSScyiSeyj+um3Y/Ec/hQvnXWXHi6UFUIQmyX
RBxy5RxEeIlLL5Xf0Sggpis9zFNylMgkAyCWY8Meca5kqpac20Edlg0N0U01LoROws1XOP7Tlj2c
4woktTTKxnVjCo9GjC4d1oMj2ismg3CbaH444sAfin2y3VD/VE+jrYjyE0sQJQZMSQKnCK3FADl9
EATvNpgHS5O1QDR2LIp21CyqzvtIzI6djdcyAHuwU0cX3CmrRzAU3KWu91+PNUQBEAxDZ8axhiJK
OH+Zutgmm55sVRPyj/0o9VC9QQ/KhnqIbzHIMGkYoB0aFq/ipedPJzovaJSTPw88+oH1o+lquq0q
GnUDQzJnxOE61/ei3t9iM36xigh82cNyYG7f/eqUSF9gu4p1Lchrn6rrmiDLpAd07dnN2V6PlyFB
r1TWc8u72tDkJQ6gIQ3cm+3p8OGUYKefZ62OLtUcBAyvzxInQEuDa2xUlBssX845U9TH4YBuVtkH
+LqS6BkXrwS+R8r7PDliMr052mwdQazdP61fWTvXuQTWaL0Nj9GIZUvGIKvt0+nIGNGI+pys9J5k
5ipm+0cCfKiV8n+538D5opf7W18Ui2bv1IweSltubkW5h5aHUrqSB7W2ML9mcgbZdi/UxjCNnqzI
U9RBvcdqzBhcBfmg2xwYzqc0opvfSR30wnWJjJL4v4oybihJ1ARdZPzk0gLlDTQttLiO5mswurhg
ELI8IEfiHuGO2Sn++1PsPNF3r3a4JPpTt1UrXkWjQdKeWrLevFtK83bmNOKEiD5K/jV75V2PMl0L
013/nN49SocEbvRRTjf4498YKa8bGbawfJuZiq4p090DXalj6pTFTyilXl+G5t+amO8lLtFonjtX
ByKBJem57Lrceu4sXHLCv0Lg2Z8N7Rr3rqG1CLtEBt1vtC/IFoNNWpGFFS9X8PeJ2fqQ0I7qGGao
283Xo5J7snvSjKTJlSWosnETWtNA3yLReFGvMDLL6FhaSy69tVhKjYjUdYWM1DwYTREH+zQN63JG
C+vIdmDiJ1NKHu/7ESHZtq+4MhpVbExT/ratOcoZSw2wedkJVjIcWqoz7G93PotforZeH0hcyK7r
cqZJYgCL1y0rf9nC5WJexxACQB2LMWISQA9WjPI1bj0ZLUy1fGtviA0rFe9l2/i2mH+pv+HrmsbN
p7sCVFwFXBsIhIOKwuqyiNVK1ShJEXkGYto3rGMUqOm7NdRlI4uMBiLGKN/gTw0RguTorPJdM2dj
Jk9Z9qUQXiZeYa+UvJNlRXedQKuqWtamHUEeGBAuNL/kUAzj2ZiIGmRKPXi3s6k4pkDKgxrMv6gP
VfvYY2rXYXoi58Tt2cWFIlOV1PfBv+pvF4nwsPIHp9BJyIflx1K5pBq9OqLaTU9c3LsIlqB0jm2p
FtwouRVPOuWjeC/H7tYYybrBvchnqxKjsPvPmFlk2/leROWqsdzZhW6yUbkpeZKLrNi9KtSwP0cv
WKJmbbEq6zC7EEW5C9h+d5yR6ZWUs5pqY5VQhZbXPX3ojgh/LLzodEwEXu8Fjf5RruE4gm9h5/Ci
UG6SMP7riSuejGQ1E8/Ywgc9xESOzsw16vrb/cJhx/9jkX4xP25W5QqmCFzYU/MbLxIjgPJBpNpb
7NWLpYrNFzrzb6/FDVX4M8vH0fDcu3pBFETvFURtDR8uZYukAN518hIQklKVbDQbkJGEFoX4nzQB
QyJItT5QA0GECoIR0XO//0Cxg6w9+MOvLe2srmkP+nfK3N70yoHBEe7Id9hJEzsUVKdXcREGfkpp
f1Ylc+QLoSBv159iFE7mbyeDlFaqTPZLczeEJK2xzD1xhALzXBnYbXioW2oCWi2Rst8ILF6THz0q
zh8OglvBNc8+9VDxrVLU9Spid9q/daTJdHevU1zlj9Wk1putS3PklmVQMIlESEwS/3VG3e9x2W/e
t+ueJkNh6sAwzBioHfCT2QiN+VyZtkkJgz3dBtfYWq8O+tTT2bZJvqxJRTnjJGkf748ziopDryOO
aBlfnXY7YHazQBYFptrTxmKj10DjIzhUDl15yHA8yGlDGO91L+R2zzdf8c/cPYh20i7qf1gnRG1Y
KJbm1xw3ooLd9jH4hlXfjGnvvHK1GuQRZPg0RVCD0qTqgT3kXA/QNgm4t8suFBKWUD3Q85XEYCnx
AWnJDLR1+Ocn/9s5nqWyIaKkjGc3+mpq/SsF/vxvzrZdZ14Tl9mMfwVSuStmzoPOS7qwuZucPIoc
JJ2zcBN5UDzrqquZc5ywoSaP6sjNRjs6GqFJqI1JR48IAD7i8aba8jgKdqVzWdtxTbS8md4xq0Lb
JXsECOOtKhkGV1/8OUOcruHw1WHvm1AxUGdw+9tTREJjl6m5p2CP64ksPERQFKFLMaDg2CUPiwJ/
QbIF/tLacM/+PtstcyE4Lzbrv5hDotUYAq0UQGERORxE6mV24ztkUocGhZws7p9NI+igUQcgt2WJ
H7+jCW8WvSEoCrWZ8ApbIdTeyHD1usjpSU0D8dCSjslLD6gwyh0qcJ9mKm2nzy2d3Oi7WcvoGaLr
H7YS9ozNVJmBGAmSnGaCBiehES6XMDG/SL72IjTG+wP+bBXqrG4Qf1xUpdxdOvgRpbrxEIeZmtea
sFC4tkeZC1PUBJMOkmABOs83LmABnRfMXRotr8+IkzEbYGmbciUkDV94WRxERbZwUvQcMQeRST6M
w2vS13pQLQiUw5TZvFn/tfzeXt9C9zja8QaEWCGu2WgtWdh75p/dVydQ/yMWNE4kDwgRLyLwZcsZ
L4VYIYWt/B9OSVZSS07IEsyTopTakxa1Ybw6rBlSlwPi37lTDnnsRo6GN1P1N8cVji+ElbqoM76Y
ip554HIzgONfdVlQ+WFuHXU3TqtTAwAq8wibUa80AWa+n96pelMWLc7nUUNkf0VxfA8tMX/OxuZY
usMUE4WV2ouM3vLAJj2mXYf6u5y/XgOSfQwYfh0gegrBE58GotyK2nFxZL9VpRbsRcplm+0BIVII
U0FW+lXTC4cjoYzT3CxARTMpDJqmoIj24KgAY0ylYwND4YCoTWx6BSWPkxIrq7bM+pn4hOyedz0r
Bi/DUcyUa5KJF6tbzH8AiJX1gUUJyWQ40ehc39uWvPn3POVTVs5qW6Cjnp/rrSXXHpNiNl39ebOe
SA9AtlZkKSiW91tn4fv82XC5DNlXI1fe8JFiKx0wWMHBUstiMTHFPx2ZWx/wWIV0Fk4EsbbYSBya
lDg3DPLvarvnfI72C0blcx6wu+6xKgH6BgVa4tDH99d2aVO9IwIIJWNVTmVua+F2NYFYLdBMR13V
T2Wz4iGxr5uaKZ8QBYmgApVe93aTev40Lw/TJb9j01bHdBvfWmGgazfV/WeVjMQKzhd2Ka6a1Kq6
M3qmyMURzgd+oNmYgqQGiL7HGKDgiPy20MCrve5l9/mX2FYOGS2ydElaHoKuxa23JjPLsvxNIYlg
49vvO9sYp5MI//aLuWSke7j2BJTiCHZ6bNmScZNy1TWXHdeywMCRIjW+Ovt+GaOJUx02zksj8Aww
Fal92O+dmZm3DrFCOFrpZt4hTnS+jydYHBgbZ+jxa9nR3teDARBpzv+NspCj34fZ/lZvYPAXk9sK
Vfvop2qi1yWs0pIr3V27fwCI8rjGkTuG6ACrGPycBLrPfbgesnHw/B6jvUkSeZnGnU+k4ku60XNf
MYQbYD1g889q5BQWSq5K24giJucDKmp5x573iFyvC1QLYx8KpeLxoYgYmu2wL9ea94mjAHAbu+uP
PTsJKHK8xEAEbedAce5joofUWIpjeOimZO6c9KQTmEq3774CKC777D4uQDcnFM2R+/59NtwiszaU
oNVqC1dwh1ZQL7oolQp7ELUmzm8az2da0VFNarGVFXctgTIGlvCiQN1lUvnccvvH2RmKW5vIKeCw
sujtAgKt0koS2Yu4EENZj8/VuDMJLMIy800NUKmvZHd9ZSo0S5VronY0KE6POH9QtErnAXNYcJUz
H7StCyOrCqF/2tJveojH3OI0xjVTHKF7cA0LOERr4hEB/YWP/BLBxV/bgVV3z9YXd8qxTQBQJONw
ZkkZDjXco84jLnYzRF/U00IUTdphVvCna8o23y7iCVbiRfNoIsVjbKTF6AS18NA/DtSE68OqrdpX
Ca/O3E7LMN2UkSkucxMLrEH5X0pWpX/QUSXICjvcuF8xmnu9vaQH2v+kqNHtfEFx04uBRLzWOtRY
505FRmxYAwMex64ZM38nIrIxmxlllOl2C8ECyQdpsz+rFqMmmxo8Dd7JYYaZlu3Yb59f4yu1UAdX
VaajAGTu4PLhHbHzxrZs0vSf25RX+eSYQwGhHXvvem1ppAwvkFidiKSFyC5imgSl61VTEGzj77uf
B8fHu/Ul1zkVG5tWsWNhmGis5Uk1QW2rRWU1defNW4gSla4u37XFzxSnRnrtop5kcBIF88+hAo4F
qO0CDGIxbvlK7sH4yqgpPLZb5oOkTu7s/KGgpOfAe1pmX9attfarVRu5wXzEI5Zyxl1UUxNh810X
RMir9VLcyWeGE2XFen29tMumEDAeQhjkQoSpgiY754ri337NBsBEY51Zp5jClzfOUCXHNkZkZwXL
cUCccPE0cwpgQQ05LM2qv1yZXCc5Ieoz+0ngkxwGsQd6KkGWFjsXdEzVuuXPw9QeowfEe32JW9Ry
vsffxUV7b2oiRgk/jNKLA4Dc5aV8W5mPLJqfDvkuwHRbc7GoL8HVQFfoKx1WsfjyQgN4NvH8+ZIk
ZmQD/RlflI5lsxQmzmjujIAjQCGbOQ/74VC3M5cf+ZOdcaqsi02ntWcp56m4hpY9a+hURgJxaDZO
3CPXBwAYdOfA7d9RaIMTu7gYt7sxZ6xdypKuDuvpyjR7WOildMrIW3WPVB4Ds91DAM6cvDV+aKHF
urc9ook4GDj3OzMs6HuS5XckOv7AKc5OXXBNHwTxety8PDeED3678Iy3Tv09Tew3surxgo/bZ7mO
J0RPKT33YAl7sPOaPNIQ76SiMckEEH7SxKewC3eJNnNfGKdx52Nyp01oYcv3t6pxjW7/blIfOTcD
kSWETUkGjs1VbAzfvW1+orqbeLQsFD3VQWeCwbWHGKpTNiodf/jMk6OboWs6p3SQhCKZx6XToCum
EuQYkz5oSdFUD/GYtk82/i29Rt0u7oual+ROi+hP4oXXnlrUF31lbJtRBlOmXOM4t6VYWoxcmPkU
AaHDCjyHQCOXna5GaDUvxw7aS6CCGGyU7k4LIDcTsjxFSKBQrlKUlDC4WVxEMXmoJV4NfHvRldKg
SpuVLJdOZ8oS4ubjH9x87EfB2YAxRlv0vgP2cvp+AYTcAOB5gx/4LPnkOTf3thVZNSYcuExPk0Gv
fkVnwZJd6Ktx36IJkHx1WwU9sadckc+DQWLp7MkRjENA1X+VIEYxHPh9g+gzW27AaNC4/R7zSIf1
o1BAxN1dHJsaFsLZa2krBT4rq4PvAWI8TF6ku4IVwMILmLirIa8aH62DxkbrYJN87e5LMK1+diS4
tSeaI9Czc34c/bRRk51IKQd2xN+wY/3yYLGgQ3l7H6XvoOLXAMjFb2MgRo18ZGvYfgjjU/ykpj1v
Au6T4AmXXfB8B/y+FQTwlkcmlRl2Zr2FX8iBCI2ErNpoiFHzxv5DuqqCTeYppZpRquPkHHmmD481
AYvLBlZWRmWI6wLFaIEQP7LkB4k4sGFIZ15eMF/Htvd1+yuYUIvxq4Nks0WXr7DR4qlEnhdoQ8b5
Vhek1MFwMZ9AME5WqGT4y/srC3e8EjS1f60A9vPzopnF+dJI8dezP/uJieB7oRgWtovZ15LAOCi+
Wre2E5l6cNFfDy7NJYMq0nxnF0aYZm/kDwcSRkP2x1HOs2unpTohXLceADAEGOlgQ+oAOr9JuL66
n7EAQDq6yCt8JIg70HsZbToU3pN4KH4jHr4fYBlWcdFmHJAH5szlPU0YBMR536C4diqbglpnlep9
Z2zOY8bUKi8JrRQ9bjMkhu5dY3zBd/kxrZBGdA2qZh/m/cFJNCFnGbxi4r+etG+McYM2gnr8Zsno
/qIxTkT6gFBXMtuitMSCblIehf7Qd+xHu/kZTg9+KtlQQTAs+imUCFnpI6wDSiWNaSQRMJgUDq/E
kFONvYT5puwDu8UqxSeI8Lg50BuramDFLga8LoCmctQBTol68sHqYoXpVg9Occ79EUp3A9LSFDG/
t18BTZ+IgbUZ1wtK/9eG50B8qNf8sVJMQx8+EGeDWBvpQB35yVgUhxZAeVuOmR5KA4eUYBVMqOJQ
XpWG0B+YL8T5hecKiEMDs1hhcOWSliADSKAuIHwHIahmwBSbLw4Cgh0Uy7fJh212R3e1sJCBSMaL
taclUNSbfDo6If3Vggtlimb7XNueMrO9Tdq4aBc7pzmYsr/NDn/M4ifoUIp2n6/RfreEDABCblje
6HBcpMf+cMh4xcUxSwiz2uO11c6QOEhH5M3QMUQ+u9mcR3/cGDzYS0rfQnh7roDWSs4P3NYzC9Mo
gZldU6atUeAqdrzL3MEi2bgBrNTfSmuOxVshgv/uocdeS5OBR7jfYvGREt48yrQINtKBjLimxV8U
yN3C5lWEYT9IeZHJsnUBK+B/9V6wxYUroCIWDaFxP05mOXEfnTjrm6tbvmcJCMD+6rIImecIxIkh
Nz/hA2KZe2u8ZEE7V0G66gkslUV/RdZWtMVE42GdXhzktzfSb+0QUl7QBVN47RllVZViH02l/omD
1yLln0ytmE3Y4FWMDD2j0bSPAgTDJOZutDvwmapPqqbiZ2xLDa7e2LDN1RdsKXxnBF+wgnS5C4Qy
iRzFeFh/f2BUiomrWxaRMTGCMrDuuirfTiQyq2105yjt5i3i9R/4ckmWiyvJFjCAyuYScz9QGT/P
qT5kuN5vq04AWYOObBQjVtPPjI5BZTZq1hbzjNph1iT+aclnNWQuX7xAWwZFApqr3sIZmB4ccEHz
h3/APS2yxIgv8yGjZjxLEI/NpJUbaOFuajQKUGV+ZYYlWnwT4j3qTRR7tWRMIXiI8JaN1AiaBwMv
RMATBuO36nEAR352bXLvh03+/H2XQH0G7KFpBznHOHrZCSp82EinRXMoQIzRBHOBJ3aM5HwwnFCR
UPm6nxoQ4/5185Dz7TMrecLp7SLBedH+wCc5u6SvaF/UOynoKyQ/IZ7b7Xq5xKc+8AJrhX90Cf4V
0hBZdSGxWppnCODfMZkUDpMycvBNXrWuaDTZaWmquOK5EEqIAIGEWvM+zRmYpXEjoQyfaokGT3Rt
Xjm9wGqZy0gUzfMeBo1D1IAzW5cvrb8MwCqeH2cW7kjes1hkyREZ8ccnjqekTe/Ii/jY4nRFEXdJ
tkiTAAracJtbQ922xoKRaK33+LizAJ7Ni7oPhth4kGZ3hXE2+ssw3WD1njcRjUtXCTlalz9BLePF
adND3EfQ2XQtlHsJ4VsnId+h3euFU9QOn8gmYV+ER+Dlwzs6z5HnW6rFLQv/DD7QNVwxeoUBATBv
4aEeF7BBH0BR+yRW8SIVeHF66vpUkGgDpcdY8COQFIyD2prRWZ6JfJkkRpRdgucAJmJgR4r+H54+
JxTkjbSbPqdTf0kA7rXIQdqdzVsZc61CY2T5rm8OedENG/FpxNyNzjBFULCRq7WN0ZGi0XetmVKy
rNbywrxKNg9D3goce4f+L1C3UKpSzZRBqg5kea3kLOTHWbl9IKPFYFUV0QK75WqzFkySsR085tuq
OGbbDNOYeYmSVv/yIynWHNAveWQL+yhBaveUqQ69ifUswzCRB9IslyEGO+rruKXPs+1Bazzfulme
mhk13EyRWlo49oCIV16plNsnCSzBjxL85gpR8xcJriqk2wn2HC5oLarVAfAsEr2o7xlDh78njUbg
t5fpAt7066X0+bg/ahlekHMb5jtllJH6VQa6xUuyQvAXO36cxXIB5cHDD1fCEphJGlO2mL/izSLS
tLi60rqGMlcpKxhtcGAuTqgTjr/LJuDO6XJWSgcGPXX2SEVHvgzMCH3EpjM3nq+pmbRC2x/8OWqM
881eO6suW+nGb6N3eDbRIsY0jmCNDGPpIq5xSrAk5oi3+W2meSetTBzGsjHOuwcExAXREoDHzHFc
Mcd5uD2MYdEbdm1gtI0ElPImzIJExvoJRkPNecg4rpVM+ucqigLJElh+9welmRmXiCATUqBuM0FK
gOQTD0WPeJqp2qdjPIFKukQO8OyETKaffliWz9IB4rgV7IqUW6UsiK03DObbBhfs12v+eVf8BofD
m9CBAGEOQmkhWuQKjkBA6ZY4nzTQvuo+AHrxXJXpjvd/WxePp1WuiD+c2dXaNTtd7vq1L7lvJyce
unAGc88VQBcSeUSpAnHXfKrRoJnvzxzjkJdRQ4oOEK8rcSsYgzSd0gLup5A5Fh2BTe5gcdxmtjYn
UbNka1DGc/1qMUBNd8AxXlJpMBRIz0dJtiRR3b6DCYCH0XgZ5CMCtuMr5YZs6WBXsyGPl7NxDjCZ
+GI8vTG1qmmGNywoc6A7u9VdmbIWsFv0bQc+MRDclHA+dmH7lXBMu1PuQL+VL5FovlSQzIgcl/EB
ZnUnsd17O2Fx0gpTvtVc5Ty8MSJNyHMz0HF3STJo9VI1de19kjbJFEqRFvCfipUGR5XHkNVY7nlN
0ehjzLnaHh3exAY0KK3onxXTsw2VKBd/CmahCiygxi46id2OoYbhOgT/bPewqOSZnEUr5XPWFVwP
VEx+IX5X0iYRv5kdtdx/SEi0yrLgFaflBQtLz2YdBNwBG5XV4e0HeTicK9ui/oFbvQ50imuEk1sQ
5lyl2pF0v9DTWINa9fFApiCGfmzT4azqVQIRcLpj3syRmZA3uVTfG+4DVClpL6w2J2cmBDpKBz/u
AstQtyeDMnfooLT7zewtoDxR6SElTvgGVWg20M0WYRWtZ2uL47KalBfRNLO45eScnv0v8xzLss0F
ixE624o+7CIuTRNFgQdSQ+pUwP4oQNZJ78uVi5qa0/0LlHYhFRsIzRcRaJhIlQpu7m2CahLNi4hK
xzfmxg/YuI0G1lKeVYrKDT2TC2sLISvGRf+W7suqlwexEMUdfxR+ob5eN4ROnfZsavhpfIxjFAVj
j6Yxa9FtQYO1WmkfnDLwbALF546CzBawda3RCBh4sPOwjVwFdqSAbl0d666+TepM9rUDKFgb2XAP
vn8BniZ6KX+hXUxsep/FwX+zK+Pd22kzJDvyOrZj2Hw8LVi1FqJybeZbiHYfN8n7v393uxvGS+zn
aj5lHtbh89bHFeT2It4GCeB3J6SLXysmSsCfNjN1pjapZBPZh56HjlKkxzHXBtkDeK7UH0xVEdlK
iB+vzQ23ZAT3yaCBjNKkeI0i9QFPe+nJ8hOdQbR+5qNMMBxvEoxeYm2mn1CpHAHLhWWAN/ogQA2m
b1MGYfW5AHPwICdPfojqnxFpIrnWt46AKtoOPdMRHO7tWqbbLBTzU3DVgZIs7QPg9MvCb1AFITk0
fR3Gf3pr/dvzGBjBE9lgzCRraACQGLPiRtxSxr6m5kZm817iJ1bZCUu/nULoy32IjuTcOiLKBVUJ
w73/iPYv+U1/q+7Q8Airyv9IndbfB9XalyGbqBucU6oRKQ/DPgL58Oq93cTpoWrqNTIDeR2QxbDr
CQVbS0bi+0Ek+TxfB7SXNUOns7jA12n+V7u2q2+xLQDeyKGXIdOQoP0YaPaQYvLTS+TYCYkUb43l
PertS9LkK0h1UFTwBA+HbGYogx0sX5r00mR19UOHttqDHI652JIO0hM6gZf2EBBP4bsz7i7Mu0EJ
ah08HHpY4DEsZpgaUDV5DKR+7YoTD7uTjs1pHujI54HJO9QIEESVeo7RwyYXFDWChrPdGDgvNEQx
rbi8FRoSt/W16yPZQ69kEgMjmhS5CCIC8YKZxa/X2Gr+hJMXf0JH5WBQWlN+V/rI/uw28yX+0nOJ
Ev3yWl7N6WbiaVr24TeqfrYvJ22/o97O6w/YBt6cgAj414rlcovxgLhT1EbqOs6f4OX7w5wrwgSJ
OKGIBtAzUrYfRKhLRu/mde2UqKCN56hyso81nSvUCxiLAZXJfb2Pa/Lc0saNYshpa/cT6bLOEC69
H6C8AkAbzXoMq5kaOGagD1nT3G3bm45fKJIxevn/IRP2wswm4m9R7Dyk7+qVEZXdXTItdrzwQ3QX
CPgKe0qSUYkcsRZP4fjko06Q7E7IsPQtJ8DNgvJGOSDTMb1ZuYqL85sgfhzf8uOJMGqkR76Xcnx6
Mu57UmYGQdhZnajVfCbl9Ytx5Fxj9r/xC1f6TJLj9A/Yt4/HQCXDXXhkGtyfIR0tUrt3QbAyUO2W
o/zYU0cdCZG4XK8RpyFYV4E1EbEKyBW/3kYkkTNnXqaSqw0IyFySKOtWHV4sm/Tzz9wW4zF+C5bU
W51HJiBAYUND9/mXkrfLnGqcidGMysLqYljNrCj1i2R0sJCVDn62jo3U78OV2aujx2rBJYS1QVGC
B3q/2U9sMv3M5IRybO5/VRwXo578eckrIt9iW1HGkABmnupLD5b+4ZL6X7MXGwxjRw+ICjlikMhN
HEtxnGdC3/trYdqXI/hr+uWiTiL3g/vXc+ONUz6jh+F0Yds1SurAOVs0pTAslSNjeGI2a4oGLgXD
AYCkCTOeAQSROWTI9ylK7MwHfvlp5aEoM7rv2oWlf8E9LLZpeirrxmOf56zcq2nVBPagwV30vI1w
Vfx4nQ8Lff/J8MnpQKOpnmuEGL4tkZhXf4C0DyiBplTEaxxL60QokLjQvYBJRNoIbkrJGKVj7+In
JBpVl2KkpwvJR/fzQoZTzVfUYWom+zJP20AR9ZIgRIteHvxujVY38wObsGUOurT2AdHfJ+FAJeAM
01iL2NQi0SLeTqPBJrpxfA+fm5TfOtvQ6eglaz/BHciLudZuB+Q/fRHXWUUDk3hG1RWJakNRKnLV
GVICbBf7QChUkWLr7R99SsteD4dBm++1eRFSfNbHxs5xMi8nTQRs0bDPWmqpb8+EyLO+ZfuEh+OT
ZNwCGbyczZMnPIg9XbbWQZ+7SaQl/BZIbhioX52GI6ltIt7UzSxHtdrLkndJJldr6dT46MhsRo5l
o9EXnZl6/WL778K+4xD45xs5hePfUKO6ex83PcTeF9fraR7Qo0NSe9a7pJq+gTDWjFHvvBrj+UDq
d6NL7T2vgV0cDQJEfWNj9Pw/LG5B+K7kntsCDh+KpulFiTazmIIF2OFfvj51BglUN8GYd7YQfive
tJK08/pgaJ0pOEKugzPAJV0/zc1QVWicPDY1d/e5/eMBsJ+10TZCKVDwnzpBlLYqSwL1Vv8J4dap
bhYDsAVL5E0gKGV9cjtN9aCwhc1OriTUpIFTwa9KQoXX6Ws2h0hkWYDDsQ1kJueQzbLmyYFyI417
1/IPz/N8emneLq+r/U6L1iAjhLh+nCbzOYmUkq5J0bs+6Ch2vY0Ep+DXDWEk/vHc5g3EovPAxF0F
Ce0wZ68gLvx0BKt5HgV0X4c6EF+ppvIZFaPPTjRBrgIn5k/tAgx56KkWwEG9JwyHcWf2iSopxTmd
8eTU8TYk5VxNdBqCkLCG7PldLjvqLFdVnpyHAbZQaUiFC9ocjubJedZtQTQXN/VVDDDtmzyNDnOE
57xYIl4NlMZYl/qbrThNQawiu21ZbWQyf9404ggBLH7YlA8Anes40KBKypz3H+rgz8YEalf0V7vh
NIWWvdEUro1dAQvaXTWSJafovn0lkbeIrr3UixoUAg6c0UFLZ+LPs2cg90qlJyNs/eBeKV3AFTJr
ccBrh8cDnmSfIY26/3RV+dAle2pEqsLlLAqc8ahcWE56U9upzBv1jRAuUPKEb6JghmBR6/U1d6/8
cay+yhCxZs1xFr8qCVVX++r9Voi2r3ywVdHaU1+0K/veeHnWTE+jq0U+RNKz0stQq6t4OUghkkbm
7yU6rU7RrQdIm71HzOiIXPgEcgRD0NcwKi7Lt4TYy9hjse/M+MHKgk8O5ArE1LOhKn4fpAcZBHx4
+qaRIJb4IxZRMTvfaW8Gkj9Q45l5t7Pzuwf0zBItLa0hNnPo7s+JDIJg33cn1RZfCu1rKVb2nhe1
vO/6Gu8Fo5vLNrmXB1PEdEK4w97WNpXTK9sn8slEkhJtc3PJogwJBIowyX+dYJ571kcJ5xhD0rie
VaZqagZtmpyI7/kRwcm6YN4uPAQbAUJVdSFDeChs94zUKoD9kbxN3dW5aOhnVlz7iMkAU0SDosrX
GiFLVpqDL7dMdBtdVSxwg37EqscFe0Ys61B9RtrRoQyYqkZZnVymmM0jdVzMlGWc/sXU0kjOeXfg
2YL9iX3HXEJ474I94v2yd54opNiPKqB3iyvQE3eMk1YnTOCxYAUuBkamVv3+gTuZLRBydLNW6Ti7
Dt/gf8mrAiu3VT0zzDm4nOOZ0HUCdiyL5A6QF2UFD6xioPv2pW6GJZmJpnPGB3aq/wr2EjGy7dis
Q0odTyaputxJX9qTPBqwQF76JzkVE5b6Jvu49kalEJv1W4DIMiDBvT/bKJXp6kqH/3dH7KP1BUZD
kBFpI8vTGw42cESYEeEggBpd+kDyA74u2ytG23iSUNHFfSyc7Mhtaqip4gMJAa13eQ/dfqPHVxBx
P8uvsF1uPtBTwNn6Vhq/BouDea1VlHvRbx75XIZ3k2sFv7gcajnAcd0tX5QADAB13CISuNi19vMr
+sx2liIMrcuEQnhvqkxel1Rg0XwJVRf62KvxMH03Qd+CDazChRc7FwsFWQL88NMX/uKl4DGLaxUL
j6ME3afX7GJAniZg5c9lDjzsMAgLOsCQCUd3AbXosS3XJavqpL8xoKSveJzeW+mlPctU/RAQ0+J2
73z1bUDsBF4LaXf3NHESMfvo31xJFP0tO8zAeEFXgBsSmpl/gMIWL6PkJt6r2PT2zkr7jDAQHxAD
WCxUps7o1oLbOAD6sGg6qkSHDNBj81LAtZQxJDp2CfVMLQhVDHVEiOWS1hRg1kGKFdGneK8nZN6x
p9T3v1nrjHwPqeQWlapMgRwivCia2XqjPC0G+9ZoycUY+nQ1T65ll8WLOWvU7y/uQH9EbPSu+qPR
IGW7FTTKXpmW6F2lD/G+Gqpq1+tPhqUL3uZd3opKuRxFkb5YEzgys5JjuzXPzWsiWyqhk2qR8Kvm
5M9UH8mpND2m1v8xL7s46a79iD4y+AgtA9pLCfoq7n5NUAVrQwMUu68KMp612EoZMKXnHoeoTGyR
d4QP+MtTLMJPiYlMsDB+5LPcsx+x7GFiSC913554dtgebR7yAhDSj0yVU5p8FAJOGnB4fdqv3f1G
IxmnLbFDWmhF5eRAQIPZm06sxfNJm/U7wE5UrQGfv9Kz+W3O89X+iCgfHjn4f/Boe2l/JEU28DM1
M1fwsj4XXoJjzeeyR+qvqr03+B7ZcTJQ31YUShwqwfw07h3xkRMMMVIWxlSxh9WPjN53kxbqeaxE
IV1Iicg9JBAX4Vtn7KGGp4xhAAVA5eKkhlAVEme6k61spb+qHuPMxPrVxWoMXEYHEFUPaauGSAgs
CHNLWDpM7SVwLKeFLoA/AEaYwhdMiljr0TNloJZsTvXuaQjftqpny+j1LxA5A/0+GRn5EeOkuOLm
zKcu0hFr85M6iUqwyT8tpWlzVzhK2e+q1hEeTq3GjOrAEETyULYVmGZjNh5Qi16eIPG8vJ8Q306J
glW598dX+aZVjoPKayiu8B6TfVs+DL6LTmzGfxcYaaMD1RS+Kj95RFmnB67T5aZY6Q/BgihPM6IJ
rL1Jej1dNn+n5KGC4DilX26s0u5XDHc7s2CiT5vTWEgAa+5W0MTCDxGdfwoVlv1TuK8Q0EpojSKK
2M9leEpLWtw+3W7HB/5gX6KUPuyQZN+S/AV7U51sFOHb8Q3+39CaQg4VSL1gh9+AVfTAb1il6FFx
LpJsn+VrPKAJDRuMWbdhlw/jNbEVx9oyZCyM4+dv66xDyTSWY9WmzXE9DbnuZhrkDS8LoJ/uSGmV
W5Y3Lw/aAGuSHomdindu0exG15A3jpqwmpzrVqThLcOyK18lFDNqABPfNUNtK0/vl8yilLKWzO+D
8o42Pn5dFmOnPHeKIGwOQhRDXbuWI1JmpudLmo+NiTc9LdzEO/CpSlY9FHwrRq3eQJ4XdcAjtZQR
ran29cC/YogNCGtxSjx0OrRVzsqZyWy7o7gtevwWpo+2tZuXf7Z5lEX5Y6PzBeaja+7oI7uAEH1A
rMLukZac3d31lPKcsLKtd94oHzoqv+7GTnzWlDbOwV7Jxa2hddXqTFrlVRi6rlRdFrHhjKJUutU0
zoWjIXfISxEIzx3wtKk39G2tvw/Cb1Cz0A7ND99hCUNOC8nkd/tQ1M+XFZXKB8rVTtPJG/K+iP5H
LxIcxuSWtmpAzuFchzbpqEmQ5WE66/n9uN9HRnxFgN/gWXOZrCc+XCEevtgF3g9nQb8XGeop/mG5
Nc7JOOq8ebfS00UKkXDvwpgLd09Ncd5wGl4PFG/V9V85rtdfZuRIu4dyDf4W+6lidhNY6INnHhFV
xn9JSzpCPwnXLqMVAQyIVARK/3MZ6MTmL2BAxrrASo4RU+1IqCILnjTC6NS8hCMMRbLYIRGCP331
js3W4xjO28vXuB7BpwYZmcMYCkKnurWDV5rOai1RD0h+8EsX/6gn3ptgGcdXUj65beDjqCFdzYzx
Nt1DfgltQK8hwGcjPgbZBPJUk22zvVqv+j5sCcJdu5NmXjoaVw2B3baopfZFjPllgc+XPSum9WpY
doS6hOOIHzYOHev+FHU23n1itb2tUutoe/3Pv35JqYGqI73+I0D8ylLPSQD1Wn619hjlsV2acYaQ
4E2PIwEbCYDy/WayxCwrZP5F3W+xJ/NZbioqpjE1luhCz4azvXqdtZpfFA5bbSjN9sdD8BYlH6hK
GWemSiF1nmlib5XptFp5TTmJ/LwNOKkVwn5vmWP6D5//ImGN84Ro3kDqK5si1mfEdg2aQUtsR+wp
4AFgc612dTCU68T8nC0kcHcMMlZKfiATivxNbxHpZ9glU1/cVKD6XnhsPv5FyqgKlkRMHQNdkc6m
toHMjgwtVbBDzLvkISpTgV3IU0rBY6GAnjZHjuWMW8EhW6sHhDKa3X346fHBn045T+mW0t/L02q4
3WP/Bxp7JxGcNQyzy4CRLoAll6MJwNPwOQlv34u5iV5RtBqHEJzYxO3vMw6BeoX09gMzKLb6gNJ3
2Oi8GDXtQ6QtHB6pUOPM2AKtDl56v70jguLXNknhht+dsfj/LwTSgXACVpKpb379rAfIx9K9He6N
ooWGqdZuF8q5eJGQ4YrXAiv/2DFIg8fYffhsAQF7Hwz2HOLNcfx2XfVGHBAXHLDrcHR3G30PVq3n
Z91NJidfWQ7jnih/UuVk+WYUdgisz19D1EUBC+P/AhgkpaSwE5NA1G9b5vpO8wKkQROLHmesFKHX
iHke0NCfCY7yfMw76Dt1jVidr6eJNTwkuk0m96U7OqKOOAsCYFp41hR1/D9rxT4qSb2Z9POYGeAB
Y2imjxGjuf3Vaw0GaBefPy2RA0liuegW1HyKluvTMGVBUVNb1zo82q5Xyyb1jzFbVFM8g2g0VeAk
TU31cSeumuBg1rZO0zfB8e7BW5ZkkW+nylAcExPvpJVZ2CYvQgsjYy8r74w1rWsyxHqnTcopvtPN
4jwNkX+u0ldXNqydewukd7lEUF4eIZfMHJhbA4DzYxzYIgCzdd7Ywe2pl8nePo1tVpXVPER6rEml
rNirPFmSt1fzYeEtci+IdMG/jUB9ruC8bHmKQs+9j+tv5M7SgCuB/vdkSHbM290p3xYxbRUkkxZz
96MQoy+FfucHVOgFsAZEvyfYw3hvyneIjBNOeM/yODPYyGIFODYgZLpa4ieUR1mBxBXorgD0A6CX
gwbZTbJ4CAhwj1lspw3dweBd1gYD4zX/j7NI9CjPkSlxeOO4ctMOH7oJENPZxI0CEsS3jsXer8Er
QPPDzcSqUve8uGoF9Kuufw0gBWW/izjinsaUeS1ZvRPmZ9MfhHNpq7wlfNTo3Y2XLn858wrj4Rlk
1UTkA3okW0s+78Du/SjCkjCF/jAXzrLTikX7cvwaM8xO29jfNQUcZedQKoWRLL75evNEL/nRRJBv
x6SxpJMRnR17hdXO0Cjos0ok7oppUJR26frQGyrPSs+cOQ33P4Gn2Kwx5dXH8VqxOPVZKXJTV0pI
jC4Htao5JymZ856meky6UuJgOU2mR1f14BLoWYD8OHKQQsesztboZKakEAB18rsBk0BGeJU7cGVP
C6/qZDy6beNsLeBxKwk4ChSiF2F4g+BZFmqecsZ6l/4mI/Fg2QaEOFrcNtwBMo1sU8Hutz9CX0LJ
FRlke0a6HICpA1Dx18D1+7UKcDflF+hXJtuK1qFaSUVAbbwJlhMzZIEhztcdls9zcv2L+VUhfzRx
4msItFR+EfYocsbU8Dto0TIRSXiJnmTIWIxJhH2AkAa5uUg0jT+p478iglpo9nwuicW5ssC5PNsb
/M16MqAJ7/TsPx2TzJ2KghT9qtMMFYivACW2mM67z7MJHOYzghee6pF5Vj4Oeu0N5mA7civeme8G
dj8kTR8R6D/VGmeN7eoMAV+1B5xfIUUH4FmGlxloql0bS6BCQSgwfGdau0LnN/71o03wmaAHEkXf
mccjtuAqXoFM+e/7nAuxyv7jg8M6rFdbouaWs/5D1+9y4sESmo/cThddhvPnhj/CYkVqdAn1FK1b
V/uJFjCHuwyeRgX6FzN6UMUNV8WyGI13QdpukV5isTP9hKNulIK4ERpp9+Q2I3/tsWDjf7W1QCKE
sy5y51AiH650aopX5VK8OOVajJk4GmmyUt4kDO9Xn2KGqS2Zr7y9avJqZP794LZQxQt57YSPRoi7
eQQkJhsrrMCeg9CDaDA3ernNfEVSapoPc8tuA3TimqxHQG1b/mpvWxVH1WXcn1sahibtEVKzkhmk
1wPXCXqKLDC286sktML2BeuBBOCZuGO9ttbrKAOykHFxyoAy50fV3i5O7URm/2t8FzfmcoTfW3C8
0anJ0Fg07KGcEg2OWtqqxbB0uied5SqyVvZMr2lYszuUU3gxQ5udwZUP7OmisRzJxHM6Im6reEX8
pUcchf3g96W6uQlkZZJW/UeJRPOc5cVkQ60UTk7Xh4wGs2hjx/hjZskVi4nOeqQvA9NWzjooswoy
OZaTd59sx37brh76up6Cl0RsGdYPAAgiBK13/ws4Qa2MhAKvHZwdhW2R7/NsZ+OHDAAlN6tv0O7z
dB5/uPFaQE0EHm4hMBhxPcZGrD/TbgOVzoucbDYHxDxi7qpNKKZsKwIA1mbwn6FGDyxc0xYJgHXg
CIIsFNcJ4MLEC/vzQMcPFwSNWaZW9pLrJaK2qhUohn0oa68cpLH82OSyzTnAN8MQ5cqEyUgfKA8l
pi2i+BoW1QDC1iFCdoqD55TTuI7dWLjcGFtXAscYnHk1H9rjE8xKczcHz9jlf1Ikb87OejMm7nyX
eWjMZSWcSh4C5a5FN2Ag/KL/bYaB0Ao8yms5CcAENBUNROWI4mobKR+T1mLPJchWt34T7I+NdtG1
FxPqKnAyKT2N8NDxVfxcrnO2CQTMt2z+067MJrLUkHhXByAmfHrvbRB0DrYSGGn4MuOfJuhpCRP+
fiXTNyvp9tYz3Es8GcTtlE5NcWgJU3pSuQyqxgJ6ckQmkEDw9spMt16Z1saIZE5zjdRC9kE4jRG1
NRrjYGCCL4/0WZe3+osVPUhLCt/4GUzAWs40hMN1im1AOy8cxYOCRGDGcZiz0PSVxedSZkiAVB5Q
MDn69sSABBv7o8FJV1uhMpJUfKRn1nTzh21ZFVcbuKJ3UYxgSLIFRH4R3i24KnYY7LO7qUj5F8Ip
nwxER6cCxianR31sZLRZnB8UsSfkPz4N2WfAjkPmXrCZniQN+ST6j6vS7/EGms3BokR7aQdY4vDS
oDtmYGaq7wRqU6dHdkDjymlRX9bv0/akq1gyxPWkj5MZsODKCSho1ySkeZdzudgEO8N5GmFSes+7
oh+botDABcUaIZCOca6rdk9Z3sipXoZxiEtyqtbQiAkjrceKeJL31eTv8IKu/DbyGIYQ14tfwVK0
wrj/u7gA1ZIU1x/21cQfz0rsAnrghMhSyAUfC3qcSz8nISaO/iq5imZKtUGfp7vMR6fB6H1cQ5UN
6fyynzbwxwznNLVfZioYiZADgrF9tuZ1P/YaMc8fOtorMktYi87Bf5ZhHs99HzQYzpMPdJu9higr
OE/tvlmFb7K3RkEd/CWFu4MMxkObiZVsmKQMaLzZ6mT1xnDB/sfho36cmEE/M2zsp2ystQ0Q29v+
yZVLeAwaR3+IV1tm2wrf4Mt3UQKdJYkCH0XMFTxw38hglmFrFOAy7L8RAAxD36/tg0zpaiYrFWdH
0RDozDPuCJrYF6WRTc7erAtDB743+YqbM07cVXpYxrWOfylo2NsczWHylBIL6yatNPWocHGJT0JX
tIE+ZZICZf4ozkHBX10Hi4z410R3AKinImPIKimsF090RYAY7auidTqGlpXOUrJXESvuXGBFb93k
tEuFKu+T6m3Di/Yk42mfTg7ck2YvpArE6eBDn/8EPXz7AWLEzpI/CgraSP8DT+Ye6gA/ZGDxTi2v
ne2ukP2HY6PRQfkxacOVT0rTcgHj7T0BpM/Fy68NTcLa3a4gTdkHtPtr2EDJDKltEzVU84OUWy60
veGREaNikxkSHOkl1QklXykt4AY+cwsleQ7vRBzrcPlZiv8kBpb/jTO1N7FmibHGb3RDJAMJg7wi
lzKRzIl9g8bevjGUChmkfCEOmYFi3Ri0lu3yPF51diZhyFdSIoeluuWe06TakdxbYOHND2/FXZRn
iRn2TAb4KXtzEi1Qj29PdwrYiBuaHprrp7Muj4Y1SbwD6/DeZUqaniHa3pOY8agmNHMfkmWmN2Ai
Kao+1cTI5JFgx8OlwAZMcswljcWxn0TaPsoNnTq1Z/E8DPVIyG14gRtFKR4pJNZ6VuuIh1bStRMn
cDL8BiGK3DAvTWRo26/yG/bR1LM4UTb0DAmulO5FfUp/hklF+MuPTPr/E4H3Cy3+I/IROIiyDgk6
dFyG+q2y1xQLAZh3MvkaeANF/odu+SPeIw0CP0Sb9Ag5x/snqGg1x5JTO49CGLuDmiTcj+zkhknc
0Y87f/DH5twjlIwaTnL9oUL6EwMmqa2m4MOrsPthU5Sq+yVOzPKm4SBTdckXFUn3w7z8OBPT3uNP
GTnVw18BYjDgXdS026/eHhYs69zWI8SQYXwt/fZAXTJrA/AU2kawjCDtQhzRVg/jjcfAkwzvdS21
9OrzUvuxbJFcjgNwy96uuESEa18P5VcM2ezwyU8lyVF6D9tuJua+bX+CxUoAc3goqmeLm8ihQsrv
pZ+RFa7bXHvuuu3I37qjoWag0XpJRSlrH/DiQnACjmcxX6LUrefJs5/v1ZPidUs+ydY077q8h0LC
CU8j6FCpAIueGPQaMid2CCDoU8KCkTxQRj/URWkYFGSGP9+jjXTIdSzkVnGIV+wWHqXVf/hKcNN6
17Tt8c97JvHXyazU26ay86zANp9oR71uBYHoe42JSMzYrslNOZjUXvZ3fybFHde85iRcw+KcVquA
dCOq7J2WuefQqkJVCbI/k2+aug0UEI6zOjJOSYHZxxW9JErbgjRCCLV4n2payn/2makyqZx+3Gb8
9wnb6xqOK0ViqLczJNEdfBl0sQuVUEbghTyWaYcTjOI7stfBzJROajrZVOYGuoC/7LAYD/XpLKZ8
oEUTkG9xmbIWJQtedHbQvRU7HnifUZi4qrOr3RMikc9/8KRGig0nQH+pXwjsQLa28g3WvzKpY0cI
IF/0uOZZr1TdXhKzT7ShXeGI2iZI7pj1Ufo9Xxg2d1nOlF9p0Bh2SP+yvekBWkNaf0wW2GVkTzV/
mpxdBCGiHSkvBtVDpokTD9LkybELAeSO1rUMOsJfmM484aT6mmnEWizaEMmpMl9o2ka3ElNM6lxs
umNnQkOU9FntAyygIFrhltA5km5UGvqBps6BgSFu4zaKu/VtqV3/WrMNGB68W1vqeVyQ1D2hW/zq
HEmjoDCi9w0BatOQ/Vu72mHPAmwHyOnLVWMwGW4e+EDnKCizRZeBh+QLeLegdVsty48+rfXtyExN
3UI8h9Cq45Bim8T45tQVxIcXBj760CcO6qfHyNS77b4AHG1Bt5vsWCv76QbaESSWIGTo1p1/jzfK
MThnnDQi+LDdPdxaiLnQor3xGePin8Hm4nPhY+Rc08if6Pv5PjD6zFobtxm5U4o6wk8GAPv5+S3F
TTmatBR0vBt9agJlvdgLmRhL/TJlVfOIutqXA6sxTG3vB+/0BTgHLrsaH///CZre+P6Z8HWyn76M
KMUerG3mN2ceIDEMlOlL+skXEspMpGV2d/Ceq9dewdG/eWfMhrh1YJ7W+XFGJ9MboP7XbWFNvUbb
/pX9wT2eSY3RDYTKwNNBesbkpgLQYb2bk6zZw7Z1ZUTQrR2up9fPmrwfBCouHCW2ND+voRW/y1GI
tq/E1cJcAMKaSs+OMbzTipWCPZx4K1uIZwyMysxQ3cmi171wg0r1sbZctSr0tI69N/BDY17I0SBw
40qfZfUaDbZFHmlnR+QrQby9PJlgAc4vah3kfSnUmPCQpIVmjzq9arG+x0xWdkYLywCAWv6qrCgD
DgL0sbRlmfCJsbVbC4KIlW3bYXjTWudHrfC+LGmvVDrumvtHv336vTdoVeN71w9Vkul8Zrg7O7h0
gKjAfNJ4esdXDH0u6pEQ493qdW08r63AKOAxyfx2z1PK/TOf+D+hQZBBRGqjPAvxfmixHmYuUFId
VjjSmIm861Bb6oqZHp9cG+3rz/uXx2mEn7RKJVSf9FzWL5B7W/dGo91w/nKlm+EHEnWyTxO6NXW4
KlyM2BZH+WlZJNJgYipwPyrh88zjESDE6xaSh6OXUHXqryC/qSkLGYIJRTZrXy5XWqVvCRxXF15D
W4ACCeERIwm2AA11Inas60hXNnZKjXhhz4zBXEtx8e7P2wmbkC6yQTLlUj8cbtmNhrvn4PE3bFBV
sY4TrmD5cYM+H6ZSL+UmgN0iKJ7/1du+Uc5TeeU9wq/Ls3KSDNH2UbgwrpTZhRx0A3OoS98HBPbA
Ewb0cOj26bCqrSrfBQ8Q/sS+8B4733Oe+RQbaonkg31p3yKZ8YukaC1HxioZucxz+MSHJDS8wD7Y
MNi9UzSVP2iTwepednDVJX6dxUqA1xvBY73IVQbk5RWrjJ7yFCMd7UMQa45p7oyY8lIGJnrTH4AV
bJPoBxhFAULovLyjK8EKKnY5EuLsjLiPbeZkxfFHz9awhs/vWcPjrukBC4aCBkGZ19rzVM5fFmh5
f+5PETslECL6+lUzTBocu7jVyuIeuPW3TM68BLWTcTXyckoepGRMezWZAnnjuhh4kfenuhu5rDwm
AWyB8vb5arad4rdqmqrU6CW7GuzYLcTtY/WLqlq8mgda1Z52TGlsar4nLWvDH2XAcZdVAJ2W454M
6kUA0rw0U/v3WzFg4qDtaNOfrnATPSxkuSC3lumwpNmS26I2gAPDdG366iTWGoYZOAuxxJQLl8IA
QMV6nlXhDSmXxLtcVbUzmdLLqRlEwvJyPlGFAIIkyho1GcGlMuDUO3a2wjutNAgwLqHMrD3+MLCy
FZxxhsGOZspAGhywWA2LQJiMT0oI+kyij7cLmQ9vQAqMe3WkvSDtXmqs5LWYnaS+mQsqQxv+37vh
VWBgHOi4pOse9upcf8+TzJ04PQJGeHbqfflr67imKXQ5PeW5+3aFwvOQXbsYko/TBRnS1hqzXvDx
MV2bhvKZ4KwH8GHuY926tseqlKMmNARU0lcQhWJt5qdqLNlLqNZS83z1jHTbt+dLhhTSpzZKhPJN
mpkiwwtN1tn1FDRkAMSbKdqW2fJZ1YEC8TzXQPL40uZHF4HQGawB8AtRkl7K9phoQFmOJYyQA1+H
ghQoIV8M3D3PJ+8kmpNLXBOn1X8dEua6Br7GPA2BtGYFS+8yjF7Q9mE8in2PsDt6ciShb0s32Eg2
XATZJ2E0XF1NfyE5mtFJitdk2OBixxrKyXTJQZbDH/5LS4Ov25GRowPZNehSsyE8USe1luLeKxy/
QaI3ejYkFjJsjenRFShU0sNIXg6wDopghAnalQzYk7NjJeCD5rrZEL/Eo1GrTzGvaRlNMlDBi0mU
n3LdEyZ/ccQW4haYxu4hMgOqMbPVpWjMW5RQruYfbUU08pUDRmayRGIO0RssbuDKtqeRNCFWr7m9
l2SjyyPyLa+ZY+QidRMMbBhmA37OYBt4FTEy4avhPXwRQBn782fzZObunU6XTWRP/Hba6WRqJPhm
Mcx18O1SFUgDSOIoZE5iXdwY52CLCrjCBQJ6JoJ70Q6DUr/Z3sXWmwX9oqsjI8IYb0AObwxBPo2Y
Ue++INP0tSo1gxe9P4kFnkXkbQ4QlTCnYq934fzS5Q9tvddCbCGo+DLUvaGvPLM5lMCQXDuiGuF5
vIJIeuZD6lpQdwR9R0rY4DJLQkDfCRIBL9sDUrOaVyzJtj2b7MImFwTJehM3L9E1gauHYcf+sq/k
hhC0vuoFgiIN84hL0F7wR10Jik2Bz7cQ/GuEFu0CvY98pKdFUYprrzJpX+bJ8f8ASUF13cUsLtuA
54EkEMl/x4nzW2uRH1VEzCLgTsT6AhaKzBQLBzEqg/LVljvl1JTPHxCqX1ZKDOUnGqGQZpgMrPuJ
AZNvkqSyK9FdwIb1ht+VN4fb7gz7evhDvwKWThll0135x6lwY+cer6phTErqc9V6/hR72tAYpHbx
FVp9Mo7G8YKBdxvfr2u8DnMyyeEDOlbBvmuHeGUfZZsghesXdHeuaTkVFzaT+aRPgSp0D5c48cZs
zsatrob5ebmT4W4uxDd6lSH+6dwbINVuiT8+SdhJghpYh6e7wvPnR+siwMf1dPh8rgk5Mm67wpz7
5RIKPnd8vAi9gyjRhF6H9sx4w4AbANmF9obCbzW6DfFMLudli40mrCsw7Gf3wG4ckXBODvPG8cdY
RXk1PdPQu8BoBjh2QlhE2SZ0SkKgYsudgCJ/DhTRkzxaf1EP9rzfyc5gMPBLlqT9+9MHWQjiVUel
cmumvNmsV2BLUMEcpbNfDuDx28D/yDP8KYVbCgrfbd/Jg9IH8JaDqnWjz/eTtVCuh4Oux9PFFt4K
2FjVD7g9apr1+fgabMYSyUlIjgi3zdSk2l5ZQCmsMqCHCYp4Wxt0XsqZCMXIq3V0uVjl1szXMyZ4
vSrNMk/jRtV8tYhcESPANm12PRMxXpfCPUZCkWYBbVPc9zXOs0FyROE98hRze/MKBc9uaDJlCsOk
tQTJUsv+YMhrQj9m9DIP6nxxhpKiPS7xRSLeF0+dkDA4qk+V25EJ8wHU7wPX+26DD4sMtKl4dLZd
U9PwTXixPcslnzcG2LDaY9n/9dFqFcX5DNNlw1R0NLMTlm3IgiecBvLNZmqNjlLJp18XMoFnGU1k
zM8M+kHPi8HlgJO8BEINs0Sh+jPraJn5f4vUCU46HdOr+Ldzo6wLrNTVJyLfytgHvZz4GEJTrm/j
tf5odoH9hsd9vRnxjjp/jsAWVpXhrOldboKmheSk0ZCx0DVC+ObFrIKDHbguC/lDbrp2LX0iLv+H
EAxESYifm2ds8y+nXHiGuP0Rpzh2hC9GsAB7/CR4oq6bNxts2S8T6vlBZQbfpeKX5NjpVyxiIuD7
Rnl3jfd7R5AKvMZ7c99Fam2kX0VCnvaCigLEqJE+0V5rdIGrfI3E+3giF5eI+XwYxKCmth2z/v6c
pEp9jVVW1aVZW1HyBp96k0hNzbxKIOJmEG/bCYrQhssnIjUMp1gKMrvj4Suj9M7Ej/sbiSClP+3L
cCTP8RG0xXa1LzFz5VdLQfVM5Ju1N0ZhyQZu26dGo06SRQT+zwMAwcBl68JJP5Ub9kmJ9pnF+niM
sM+/ITgg6pyfXNgnUg+zexSQZ2tbVnROlDrtJX5Oa/3zLBsOlbFWwQnovCRJKLQzuni5yUxWc4q6
r6BTyKyWppBS3l69q1SRBVX2l2+/SXGGL6Bx+dVuWaiNk6/Flcn6BPqoak3qICYXmozL/7o6RKvH
Jtft6YmFYk7BDv7qbGzkBSjW6uVM/tegIQMEfSkla6GWprABmlS366pFRQAom9I2sRfy2XE+Hyt8
nC2xv/mxfbNFFUBYdZ+K9qAUk94aFKUc5yMFAqX7a7D68CVAe/6oxtZwMszAPr0cr3lrgMw758QN
5zQm/WnuYvQkMFpR7rEgvK3Um1YxpIRLOSMkxajhftIx5GNUqi5NN4X6g9f52pAzbcmKG0Dyb6yw
CGB1n0b8ZLmxjYN/GE5Zob9cCtKMjC7doHgp5IPvvgtz9A2R8ApmW+1PAVK9e59ABGsRGMmgFGS0
sxh3r3VXE4qifgAtYLc7bDqYushsZeYV01qW94/GcgM6qAU5JW87OuTQXpIxMDuLm9KGaGCeHSXP
NRJlz1rZHxBOwLp9LfWhkiq0VawKdQgDhf1aCNCgkYbanFeVHb7IKD+wHu/LYH1F+Hz9Ci8Nhr0G
M78g6m4DofKnHSJFfmSa98w1jlFrvXkooFgDpTLSV2d8oiqwUjlQVlw9btN3/9u1UU6Il7V6RD2a
Q1fJjLyy/JHLhnruWEN3N47/4Qk0vs0ft/OneZpaGbULrOFVHW1BcZ+VlClRkdtTpCEnmWXs/j2N
JaijNF6jKoJl7iw6F9gYHwKfEphU+XhgxpVxmwMwmf2aZ9S9jAZL8E224un0GY5uGeSRt2uwm07G
HZaoNH8llFu7T7L8hUPlFdVx2+7ugeAgAzRwevpJ/1XcBaQ1wcuM/fpSzUVnqwUcjXdhB0ezsD88
lDUx8buXI969/CwLst6oPKdCZVbEIDgSI8FLNIAsOPrd84dciAhuJIPN4CGouhenLD+2EDCPhPVr
Ps1swbltzODvCoMpsNtjNV4T9S3HXDLwR8nmtb2wsb90V7DYcpnyaBB1hL6d4jB6MdGZZFfGeiq3
P6nG057ZamDgIbUuJ/t6vWKrfD823/Mc+4MqTQpuXZHZ6Dd7jHXYG/L5XtdSJSjx266REhOxiqKs
hugwZaqXzp6C2Kg1T3RO1D4YO5SUN0Del/1dFBC5wRC1Ni0jAUwjB9yLP/V+xrIEeJuds3XLi9nd
tVU6TTxCmnLqjK375S+MgPorCIvbwhRMyemwyBS6FMFJRSRDotQcxyGFqCC1Zc31ETiYZaRpzTQc
Q9Um97EsAsQp8PrSaOXoRADR57REnwsPCDOUcTdjM3zQCYKBagdASaqwT1XYxoiHcXi4oY7bCOSi
SZzLh7GAOc2Z9+N4uFYbyo6SoP0TSo3VCJ0q5ZNUPIHl/k/XNhRiQIRae/ek8lRLbf3zgYcUhoNz
v982V3A6MsAoDLIJt+3STRcnhK2WjyYbOdUKHVzWb5mvBsMdz235pikly6SorYwk8a9rFxR1oBkL
gxRfvCRePBCIIWFtc8xscCqoRNwfnJ4AEnmJBXzItF255in9XIrh1iGSjh/tIjS/DggAH/2m/j75
qLmnpf7A0jo0JnyMPsFhCnHHS3roM8Zv27D/TztFGI8hMBPD1HslvQQjO0wyvVd8tu7fJDPjToke
dRByzdLucADyPWxXFlktU+5ego/rsqeVgTlmVQUTo6QMpUtsuWNji5W5pb4yyc9UYjXnATHwafyC
PzWAcq2jBQs73xYRvd9mgIdwjg1XyzgDJ+xNgchputEbth3vF81+mlQxy47Wrt3/0QGrLlG4BoFO
Bo9Ybz5cyOFUPyMKotKnWS8exT8WCUI4Xqhxg2zUVQM3yyOygg2xnufGxOmAvHM1mq+4YTyUeLMc
sm/LsMKdI7AvZVb2kXDfyOm6YuXP/OYcBgTa5sdcsHf36jqwEseT82epYttjDJWzlVl+1r3w1geA
j1rS7MNJQrvWZ9+yRElyvU/+tjjhbC4pSW1o657UDDUZxfDq2j3pJ96kM5KskAB4E5tDbd0yPEk0
XlpMXK3KvnGRCs3XhPBExJOb4XdLwNlsoP/2sp0SD7Enx7JlhXDPnum5oa+FKBQbyKqKInPoAUeF
EBhYPtRo+iTqK2ghjFrPdDCysqVnEHlYu94l/gD4lF7W1J+nZ3sYiGVfg7Hq/ZGCv37bDjVZLz5r
o2hOd//zFjq6owkxcWcDo8sbIKDEd5kddh+MJCKg4VMeEwuH8BAGOX5FlL+uCezJB1etNMbjMvlc
9WoILRcK2ETdclG5IliQ+yIfrZCoy4Z+Ss7BMMxVc/A9aK7MmXcO9a4aoqcH+8mSuUeokOMrw2zA
sA4TAyBokUjLkJdrAose1wbZkuFeTGIUeoypw9umwGdTBafwqWkZRPif+vL4lVPKjQQUJRn6yfC/
aX1SJmjMtjeKNcTbkBMZCvbfbm9oHN09zxN7NJN8z7OuKc1LqrmURMUDnde48u3N1ZeGyxqtJUv+
ElCKOnotdGc2cy+m87ST0xSdA4ydNCpqvp1F/YBTdkBSjTKWRl5EBkeMyZjgBNi9YSibK1Adlj+x
V8Ij7NkOt0uWDgE6L91iY16Ba8VyjDv5mxqQJfLMXINi02xhS/FZGDEjW9uKtIY9U5R2RkNp9hod
+AFBvcxPU2HbLhSfrPAKnHTFb1B+hWsKgZSEbsia6DpvkQC9oLVvOlgmWxuPMhT0Xa0FusoywlNV
16dgPa4rLPMoZvPBrQr1LGyHog5qtIj8pKy4W5y4AU1E/n/miarpJ3BYr4B52gsU8jjpMUeAwi26
xy9e/5I/6Hc+wcikRJ1sd/AZW3KkNBjybiyrx7iDN4PX2PQXrdQqJrhT5vPQ7OJlE/fVw8Taypbm
6EVcLaCl5WN+Jz6dnP6vNhMJkIDZXA/H6Cmrwm5067noxIomrqxbmI1WtJ/hGgl5K7b9EoyPwTh7
9gnHru8qMbPhSkPKevAytAEMvLmXlUt+qo3JP2xWb3wR23g6NcE9ma6ZhXTVA6jPDcl0OQzYzbgA
g2H9vBAkkYzvwWNHKsnfg4rpe5iSXQahFyUKpR9IiaPcI2VensguExZXndHYSARRlhD9WqqQZNg6
kLjkbFt3vyT9Lbe7S6HEYDDL9QaUrXUZkc+pYKdIAUB1N32BWb4x0T0od39Pk1AykPR734w5irNL
RBdKMCWPplo8Iuk23ASCMrYLwLfHYAVLkjrk5eC/PBZkUrZX4rdGGkYfCP3ahMRx9vw27mAremj0
VOoJl1wYttI5yksgyxKGkbsJrUh0U+PI0TWHzdxNEo3SU6+WGhUFhQcYx435iErX5+YI6PHS4aFb
ZKxx5xiNkuro7QoyiHHyWCoD9Al1/2xQ6nDCJGA/hsFKerMlOFG9jFuzyfJpUfcJ4vnptPKK0sVt
YCAMW6r+lN/u73AU01t6kouG5sjhjkH8ByTmWbGx7RuOTcRY0qSzMR4u8pFgDXv5XFcL4qk4c7G9
wCrC/9+3NWBE4qEMsw46qx7l2gjs3ip2XWZ7vfGlfiuzIBEYz8SzrcaiubknA/KAyG4g4R9sXzVJ
/lyx05GlHAzBIRpgk8ye6ndV7Cj1Cp6mhsEI1ppdvXYIjDqjfrHCmtewOPRBq/akfXFvKaqxYKoi
cvwGNwrvbwXHvCOx834Te+RMB+DwVK/G0+8epizw98/BYgiB4rn1yDNER9gSyaCovukxalgLQRjm
lgeIaf0HxkJuzD4vg8M2NcIsRXRl8nFh50OMAv0INZQVV2084i/h8dncnt7SKEN2TLtW8SNTJVEB
1FpibkfCY97h2hod8NevwrJxDzPhBfFj7GadBq2vhoZ5CHXLHvhJ8M/KHVhdt7H2LNNfq2z4bcT5
lfMHV7UF+3gWnRNT/2ZK3P0dqRUvlqA+Ngeik592PC5zDG96JfQA2Y1MVFiQRcWj79rPPibsFrzA
tKhLSw7iMHHaAJqToASQs505EC9cY+T18V7VYiGLqoSR4CO6iwzd+/2OR39/w+OKid8SzYXe5uJo
ZkfaJoyZXrV3eccn2MAabW3oqpnslAzoWbOSYXXQ7DijA2NP34f/jQDwOlLi3pwnddYNINXZB6N8
goOQMH+lFfsxBohX5XXmcutNyyI6CkJa/XubGCrnx7RZBCOJ6bph6S49Rj2iZJ6x5ybRoR0eqSwC
NsggofGNizqMm827KoAqyW/vDZpYEnjdIT6hxLRWLklZhN4hrjx3Pj+f7wPRWiKhQwHyVp33y12u
v0/7RAYpHWhecudRCUKrOlCVv2XgKPV/+mZP2VhU7kWFXfsR79PuFZFEGwnW25FKWZ9O3v0mTQtW
5wckWWy4jb8/w3e7vPoWFGeg/Z45+ubzu7MAbueutLdOGKbUhGKlPnt4cYUK10T8JIYrPKe12cpn
ImxOEpsl5L7A+Jt5W77XVJHfSTVB4oFyAF8wvGe5j0/LakOMOj3zI5+9W4WcOZeEK2elhEWx4kxD
og9nzc0mGeWbCxLgLJXRaX3tY27+bj/t1MG2Fvt1sW5FA/vG9jRzd35ouZHxkeRgXMWIy2jYpXsu
iJ3RqLLn2nnLQUEGn5eTHJpCyC4rfgxYijaAGqJAvhigWihLh31HO2a9m8x0bUTc7fDi51BGuPF4
IZMnQyKfiOdvv23RwIUl9UkpvCJqUjloCmQXTPnALydWXQu4zvK7TnakY6iwaNVK7xd/t53qea1B
NthPmHMjSqfMtiUbyQ0mp39qVWUDBzThHHSQll+11uGPGAmSnGYd+k3/LK4E6FBAF5KB70Goa1iR
umqv2n2V/XDp3IAGZ/yUq1toEHthBumZrKHJ0RWwZebPvRaAsuTWRx2ftEq2w2XGyBWAew0zjflj
OJoHeeMcLOXYPxb0KwKpfS3sYefmWa1dJNO0hYiPU8aABQgvPlWu6VyDGCuDoELQKiZC0hhkCrlk
LBWDxnww5aOXSqdxn4M0xuX7kz/ZExJ6+hB5gzSRwZAb/4gLC2my072euCHqjfDUsjjUzag9Wuxo
HqQTBcNVQ9MGEjTc7K/pGSUMkoDzSngRDY7FOXt3wvDOST7i5tUFVif3S+ym6h4m1kYc6qiQG6My
PdTtm/m8Vjx2o6zO3kj6eNf6qiX29XmaGImm6HlCW3XPYQjttZZDMyCkkd6qkZ3vTa+86Ky8hHm8
wXJQNmH3hcEGRZ79hlGtl4Ke2aevRIzbO4xVCsDx80smWAEvSVV1yEGfE3wWyNYqlUPw8fcw+oVC
d+fgajmsS1x69c/oVn0j/Xa3/gth9N8McTrmD7eGhgFI5UpNC/VU0GXQLTaKKMPlRKen0cd3d17o
86lQLjhlgvcyAH8TDFPYvdtaIKOv4SzYhbTbgvHu1is9J1USEviuQpl4fGiIg9FBmmQYj/aZa+3J
/zl9CRLt+8XMLsQ9IP9ROPXlRx2S0RgDIsGRtrIUmZhld3E75ZfLBGNeCLGYBUai6o3EYDRMpbvQ
Bt1ktKkm3CNN02eihM5m4CW3tzmQoyLWPKRVWBXe6EUGv5c7JO7gAC6897elN1o1whBLJdERiMkU
tcLZR7RauOaZcCHUtvqRupHHgDkFvAkdc7RNR4SrqRZhWsCjLa5tFIdVD6OaFzdmU0i5UfrohM8h
shY2pRbhcvU1dSFrxusGPzTpXUR9fqSfrub2FpCprGIOLHwjsKh4Kw1m4jMVNQC/ppsUalHzVlH3
fGT/rqAzFlMjaSSrGIeC6pRzzNzCc8rYcJVAROWVYRsB102qj8A+9b1U0W6cggscpRO4aELtTfOo
/2+atEMYbJnrfBjIuGpop0JAhXqMO4Z93Jj720P5kJSbVXX8ZxwV/HVk5Uy4cafA1K35bvXK8lUS
vDl2Zta4UPUsKJJ8tFL5B2akJ5VpBvhJQp60LxyjsfJpZRg2sXWjhOIqGhzASvxQjQmkkjWCpdCt
3Yd2J80xlP//LFLIdXcBHqFumTIb1mPdKcMHhSrPIo6oNKSn+fm6YD5KW4ECc0jxWTPMz7Aq5lrG
EKhyT+wEPX7tw1KOP93Bh2t4Mu+Ud9e+RA8/pkNPGTAwL6MlFstCjTfMZdDrF855LCRvIX/JOrLd
ROA9qdrcJOFtv0lUJNwkf+SqnQv6bGf9Z89FHHX0uL9i6SBQj8mW2H6mYpg0ElDRkc3iA44qtxEN
ulZDHvanvch6UIjEZ+TccBYOIRBBAKExoiE2G42Mf/sOamvTFMcfywbcvnAoC76vocMYaprGrtyy
RQQZ0qDEcNhnYR2GHw63Abu3/URgFM2k61zwfKqSc+dJG934EGTGKHdGjr6qd3wekG9Y4CFqaBMS
ilSYKLrSOKWu6Ll1R2SXBdb9fNwy+I3a4KtYEk63y1GkEtQrmVUp9UZNZRS1EkHLw038PhqVbxIb
9cKfQhF+r6mkLtjTk1ScGJUX+a367b6jI3RVzUfU/JycOEEPX9KkTzPnpmiBaSNcauhLGbPGvU6c
5R3voH9L5XDkgBkLM7kO4XIvUwV9JfgaYay/BgUXGIoeADyiPGKcy2lOmoBChJqp4v1ONnREoldt
6qohNIhntvp6TqEZaNtFNkAJC989JP0/nRvmf42ZDwGhk1gQA3U89V1jDKiU8YMFVupi7y/xYegq
OD48+b9JsuljPq8NPV6i7nT7ozkDd/Mk7/zBUn1qbLUwrwFpHl5/Zd/FRmYDGlcVSlYWfzX2/Jas
eNTM9K2N2LYxWB751wILfOsmoAVBDCnmfNVRjgIBmKCurWIWY69JB/Sdm5dkCG9BtYX8KzsES620
kTOQvGIr6DQt3KbkEa9dW/vqRisBjfQRcCNSqO7ezdIq54s9q3gPdznThNe8kDMgDVr1iw0OHcuM
T3fCDPO4UCKY5rxtU1vhRg2oDuzy/CeVdFni1A+q5lBmpK4rHS4r1e5nr6IZctSmnHPVUW8pPudo
aQ2T6H4zfIyvXGdgFLNVKE0n/JpaiHc7yAmLb8AM7AafoBiUhQpibFI99LcSa89G3BPqWmtGfjf0
9SwPQ/TA/EXa/Ax3inbUpsidE98TIdTa0sIszuwIX+MYWsyA2Bg9BIHHxfcu2hQNS9VUUHwS9kzz
GlC4prm3TMcl0y7QXMhdi9CYLIX6vaUM0sVRe3ErAwFJmrPpJeVxQT43my2PyRIRMC+ucR//s8I6
T8Quv6YUuXdL/h11nsqvnNVWwTdzESDzA5Z9C0kGTbCUOgGEB2tl7NJReW0+umAnWKHZwq6/T+xn
c2WcovTMiwKnI1ikjkdxRIpbzGWXcY6ufv3hX/Ruk1iSrEOb87XEH/UBMrpRetBsrk3oYjP2oGcL
pFwG3TBtpDl+Y+wGlXF6kcZhAn5wuFV6LKYQto1K+tbhJnMdzCervjyDMeszvmNGiycyWiTECrUz
7rttSzcFt2rBmpCm0+TOVc1FjGD5jcHQx0b/VzO5Uzroy3pQJMpz58ivQ24hmBEE3wfQZFZHf6RA
H6SQ+LGPX0hEPaH3ecL+ar8cRQOpTrS7IVO4O/rm+/Y68QSZVfFaYNoq+XqPI1oGsTzaQj9Sk4C1
t4qNGcHhwK25KfyMBcvSZ8D3sCgGVnWbABdw42IYJFPKLtLctKSUaeoWYNllEjUVaOvNSAIVdMZO
7rpfFZ/2lHL0q9sJODM/NdY7XNBfFuax075e0VK2sw6aLT8WvLn0CnDuUOu1jqNv1WsPl7dcN0kc
yXWycqmjc1H6ijXZ6QkZ59egCOakI4ksb1lFZFVzewEZUKU6DTf/pi6HisjwRbn/XBb+M3+wfPzy
a3eaLdhNxJu/ZnHUlZGbw/30tRQOyjMll/ORmq2vONhWZ2NtA54xGYLuVBvcKln4eexPd9TJp7eC
PceRzz21CfVZdE+V9Lb87O6o6NyCxM+GVj0889DlEQzQdKZAzGxZTg9BD1RtOGfxHsz0MfNI0DyD
YOl471VK/9HELUJLvrVkV43CTE/lp/hIPCQYdGlCxrOw2wZxcBDoYzPHujBvMzJ5HQe14kj9wnYo
fdc0MUg5FOEKnkEHTEGH9JGtuvw4xCxTj224BEgzZ5eZ+/LLR6AbK2y8LHpS2mOdgWoOdjXKJr1J
R1kpRfTPc0h79RYI6Rci+tMoEc2w45lZZj7fhhluAu8jofAWpHE6p5d4i+HGU53AaM+I7i/9vKDY
+cGECbSq7sYqSCieE1MkBBnoF7AmunzMxYEvBIx4Lj+//OfLwGWYwEHVr1f69iD/eeDwrUEF5bnN
m9OADobXuztOAv3oENhG8nxYHxZQrt5Erq/uRZFeBGF1ErdqZ1zjOyIgo9O04n8dffZDe5okMBVr
2wXLT1/UuIiPsqzMFTTWgdYgE+cRLEGFk/3bW9liY3ijuN9SSM2sunNqVQ5XN7GWgJnQnPu2t7ut
oiw+FpuHXMhIpZpXYNNdqKNmaj3B2t9P5z5sotDyvMhuzhDLtBsaDSjTKFoqbwo13k/N7MEY2fOB
rCl8TISAun1uVWdabKpds62Srsq8ge0tDBF96BfBhzbHnq1BYnZcS9VWj9jj9AsRuaAYbo2Of/y5
84N2t1rAtuIlK02/YUiPPr4UJqT/2iMa8+LmMi0BnTNxWHwnm9nalXTJx3yYjrkCgbWddHzw7Fgh
Ycv3Kv2zHYatt59lK4LSizEn9Z5PHk8IjhO5zvFoBeHpkeMGE0rAQZ3tF5d0+vB9TvzgjsROA3V3
dgZsXqYnado+0sv4rRQt0VWsv97ObfoFCjMDudl2b2d6ggnyqCH912H+UXQWlvGTDg0k4qQIkl0g
/46LGKJ+AlyJFm0CipTncJkTbs46kD/79eAtcwoTv/C/HNxWvDzRUgR9lX6on6px1dEssF3dkWUI
rfkOU/RcJeduddB80UCUt0gCA2wXTA5Be9d2m0zyrToZLabK18J68+G89aA20Ad2TYG+wQ+7GKfh
p/Cw9/QGdJHHMjozJFI+gGZWtjgZb1NM6QOdNhewHOlNP5/XnBxIantesyTk7hfnIlPy+odbePaq
l0NeJUQOJaQj94dJoZEDG/ZozJ3KVRf58fbsQ3D0yInCdJNV8elfHZuakB0aU66dIdsf675AdkMa
jpHJMNJXHoLHsamtSYy2nsLFfQ3LHhIB412ySQt7x+WkbjFgHKXHlU9kZETtgdlpngU9uQqHDoy0
LOZ4YU31lHhYHJ4EbLIgn24jIXfKeVzPEBduhMBNeKo865U3Ec1H0gIlF9FuWOjoeh/yxjnSyro2
Y/J7zYgNNXfRioDU7MX85xVwH19sxs7v0wuWWUuTktMNEjW6k/IXLFjXDlvzS5lOt6NZlwtQzInD
9oquqJWQG+nGaZP3WR/uk+pgGpIAuFRRHm3skQAt/06ID/H7TjIwOHc4agAqmUMghrGEtq1eK8TP
s1YRHN54mtccGy5Z2fXF74DMZC5ZkJgIPTsKCE7H7P8PQrV83gKKiTe3JIg+EWD0G55r5mBtNvDo
v+pDaW2zRWAbwMqrAM2zcQ5aWHBafexBxTB45l88vDaszuydzr1YnAS4SLJLeN1dA6Gcry+AaUNz
s9e0baxjKiCOLML2aouUC2OKi2PFdNPJWY5z20s7oHuEETCWzpiYRDF0qW1++94EjIiu7VKeTN+W
/NhajXOUYhbM9IXTswKygWx+6FRWf5t93NZEvirOHa4+jukTkPMHDxmERZ1nTuI8z4FT9MQ7o+Rr
B+eWTXGL48B0CdPptOv9G++PsMKt6UpbbOooXuyc7xz2tKeRyyDRb6w7hfFVzbMU8wOply412DBm
BwPpUJA6NAvndacskyadFBXp8fTOeeI5Urf68OtlZBakJ9L0xsUdCT3qXy0qKruy9owzZU+lmwrT
Tuv2lQIAdNlcJ7n20TtiIn+302kbZUoC7i2wC7JOooyv+vyOVEe74kmAbvFMjdyvWmdlRNPP/sbf
7gPzjYfmxxsoo8dPbZefdrYV3Uj+0iyf/hyAFVEUdD1opStN5uQdZrh1NUetC2HfBUJFyndNDUAp
6xU5/yrjTgKIELjT98hM3q2ib51bihhXS9Y9NfVZ44lJ9FAdvuC2NVYZYQRmgo83MiqirLzoJdL/
Gq+oobNibHugrFudsYrDiv/PbyJVTlgAbnkuKp6TaB+PYzirbIY/1Pu+AEK+bqnbeLb9VPdWHGAW
xkczB/T5qCMd4lulwrYAsjdTwSKOkSi4du9bcwXvYsXthEjvLSBmyhHMcgYdTj5TIlQ3T2hJERAO
bWDnfKaR1PKC4GCCGZw8gU4UsCWLTDB/pjvZwJfOuV9xoaH3aKIjzhsZFZ5skkQQSyLXlIdp6x7f
SSYHe3fXBZRkcavNG5xaYAnFot+KRwHF59WcbTrvNbIOxlVqTIqwvlhOMfKt8P5MRy+Dv27zu49v
2yGslCpAm0rcu0vhRcWAtxDoiUKCos0nHrli5m3spyU54GwOAE2duPEwHhC1Lxiera9OP/IaCZVD
AjPLBgrVhII9m/kY6m3ugzfBIt6pErg2z93zBwouNXvzUaS3LhuuaZ/r3jqvDMB7irhCNIPlzrpw
IbZpOnUP3dyHH7AKMXhUMDPvTcf10S0lZRJMug1Wt0GyGY5HjWlJpyY7x80n1/JdJHXl0MuKPk57
I1ZDofy4jPFkIxoNVyXucsn79yCibHg3/38n5ZmRrKccLdgdcYa/75FxQgE+VKut8HVPVI5W/lhL
kaa8TdGPmv5qd5HJWlAD8crJI0zcN+GbuBxTXRxKGyOu0oOPyWy9/qIq8ndZSAtdFxsT+fKIKdDJ
f5M7fcfGfPwk51pRcvWopPhF5pG5Guq68TF5pOGU3Qc4y0h/GCkW+VVdSlWy8p2Pi83I9NtXaDTa
DzEAvPWrUS6aOD+NrGlB9qPpwzYtjuFh4LvBJjKNZqKH6vtMe2OkGSCdihrlRrUFDb3GKHP0+Osi
psJ6jWCCUkUGPri4guqVE3DkYHEcE6L9UqVe7get9dRdV8MDv3NfoBOiWvrS8UkxSzwFo6rlNx4I
R+JqQ8zvkP2KL/N+y3pRlSUaA33ukqTEI71l9pF6tIgS/x5F/AGzBx41Yfe9lniTDmvLauEnb3HI
fX5nwsSQteaz4XPv1y3zz4wH1vVO0k2QPoDDV6UCai7w83e56YUGhdIrFl+9ou1bVaO6EiNzYKP+
+00rMUe2/dfFGGxX7cujgFVgk3zn9DXgNS9FD5Cq+H1o5N2GUgJXeZmPFqemlwgBh1gRXWrjzSEu
g9yHZh3EKI0eM3AioOhNzwkwSlX8o7YN9j5ccoWN6ARqiYskhWdBFqGguZpE1ukE7/HSTi4k8FSj
aRup9av0R1PTx3EBukAW1GWbo28E8OUZ/OSLBBglu++6GxrVIAlaKw3n/tH3Y57qATi07DbgLjIv
3fjg6as6hMTd+GiSBVYkfqa8l8BkykmDCDch4tRv34QtxrhY2o6WNQqxQnnqgxMbXAhbj8q5IKhL
vB+fYexSO9as7ia42ldPcS2e3a8eqZkcu6aogB5KM9eg3eMSjog0Rmbm5pKvSQkoMdVaB7xZafF7
EBQAwSjuq0yBapcuOtP+9zwnKx1mSpaIY8zC0OFX5sGkiWmP7bdycB7l3zRizfLJKsuVo1HJfd0L
kGKKCI3zsrsVA1AOR3iepzd4xB6+HM4uEW7sCizSmQ/hEqtpx32RXNSDOtfMZYUu6WRxAAGGPYFC
xfzhHU7MJvhPxq9MzxMVzvhbp5vSMT6sZyEJST1Ae3kPEMHduhK3akp4ry9cCJciBQHQhLKRaqk9
vxSMBzntpq3MoKyMWCbv+KvcdBARFBRXtKZE8eStITrt5HX+ofetSFBjjfvbqTz/5F60gdEffHFa
QrS/XG+xenDIZku01hafiYueFezyBWzMtX2F+iAep1abaautSklTgFe2XJO6rcryCSExgv78XhSj
klHaNFZrrSS6aNNlhFSk6zcSM5nEiugcFYqnV+8jaE+/UatFhquA4jp8ekaxInbchvPxhA3jVbx+
aQhUYXhDw18Zin0qnz5Lf41v+WO9HBdsQe0+SrurG6C70/7Yxr6eHVAjaPODg5nEwMQD0KDkIlnv
wFEWlxY4mUcIa83Cu8iFlJihwWth838U1BEjAD2yA+fR/pupqg4QobDIPIIU9U5xnzRk/aG+sbtB
viFvmkIWqfIAEZOvLHQ5MyyKOXzczJKMEw/epSd2fASdcmIlHOrtwXj8KiafRlevdYI5PosVNP4K
8cMgmLBSzKU89GI9h0C84/qsMziUZolKA6gmCThDOqpWuTtF9TMphdd3EpWA2nwbXZYWWmV7keMI
MC1ckyeTqT0XJjjsC956xWvRZK9/GN9VAXUSXmhIHUkuDpaYLx9eaaq3kprMY8RT/+2iH1RLKvJj
O1+gjCeSV2Z6jlcwnSkpHrWcHpwu4WW7nR0aFWtlo3PLGOp4Uw97TGOQLnPaLXzemCKjxEvXNRic
c4L/V+a2igIiMaW7px4mRgZHkgHxU3crf2sFaJ3PxgprDo1C6kV5vnMdlSHl7j/y1+soW8cSy8xg
nhFLnNM18LvBX2XzwY9i1mh05onxyC3rrulOMbOBicpAjyxT+KUubGNWNIqnC/JDtx4PMsLiLIxT
ha0GpIPe5+wjp2xhDBzxlZwOBopf/1jjMhVpeYKah8kYxEVt53xMhZa/5gwcixQv/BfJEFEDIKk7
MErKQxrkuBeSa1r2McJyzJlUmiYMfpzTmtYs2k3OF2xlZwpGMofvin75B61zH2vRl1qSsrcsJcAd
uZzgDm8jKBC8ZcxlHFs8XM8CWjrd2NN5IWg6z2mfYfCZ1iadJfWvYfCrxodO0fLgGPPtpPfXGCQ3
DxnBp7xZ+3u9wBGE+pfLzSEUo4IgvCHzsfWICR1jgVh0pLH3OXnI0j4qHGxJbMqhw50ROnkQHnLx
hlDAfB6MgETzYBGmlObi9PxUnQzs/AvvS0wAj5OWG00P10LbK7rTsPbdwxEwoirpdX8rTOeKJwN9
QRdH2SCSMGgh19Da+E6QMTwNVoLWcvbLVGtsMQcDArztYYCCrHzkNdD7B1BeAKvsJLW4WvsbB8v0
dcQYkdDmn1fdnnmDsrdMygEkYSx5l9dtu3cmXYqXsjoP+ff41EWs+imYxaZh5Ekg2sUMfcseEhNd
JWfiNJTO6PZkxh5AuQ3plEpCXfQ2ltupoJxOku9/qAwrp4LJZANrAaLOHU2w97ppH9EQ3XzW811M
ejjJich6uGLB5sbWf0tfd71w3aOAAG9RtO8lE/1GRnScahknEhr9zzjnesDx9mtiDTljKQouZl+m
npf9z+wTtun5uNbB7Qpsg0Zm1+MUY6WmlChJLHiD/XoUY3TVwtmr7b6kXOPEPXmo7zq61mQlZvUE
cGxX3oBb5uDTbUExBcaf7xwnAPM4Y26aThIKNbZWlMKt1+uidKfVFtJnFgQOAeMt4kLazcHQLj00
0CKnd5b+2uy5AlQB/ipCDTTH9Xfql77ZVR73d/UZ1vXl1p7qGf+P9tFYOWfHAqJXeLQItyKacwTN
k/xkP5fmX9aNWViVWfDSZuwzecEOIGwxLT+cZ+YvOVGXeK3ggUeEmQiydr1U6rzWrCqIiCr4lKQ9
QW0GKibq7KgFfAeG6t18jj8T2tFj1NeLnEtcOexQ+N3T9Rc+5mAKZ2I8gROwRMUIIRuPPBqQgy0t
MmvRJmOb1vEdYbGft6csVNiHdCrhAoLnLMZSm0LMF46odmO+KAj8ay+ZnwgaQEVAsC+RMS+RlJq/
b+dE3VQokDbicFPCLUMPbWsMcwaiVo/mSWAQJHm1ZCKaoh0FKB0WISPezJyVzJ8eiZlqkVL2rG6c
Y2o4TuMzC1asi45ziSUwA+fYJZT1WtiluGCObcmtl3txzXe+ctPRK5k6dXjo6q2ol0HnaV8B3whl
ZkWWil3Co9X1XytmMgmW7C3vfzgE3xey48BjmvqD+utDN/f9dx2WXnd55RMFcS+b5QfZQ3ssLS96
uUN3ibFYK8/FmF4SST4bqOIa7fhdH4u/9gey0Wmx3KDLES+2FS4BlemsVtCU6NI4ggTIiUDABkZQ
1pydILR7jpOnwxANJNLPNOjsmrwFUTrL6tNfpOwiEOivIYy5NpOZNWnXAtHzOSeEaD0Nm/FaYKzQ
kO9MxX47ws6eZG8qKaX/stXsx6P76SGwF5TBoNQeqdNFEqUOGHVS+9QwDedBoBSZw/0vtE9tzHpq
Y7eAsfD+dkPVfU4ZnAlaES4kTQZtA1QIpTSBEeVSkULwsAaLltB81zzzjtRSuykJmPA3lPxNTYfB
CDpSZxSoVy/MaNk0upoFknc78ZIWZfRLRGTJ2NYkNznuUFrXEepMru/OylnNEXz0Gc3JcZcRn4YO
JFrKHN0dpxH+/cyE8WR8SFbmfalwz3rcNNwm4kwokheLPjsX2ZbwczZyjtu8m1o6qhaWTwQVehhd
RiefHg/kTsoGQjkUJa1XPqyX6j+5XK8rbV/yc82pWCLiQOP1y5c5UNiXasJ2sDXhW0I9N4X9FIhi
xzL2MTwgRqyC9w8KWtplS0g4p3zmtve4i3f2RTVGVle1Ac0xu7rRT+4fzLKcXvyQ1C5g0mtNW1VR
F/UufgIkI+u/WD2GKK50Db2KFO+uKTXCwFtaiQAvoDUWnTlpiXCHGMBbMik9qWJHg3+fRPlzPjeB
bJtxwipm8bT3iA8K7xnsKpwCFFIJOAIbo83m4L/V7+MGjw5xU6bk8bDfC6aWqsCM5hKCzLRbepgv
IFUTYiahLMqp7UdsT/BQs+ExVDzjlUL2KZWAxZpm2wyKuMf4KaYUMwvedY0RyAvFKew1tgHrFLaK
NXKWucmNo5vFq6AsVOxZwN/lT7TX+CvkWgnJ7Fp0hi4cwBGYqlO2mAAKHpU0E5oLlgIw7Nba6vpL
4xnCGZTVwTJ7P1EUvXKj//H68xrttLzP56PW18FdwmQS0at1jWRT3qOUUBbeEKtzstf8l83NlzXQ
Ub4J6WweBZwKDQb+BCLveKtGtYwll+teDIQwIz/UUOhNPtxKwHUhBJz6vSX3pVCHQ6WCdTNvo6yL
+4epUjXZIWpyHFBCWdXPeHy/voeESj/7KQDBELYfPXBgwS5l2+cJyc9bDD5YpD/20+ProphIckzx
cK2LbSNnMONVul9JOQ4yuO0ovkrBDHC7kemfajQOFldijQA/Vm07cGRcpaeZ+sLd3rTNH3/H6tZD
KsBCVDJ/cP7J5//vE6BSLg/Ubq7cdFqRLw7+jEA7ok5x4VcW3DSvjdCKCmujILFj6v+5yjOtYBNx
LtwS3C+zE++xSNwNuM6lo1pr9p52nZ2PxdKXJIv16oMoi/+HmZjEI44tvDjtlvFvoxa6vxwzLHw2
Ws0OIkHbNCOreTmmp9It4se0vyeiG73yz/HNJpOHKcY3gMdCoclP5+l7vCHiuaIobEy7wTUnleLd
zMVdi+9oaV4uQMy+UKoKFm94gXozAhPvgbTDu1uTczcmAjNHJNBHYFBgJA/gMxkCB/B0xeM63+EC
TTf2d/1u6zMdTRn5ilsmem0PVoTpHOLo/JN99Qd2Qu6Sfpfg5gTrWhjz6WwloQB8glRl1b0Y32Fu
xBoEzndYbKCtdO4DcAmIdhQLwTU0x/iDjHu+WbUf5u62T1zECgytwTqgAizpiovDRrH4bc8vRTOL
WSmeLQkVTLf1M4bgGoRqQ7XCOh9iKIAplzSoKiqgBRGuD+Uy6aNSSKoDEsJ3KntSA0rZgQFQ+hiy
I0GdptL0xtKi4cvGlKTM42tV/Z2Pc1NiWIQRHvRqvWROpLAMCdQeJfY3fXhcs0OrDgBxSuqhKXz7
/RmBgthU+mFQfYFXKjvfY6qyzuBFHFgBeKW0RliUTT+Aj8X3WKEuHQ01rGF/1nbhw6DkJhqJwtvL
UQDJW2vjl3ikdlRBFFEw6+o6XM7vTO5PpfemkHDBKyh/91kgorzIAEjDBIrJdzH9kgl6W2mh+sDd
LXJZTenuTumn1Ds8DX/TFIdtqFoV4CvvgRRlr5HoYpuN9pxN038uN0akiQFmVtGpOH6t+3R30TD0
ELZ+jcwtuOQCX3N6W3n/rCbdcrCNJSSgOhfqHEuUmh8eAG3tUrCPiyk71UzEClorP1rRBLXPyu7N
H5Qc2QI2YuE3oHeb1bLsZwsuus8k/hIm0YHhDy46+3Fn6u/xMy2jMp/4/qOfXvpP5tlro9JEbvVM
bjGB9Utqh1HB/0A2juSfyK+e0zfnrFU619C6yUY22CVvy7/Fn3gmevq/6r7x8HR36ZA9+1KViPwE
9UJwtLXmJRww77zZiIJ0D6R90Do2mnqc0g3n+egX2VjAt+WWTPQF6xAtlZi68XrvvYi+GbVu8BBO
Uc2OVRuVNKe4LMIZbeBDewnAUQrBHGFqciHwZCq9GFauZFKJOgMonLTrSQNzYIK5nDDm1gcEeJYK
KfvWTsOTr7wjRvK5WBGr89cxtSiigB0/UWUGzL2I+TWe/I21DUqNaP/3vl1x0UfToeC4N3Q9fTuP
vLiN3Fu1RN6hKcqHOykbR2YHRa5gbXA89doKbgLIEUceWd19NbKd3QFAIhTKrvBmT/2BRTZknZpW
uUIodaDJI3isb1ra+RIiuR6Um3htVdxLu+6PVikJ4Lwk58QMKDH1CneHWv3XV5sbj7/NskjZy3Vv
3Y9lmYYFZneXR5id1zWp415np/7PyUmbCNELS4dW+x40mInzrvAII7fCXWlvc66JtDyF8CeVfpQ7
r3kAm5ePq4Ns6tHnBxjm3HQipsmCeNEGquOHAxqS+jVXCQIQk+3K1Qgvstav28VLzdyD6XvSbPTT
WRV+VMAc2iyI5m02ygCy0g0Y9HTgkFq3Ir0KtMo7iLgw1BSl200YA+JWzDO1bMopnAH/sZMIXxAD
Uwb8ZtQBBaaOOtg353p5Dnn2vTlOHXkbu7hZAfpH20dcCZkYcm76FGUNX6jtxFrCUdpCntJoic7N
CpCfhhutZTqaeN3e/+F7oNDEOKtJpmmmnXiZz2aFa5zxVhxGjkX3rldLQI2LU3eqqwh8CKrHslRt
nZkaafxqJfR31O2Gw6R9VQYcgc69Aze4Yqtl8qv9wrNu1mD2cMmT1VipJA8qh3rUzq2dCxZPESVF
fk9k5Z4dwKC/r9/XiiRRATRYBdOQV7CYuyu7ykN+GYfvnAEQkrCFMiJl6TbHIQ7XbJPMdudEzmLc
kCfmU6e6t4zmSD09kjkkbZws0FYoaZUyu59Y9jAqBdAlshZjjl5GCY1JyfE+pNI811UbTOqYXQ+8
LTeN4hWQys6oc/ec4iHbRwpdTBwFlhmg4tnY/WPMZi2v10+KJxb7cFX0aNG5GdAWq5KyCoVGGom1
fp7Ecl6j2qhg3Q3ugbdDHbohpv5gp0eX7ynx4Zc+HEfEnayk2QCpo27Fv0BBZtrkIFDKtT42qetB
i7/bMh1mFMj4HkDunkNswPMKcTUEUxa3Z6aJOiJ7+XVSLr2g9D2nYjGXrIMH7u2CGybXfJIM0Jn1
F7u9a4sszDpXtR7qWdtHIfwcBh+fFBskpsloIGMjS0AkCpRYV4+zi48SW3mPo6MMXuzkLdVEPkE5
xb+ycxudNxFXduEXR75Zjf1KhrQsrsncc1sCZDcUTw0BYJbIZn/OOQF4IY/axnXWbd3pihSd+RGD
AGc8ENkJ5LV/Z48XnqGhnGVYhz77kQbmTlJ8IDy6Eko/lPKe8jSBzbW8mZGahj+fC0AMc721Pbln
Ci+hQ3SzJ2GUnOpQI3wlZPtwrfMIx2981EJZ5g7v6Ja4Ypc21rxhvQByEExfyat097TOlpLs63YU
PuaXjHViK2diJ6JTwkXa+Q3IQPgBs4cfBvURdakjnWnJrAnAs6t2dKhSyIF4eNHLjFK9mVQ+FMrI
2DnNznZ3MNgn5hDf786rLq2OGcRfN5hYO2wKE3ElClvAnLgGa0NvYRp+EkMMPKExZyHEYMRyahmQ
bIv4hL6y7fP7s9sCkzavmG5vkk3GglpAbW1j9fxo0y435TcnwgRSFTJnNhkCDoVjMGwBsaTP6fJI
BGaeMFgMKigUdijmMZOgWTkQXuusBBgxtNB8YoRRILGawFbrIE92dFb3fD60eRHqW99CQxXXjU4d
jXnRnfEV6q915dwlcxH2ZtsuU8Fqgu+z0hgTM1IrQunq7N2Cl8AGNrjXXfuPAUtC40hZM28JDQ7Z
s0z7bP1pbjDr69iyElYiqzxJnTVCI7yYMhi0Ob0WMY6RyQWoMb2bI63jW0N867rKu9gGko8j0apd
jD0Fp8/ClLH/jvF2X72dkqVDaFOettRN5MeaR/mWkCjYfpkPnbsBWruyaJEexsmWexhCeHfsYSFr
CcFpshdWZaQNA9dbzLlnLOyNsnW5hMJbybukXSzDTEl/8vcFVsjnT8UVlUnePXtMDShyYWMetO7T
N6RQNGpaLzq5YjkIMJZhGgtGflncqvUCEFL5N33QgVZLb1IXG0QoKbYd2fR+6CzZtTg4ClVlxXxI
Xfzy8QLpEFwRkhbX21T78JNbjkUGzqYU3VyocoXoBi/q/lXSACACr14z+jmYuYBAeE4BiQiX6RQv
CYy81HQLH0FNExek9kDBIKteT7hU8ty0/Tmy/UKhjNlr25gbcqQJzRz2+mqfQ29G4qMB/Lzl7ib+
jPHVVXXBQx4zh2E36sjdR4qW16bJ25icx9H8aej1BpIyZbpUGJOXNdcWUujd519fwxsAoxCmKRZj
zsPlFiLs1bMrdRnWXQMbqIH5kua8ARsiczrKZwXF9nGI1enXXTxDK+5gg/Pq06FCffz6YM+8N1K8
1KwsTGg2PxlDW90F76kzL1BWLgqRyeKBP7c5AxqdX6mN78y7eETd7Cq+yAPs12WZzK1DIMsG8Wif
VTRdqtbonAJ2qMzMEsXJ9u1UvDiiDa4QLptAPourRE/lmMVMHboxVMtWh9W5jfaFkHRYwqOIrWas
EeLSyNdiLiP1Q/11WS13Kva82Ns2MUKydf/AFQFbRRgBB0cjntgyKGR4BAtzVG1NPDNQhY1RYsQM
NRbX639V+Z5nEClQZSMRTuLlkAgiJIWQzGz+3Nzb2nxAM+AmU9bMHve4kOEDUHr8aaQjSDXUl6Ll
6O0X/HEaEmBRH0gObzQ+uOUm2tRffaaA0CvCrI0gEO6QnyawebXdE+iPt6PLOH9S5MYuzlDTbHUE
1g0DOVkJenW9iJSkBceeRSpo4dsLuorI4CC7mxiEM+3nGqAxwmP484glPDIALDZ1UMaV5sM7lMJn
e3q8Msf8vt4ZlY2GASo2cwJ7IEwjOx06Ui+L5updl+7lr7iblAuqzNqQrVFbR2N8smgjZ7MyRN8h
vKH4RdmFoBKH5DKSvAAIgXDZPtNGGTMv+JeOe3INfGWxJzs9ONnRMj1PHPGFVRi1SP8n/rm6A8xR
ODWqNnCmqDiM5cthv23+Lg/luWYT63nFNhHrI2W3PUJissEpvohABE+k7WLA31YkMR0Gy1gCxZ3D
8ImdeTR9pjLOeoMfGNYsJI4lsv/6Z0ivyjQa8f4q3NwlrsobESDjYNm67yMlF2/p80k4rPwAPCZa
gKzTyXEkah93B4o4iYadlPrNIpyNG5ONqxtf/wXh3JTzji11kKyeQsa3EqDw93UhyUSpF3kekb0U
nOCdNUE2LKj+JuW3s0xppRHmclbubN+FO81LPboJkbBn6sIasK2f4dyMrqhoc6q+OokS4O/zqbUn
1xtg1Z5p8xYHT3/DMCaOWbZL42gffRzILQQuvvyHa6cTim18W95TjXhEivQrnADsMaeUAP3q4Q7K
spGqFBsftF/dgbeJJf67yFcE8lT2UJbSU67Y4+Nt/rYLDC8P4x+i16mCG+fUJ8osQGIpjyPY547h
ow89GGaQgy6xcNYjcU+d35c2ztHaMQCwowYqVry+Veunai9QndoXY/vjYFteQ8KTIv0ad3mGhOVj
It0icw7x89EgXILrQOopRRVBL8/Q2h2vtV5wXeYM0gEQH/7/zfmFC/MdvW5X/nZsVQgZSQs/Hmds
aNnmNrZljCaRso8c8SsYAFBCf/ZHyaKaPt6vEka+wLrNlmlyKNnsao2He5ztw97RebV45culKA6R
4drJx/ag5P2HZoR8/wT37zwERLWLNTIasIGZrDe4Kl8NHPZ4jWU9wibo8RCaZE/InO+OvDxvrIYi
/R04z9f7E0nI7APzhzmZzrouiKJ5bGoT9WHNVK5mVVZkIQRxkAyil42HmwgP69rEA6d+Dt0KMUuA
r6PEREmTbsV4TkYtKNPF3FWkEltjvDipccffW73BxLxdZe7xFBEEWJ7q2BgPMdHiNNBsrlPP7GFQ
jGrxUBbT6RFwOizGBxFakV+IZ63jccldq9m/r9BZBTsFY8PAwdBOuWyudn/qqr1dTmC59Z4dV5s5
YzEjq+y/agEZ/yxKSbDXoUNaDgL13aGy9GTvbtimT6mXfbFBpZGOgwCn8T0QWqTojLUHYWxyipn1
JFFcI5iQlHP+fujVp2UbIMMVgNI6c6qi8jYvHDImTEhs7SkZx9TLwzmCAq53WIQK5HhrDr8SzeO8
fBdDJL4f72+pR6f7Py77+QqAeuV/+Q5o0qnrro5LsqfdZ8qrROxMdFRkp5/lChL68mwyyT0+HmNF
AZAtFKp54Ln/FzKJO0+1kqsLsXW3l2Nn4LGx5cg6Tqhvq7syJgoh1TWplOmd4cJpye+EsxRqYFzl
FdvBIlGYc/IeqGXOqGjSEJmroD3PC6vfPeEpR6EriUjK/ssDy9voHGaR71pS7TMCoRY3O6vmerYu
YY70WJpU5wRMxa7iJ9+f3RS5JQGrg+VQuTSCnY1x4t8aoKJn6RNqZXJceFdYTHf27wm/ucUnsaYY
sasz/sjKUVTuX4r15CV29tiaS+/lPtnJW3j7Ty0MUqgCkEn6toA68FUHIWo1HMdMM++ZIy0tcJpA
IwOeWjs9dc7O8tvplQev444hsfynh3HPnxhDNGaXnpqGilQDANqAL76K5+w4eeqe2hykF13oqIdu
qpfquTEG9q2ENqyMlmTya/PyLXidDlb4vRvOEqXeTGRGe+TU+sS/RuxB8jfBXRkYzBd88/bBh7x2
vAkQV9XgeloekjHFh0Vz/bynUG2fAqKJYjm6BeCuLMryAQGQ/z91adEP6N8JEyJ7Zadra+s9z6SM
FnFFIiItfr+Id8LjtXiQVCHLrw4qtACGt4IENUXY9sc8MM5wP8uYGNwKuDzwSoKQCImg5Z8pKB+F
k3FWBR4mDVbBIoe6xr2eUzSFDuBA3P8eN3idg2MZ4nDrGJ8XrpclungdrQWdgt1iPCBj+M3ZkrKR
ewpNbnWrzgpgA4XMyCkHAZ7zwWGNlITIBBOJFVJU/k1PzlGwfRyImk/xHE4wd5iG0OfsGuMlEQTR
68YkWCwwEv1wgW2GE1X8eTCNO6N1huJznePCJjfigibOUrCYyxvsuk8CUipxQ1AZwMikeLQ+rSe0
CRCTYPPp2qD519RejDPYSMO4v/tZp71OlV89kGP07Xd/6MIlnWomNItvZ1Og77GmIrVEBqtp9zcg
h992GWmP0iHve750y0wGWj5SyvkcJhNqTrbwigw+lJnhFJaFwCkIgPPtkuH7ZsuuxQSrjeV3FRMP
P5/hWdJbEV/X/4vbwWXsQM5bcL+ypTMRBoZlWJYKso800T4sUznn1ulQSfvswAH7frqe8JjyKuKe
M9MuvrXxpuctR85UQ8uLwGpH1odzLMJMlCvLncLxC9Whl76WzkG40eFDsN+xglLS5L/eHAmSBH6b
dYi4G4KwTvIvnf79Nld7Dz7p1vp5y5lsquZaVxbGlEBKcjEq6oBCpf+UUlSAwnLGvkJxMYAvMRwG
ZfNFrvlwCI7gkzwYrhZBVTPEV2bglxKYzxW8CjdA8TxLOA3C3mVCi2hZpb/tYJcuNAZ0QAUEGVmF
oFSvbKA3fd/h/iTUoGLOUmBJF57hHSODdGn0cUwNJxU0QYHCXXeadplmboON+Mj7TjoJknGrtI43
NnIdusQC/nnyYcRfoQanx8LdRIGWWf8schX45zjkI/DcBUZO32M7FBqKZ5qWM+uMeCPJKKcUN+6n
nkN8D58xV7IlavwhRgVuvyztSijv4FTl4Cxk2gqfYaGKfB9cHUBjbaLSQm5XpzzqkVPng6n26ChW
3FMj/9cFJsU+hgVsg4SAqRRDId6GIQwbImLY3DFSmDlW5oQHKJY7zRfk+NwGcN0ziFDK94ES4yeD
6tpB0qh8dd76Tc/jfOAbNIF7LOSYGpSD0n+5eOcnqAT7pw0xvQuRK/rLb3lCkmPa9fhDRZttk+pX
jZJ8exJNM0RkHCw255tvfFAONef2L+cTp+F8TFH8MHNDNl8cUCmV7E4zIxuwTjkvcc7flrlrni61
bw7BS3yHiZiOQWjA6bsnDMdnzTJ/0rBbWx76gbPop63i8jTSTQpGf9NK17MEZYOB1+eIuAyDfh6K
Q6/6Q7z7HBzS5bbnvBT0md4E6dAvIV3p577zNGkcabiO0DBL7hzSEp8ev9Y6rTIpAFe4pKU1EtYD
bwkGrdUOb3GiDhM2uuyRPyWdauA2MJPKjAhMs62vkwVbfSm35qcIV8ufJfbYR01+LS1GiN4KhC/F
KPWgEstxX5Hw9hTt0SdBJahPmihgbIQ6b3dytQJyfTP3QEFZn67FkBlBUXyrQbhmcqkcyimfJk8x
CbT1b/DVHFG+7gpqcskBRejm9H2tjFrLml3Y9TNY36mS7T3CSkD/VO93c6NFolddNVoJ05SZePsJ
si6o5PgjRmXi9M9ORFhS3TcpqfymlyKllezDbd3C/dQL/jPafk/vgP9P2kKAX5SA3XIaHn6Kx8Cx
iDVSC87d9e9aKOiAiWOiHvqx8AIRU7r3FRxJmtKpTli/+J9jaVer4erqPExCZtEEYdQkImDPBuOw
1RHl2XKH5JEE/P/b5cbgtJxo4ySQtVpjBvs0Y/oB+35RauuEdHkuC5eb7YPOpuf9SQ/egRdVuS4Z
EZ1hzCYsEeS+CQ74k3pp0Az4tMpRmCfWO2j3yoePhz3/Zk1+qqpgJKjNo8j5dKnp/Bg1qYAQxnUa
coJNFtwwqeVNS085vfda9/GGRm9z/xvJQN5ZSmKRr+78TJuOezJfTuA0Fwwy2gUHkpbpNL+V+V6J
OZDac2PmQXqT05KrLYecyEhQg6sgWoq3QLYjGk5aIKy/LlAOnTJK8F+5x/uF13LXSo397Xa9jG2b
ie/OvrYmbL3Wuyq5Zb/iPkNxcjWJ/q5ogOaATc/GNsSZP8rUMX8Quv42U4lhtQqst/tLBeT0A7gf
1g4hKmbSuPvR9mwKXdzWhslKYAnLmqmVwzKpLFhFkycu45xQqOxKJ1hQqMIalSIs/ZX2z/qyaeNb
ySgPx9j43qZcB9+nEjBSdbyMPhWoKSklQzqFVrkphUgbDdgc9vgMkx3RDnCvyJCfQglTCuxl2MXO
S4EKQmc1p3+KEShY3OWSJ96yJqk2xMukuZT/XrKt3ihbmyZIMqE4xBWWlpOvQLpR2+IIDBn3cZS+
KYj5F2mzs49XbQksFUDr9RZypgNJvnvcHMFAyAAM4mhCWnOuHFj9qeHzk+rh5NWpm8E7mqAiLA5T
tQrSV+74l5pXPYTh5V+y+ujx10lsXorxFibr1jvHuR5fVvEGKYGj2SfmrcNfXpuOVAyr5TkRAEmA
MhnjyeLprvRPN+OxWMVCsroQxIttShUdCxv0eXVocSdA7psJismypXBsaDJyLqlJbry6fOdiVfiV
2QqsBmT1xm3YwI9GHGJD0Tpte0PvKjJHWY5O8EWwrnf+DQ/7Pi7H4yVwVo/RQ15GCVksJX0Ap9dL
8F+nnJNrtUfGSrtiZpK6BRl5PqXMXGS0JwtHLRxSkPFGn/WWLguUUIlOfGhuPrDEPuTz/+iB+vPD
uTP9dGIDaMXiGLTQSmjaJCkyohN2Sry8CUAyyDDkX9uKAPyURLXuu/6WCWT8ribbbeye/Ck7BLAT
7k8x94tJXM1iSa5rdhQb146J68OjYLsUoJQz6CEmZoRcBUNNwlHGzr0hLAQ5Viry8j0L0LdwWSIX
QtWVL4I8l7UViTHtXg7E4eAAZ4ed3CG0zmwncWwbsXCPrB7ol2IYy6JdxxSV9TrV9QWTzN7TwZF/
UGOFkPRW6Ln8uMWR2pYRpfDqgVR1dEb6i5thBENuYqLdQe82X7ZeB7ixCdpyvlGovEmjUFeIax3H
5wRpVM6UUnKKye6QeWHT/rZw0T2+0Ck8GPNKHvt6lQkQ5nlsptF2kzG+tMsLOP15c8F4ow8Iqr2t
bl0mDcEbx8jzXib84F+hil7kVZMyRu4ngxmDzinebkNLfTpqXBkjNGWef030CZrAIE5RxM9CU3Ip
WYYqFEuEKtSsghHtaFrTsX0s+5ZSuTdjiHhXWc7Jyzn/+Wd3iI/9ZEhTcIp03jag3fxxpxVBrOjT
dWswJBg3aBzuhT80DxsYYp/hCG77dsAJ+N8TRRGt8i8ciTqw5QAacgo7Ehi+jjT5z1VgfKI6pUBR
rcJWKcJOwQw9pt3WsbrzLuiujs+L5GTwjFHVgYEiDbizxKFYRmvg9i2Q0QkiP47ayTVioXyu8jZT
rByV1BhWy5ciUkCetnNZBPaEArlYxZ1Be5w3D4EgmPwK/NkTSsPdYTzIreIqEMIRQl00cOLkEPwh
31fXXtF3qW2IfIKEETKPUXBoXPN/EQgJBfsPY4rwVbmw5kJPIJS/1McYFrYwOP+ejChwIoALkjU1
z2qCvgxLxc2iILf0zyqUehdqJ9SiDfJdWbQn8FHpyISuh9foyj0CuYdpCSto79LGRFmnRmGkxJd5
1lDbwMrJntSXUcmMV9fNCD+/KgFNwOGIlpfW7u2zDaGPSwfK+GKUgs9jeKxtyby+LeO7FumQJCda
AvcBCFVA4rugU8Zin+Uu8x+PAhgAx92DwlB+W4X7duqWVbWf5xvTXkffd4OhAKftzgCt2Fr+QBn8
bTHXlMXJ8x5671K9K98aW+vOjGSXF4NpSiSLjE/y1FxgYBCduwL5w/NK/ncg7bw/KxBGZKZfUfyP
yZ21sAqbvatqgzHHxJKy793GN1LssTjLHnCQLwOSSnItVe1iqXZWBvqE2X25bOupcn64n3w3qrmF
Sw8F0rjEogUydc/eTCyJolztsy7UKAMn/NXZVS/XEX5HxAV4RGcqqKMdj2+HCCPMg8KT+At6RL5V
8f/68Oi5RZCbeKntV9cfahKDGrCQt2uH/r4IMIFr/n4wpJ4oHhlTyS4Sq91mxukdOXEbrXdvbXWx
ErMMtL6HudjRIUmDz9TW5SPcOELHm7QGh4dwGXyIvy8mttQWIbgJ9j/lqGdNtSPFMY7RCW3nshCV
EEgrODO01cLivKGvZdCb10NTNFVtxu5BuCDEeTRbmkqlfIexwDUa64kGpDWZW4Q+fZxaUVGiEnm0
aFfSlerW7Glca7atAx/iMe+mrDT0HtICDUqGARF0o/fCyJ8QQZ0bZBD2TndWYuFuDYjkJlipfG5h
m4Wbw7VzxEcpwjFbsEToKNdg1GB1Ci3xWR24WS/YpDZBT9jvMo6E1iV/gunhnGRLPKgxCMNZk8aZ
NcH7cpaMekSQbK4oujEmx3mmkfP13iG5kaYbONhe/62V+adRa9EO2hTZ2KCXwYWVHR+oHp3AgRWW
OLQCBpzxvOZvZgGo3vLjswXqjbebOo2J1uviqSbUr8RK+nOD5tEKpkFdy+Y5HcV23BLEaS75R4Ue
EuXX/8oNdwULflxHpqan92Ua67T9bGZzp731oNFnAICXUlZ6YwdsTcRmvAw7QE5Fk58xXJnSOkfx
v6xZoAGAA2L98lVoLnYuk20h93I8SUgU1j1XiyJAfMe/D2DIWxYwYUjNUgAqCC1j32I0qXlgMOmf
9DakpZVZt3jak28TjDags0UcLDu60GBuCRygUP/HUN2Ru2rsZG5sQDlqEZch2M8AZ3wTA8Nh5mM/
pecvudxjvhZl8OjG7pC1NBk4HJSsLa/DfLJchLNQk/9yXx5nlUEaF8a1VxOT/vvgmcCfdj3UB6Nk
DhPfSzJU17vi+ZIpc96TmLX2oDIl2D8ZejBlCoc8k+TWxOCdbzC8PDgT2n+VUQ6yL28R0qd1TJUE
Ic7dki4dhcOQ2JzehFwSjv20ob2LlDcMi+S5ogQ+sQMA+RFJuMD9tqRTSr6ZW/oRtC2o29QcfuDm
zFVSNqcSTdk/QahnuGd3P9utudS0U3aEHr3zkoVGjdNA6jMu+RRuaMBPiOxbayLrJi1mSe8qCC8D
eT3ckUXyIVejY3XXLaxg3v4Ja1hAGove1vdDLx5sXlzOYcNfTA7IqF2xSoDvETfp1NL9K5h0Vuto
v1tjsHvdTLO1BYhK9gXUUfZ9LOufzJSabflzbhlPxuUPDxtc1leIIV1gyLDL+DHvvGp+rXF0Tdl/
IvpE4HPqI6+iSAYLvRu/Qs9zWi/fnYZhmLrr09AGuxHxYiCMNuBZ3aZmJSetxSPetJJU2E7vCrzh
7FQrPirN5f2QOeeiJzZliksbNdX9uc1KQUL11aLTsrIwaXdjTVLkCAIoaac/dqrWHO01uA5/vjmN
tsdahqMuWh876BjMb9d+7KUiLFFmEzZtAcSdPFS2rPPu6n2I2rCdw7iJZLlLe/rssQIkKlX9OUMl
oK+SoQ4HckYyerv4GlyQ+x+ew1EQkTYXNrQv80zVT+qkLttiNnHHbC5eIX93Tb4fN4i/gVmwGr52
6mwNNXI4MMN7srLgtTXZXT9YsvdMVWLC6QG2mOK6rNL3zzo9sosPtmOdvZ4B8PqKo4DkAaR56v7h
wxsGZjKQU9KXddmL6Bz2BIa8hTymaNFfRhWgl3E3qIcuCsfb5rsJlMDmIqjvXyGycIFxxXovPlZs
76fJobImwiku8Zc5b7cUmyVmCBNEsAoeGgZERcoBEPrRfb1oH4zet7exUm5qQNoLn/17ndjsPVdU
Zu5B72uzj136yrw9D7mSOvMVV5s87SwJKhdJx+bKm65WQCGc6L68mc7f+IFAqMgZsKguAWPHFc5g
CSnbIKj9hUT9LjF51vnXnMLCPB8jigXpvdommqY2QDHhuJkywfy2XbUBbCa9qrwkyhpWMmwnvL8+
7OblSBYPig2hOq7iiccOXzjaAts9rqtOBn9q1CE6DQygWk698NT1z4RK88qroNX/JpHTMnVIwkw4
BpVNX78HBanPXAcMQ8/Tz5jPOcMJcdpF9UjbIy4KSRKgRiaN5Yv16BiXZFom+ryFRHytN4ebbyIP
j7Mivh/ZbKWmzQjYQ8MkiFKmtbtEAOUT4/kSvgnI/4KACEMr7dNZs6N6bvcO2z+tfSl8tW7dadn3
QNP9dIoaCIbpRHr8VOTutvaM1ZwUS3ZAOIHQj3JJIib+aYOugt0jA1I/7KSul2C15DMQooCJMr5P
91zYIczl18PAqTrSCWvqitDjrZ7kX6rEAo0NVX3xz/N5NRgnlC+/BWvUOWb2+xK+UvRdyYIj8TWm
4NDQvBKe3xvHuecmjs/gIAjzW2N5vjEyLTsI5ajLIt1BfzHEHsxhnvC050FDOuMSHnWJnAvDH3U5
zbHQPFB+PXN2YcEOBhEQurnx8+YKW1kimkjlJTczbxxPDLCr8BMetYvAxjSGCHlRKDCVtgxBObRw
H+eUVtOiat35fR7zl8HuHZNRSVIQSNdIxK9PYiaFybWKpFRpU6J7vHym3eGBo7hdpJpVlaP1xUHr
PzR9c+gFdz3Ft9DM7atW521VLNpnVAuSbL4BplNoD/eDOKuMDR8WCeS7spBcu+itYci2mnfMeqlI
D5AJ0Q1B7E92MSMQ1Wi8Ham0SvswIddLjyXjgnvXRZ0UXEh9BoKZnOvC9j6PFXIBQ5xSxvQ0WsBQ
fen+zCA2elEIi/Oa7u+9p3e2aRybi69KLHyvj8JYsFEBjES5qx18gjrflifIXGI2Rmc5QKtLJmgK
wk5CTXjYNCcDz0EQIGDM9fZRfySAzg6hnfVcA/2JDtJiZ+INgTG4q0YrMvXKBT8Tu0lRSl1pbnFb
fSyzpmbdKI6Ptwat/aBCtGqXEWuOX1ZYMHIFd8Uuv2ALNOOxN0N4kZuwJeW71iAOP5w3B4MhXqOX
v/4YAQ1LgsBup/N4qsshYBq83UA/AKNXWn1hKKLwwTuoX86wiTeD6bMP4vV0Sn1VcXMtCKO4bVNp
f4ySu7pL92VfhkF2RW+Hp8KrUAts55O/8SkZLcZFzYHh6n1RWXCJGlsj4YqKhOpJNwd76sh0Wuts
yI+2bxwyGKoGCx3v/C/h2ZL5aVYPXzrlly6fEZrBqK8PgmmdQaHck+yLMlE8gIbMwL0Bzqfxi91L
6/ehLaoj68fJBCll+gP+qmtV22ORmZBfRU3A4rjevSjynXseW2Qjw2aiDgdD9QRcq8AAg4m30PQ+
HuYVafC34dHCtiWERnb5cLRHNuiyiSfKL2ubx2+EFQKd32GwbuYarGhkg8eyRJBOXVO8cmzPn+EH
RDbIkw+hbyoSI2TBvaXJyJHMgBsOXR79Q82FNVSX1PuUhNkquQqUO8l2muZZHveWje12wKoVbsG8
nMWa7xpAybk6kWI9s100B1rjlfC3vE82ofAoaJ5wqwKE4G0LrmDCQcaZ9/ykm5QqKQijv3EpVam2
ierUkCb3xQzt62pSAp9fmKSpN2ygKf25EwED1hW+iDXmvVU2R3xS2BmKyBYYoQzXA4N0EG8FyjE/
ria8QawoOpvoIij3XNkJo6D+4GXOO3FfO2cj/8Wc67/uK2HH8NUnM1wnHPBUYYJL6S2AVkQ8iZ0H
4DABLf/pIGSZS0Sq7WeOjlVPzJQDOXMCt4sMUflj+m2o41nErEYvdffH0LDF6zNJhB6NxX3gruoZ
zM2mqO1aCQiMjcV14wQI5t5Jg2k9wf8sEUff3N+tjweJVM+Erwpbb9DWXjBRwxhbbcrx015+YiZN
Py0/iXn0rFQIE1oiT5MpqjD1RA0he+v380nW08zKCKJlzIifhL9M3aFFqlOZgYngOCH48NX9uGEZ
ku/nN/vt12d3Z91Ypd5tH8khiqUVhAr5gmCFAdKaAz8BR6EKPLYGArP9VldF8jFoYuXAbj5R+1Yi
EkbfTdk/SUPFRlU5VeDHxDIeoJnztO5a88aZ4Ivo2Yw/iB/0BX7ZNfHutMxYEayDw6TDYn1GXsy8
FCTj9lvzuggf57hMbg4zRjUtrtKC+mXtafvQxk2XF4qGRXmhvGP+th2LDA89RGN+59PeKzph+t8L
YtzVDQe3EO8vny3kYyKgP4jUXyK+mrcud6iBAjXmsNAvcD5WAyR+VF8MhZNleRXDwcCwRMhnfh14
QTWVwR89XjKPtwVXFVnhlTUrXKzy0IfIl+AKef6Mw1CaBcCFoWSe6GKfUOOai8RocQmtqGC3M9MW
PfD1TGn/aRKTXZ8ZFp8YxaYqq7J3PG5fDila9okgea4XJjbRkmpvX830J2LYEwpDqUwFHByBRq9m
+aQaYuzYqLl+vxo3Zo3AfLbacRLng0BU109SpBuCgHrX2JnycQ8/RVyplxmmG5ilDeGDThzuDRhi
YQXRkxXJs8h1rgxzBUFO1jik9kguMR2WsFPt80iT8NUTu0ZYTXYMnJ8Q6yG8lwVL06JXVqpToc7H
mWR1HSZF6IehuzgfdP8PAWxj0YGd3voJNkbQnGXzvfNdf+mVkiOLe7A5tcTLXNGm8bhXONg+2YCs
beahXNDctf8vLe5eEleNigOdetcLRoQ2WnZOJB3ZOJbS66A3/zah2mTcmbQJFHAWxE/9yCFIFHDa
p2FGudzXoCY65hq3XB7w3KbsZglG/tLPqxznhAsewJ7oItqxKCDNnJOCaW6bC5VPSBdTT36kZCYy
CKyFvQYZYINRha8mEr6DMzUkpCuNGCZDy9BqXoTEEhDoIXYLEmNZ4NC/m+JF+RDj4X0m+13CejHx
lqxlL+BdqbdrgMfRlYFJk7mxhtgENVHEx5ZGeBl09DvMrBIIRb3Y+tgqc07WKBq8nS0zd38Mk/tR
0nGuLqvLSqxXwD77lgpil3Nl+eY5K6JTVWjMBYkkoALMwcZs4+TmgAnootYh70wMhxVLRLBaA0EM
JRw11/6kVT2BSPz8/7fRdt8+WBR40Z5UH9tOPoHGnXnnpco3JNIC3ASFQ1ntBM1Zy2QOSAazycGu
3UBISPR9FKAAtQfWJcAlawVbWlI3QcFjX1W89At/iSOmPk4AHTzv14jfnY0+RClkxr3iKpzRbch1
tUT3jmq4PVq+X5qoabKr7O19U2ZFkypE3BKu8X+ZDRUgZswViUXhuVVRROa5mDC/Ua4ogjKlfVVv
YzKL+o10i6saictAvnQ7B6iJJNCbGzqkk9FPs/kiOcIn+2NjDpJf0Qo5J8aLDVVx1jRzFaOYCp13
VV/l6gPMYljUt2Qtn00rA72VKKLl1iUN2QLJPzlupvutGA9xtjxB/GXmwog4wh9WYIgJYrFJL2h8
fZnysZQXkesiUz0nD0FwECrkgtj9WSV/zbmhSgwvj+3y7Pq4zxQuOOwPNRfDeJmjKzkIOIusEpEo
rAEMpVtema6UBXEGC+xAR42eCGVKJeM2QEhOj/1HQDSzLjhMOnvsiUq9xqWz0kGwPEboOMbn0gLS
CSSCiLhA6I9nSnzOaHasQAUPmPvPOpNx+onG+8cdfg3rSz4feLY4Ahem7McpI322H3Dg8FuiQ5eo
JyCCy2YGzx4+U5m6a9G4SZJyuhSEMijWmB9WemOLIOJjQZrxd8R8AkvlSaL0DoSVJPsBuT8tFN5U
ECrXI5Rd0dDpmC5ghQIrSszZb1WCcFAcRCd6qzPttBsNSsyeNmZOxatyI3mtNYvzGEK8X+YkK9Cw
0ZfdG8ioImqqYq414edrYgaWVdpQptwensKvnRDxuJBSNi+wY0CxOgc78XE8b00GU5t86RZrm6wU
imRPbOZVW3A9TyqABwCiryEcFN9fGSylQl96LhrUFibcniTBL2gnnLbARdlvhSnKLdeMOrYf+8un
eFAmLKHYs0/dY8cXRaBEyGWSSsny394G+N8dRku2l0mToOdEnwGKodgnjqfX8cZejAJb6gZGSLvj
04My4qDA3WpQUB/+DR9kJqRRW9A8l8QoR3XgAPbS1FQOW80LqgJ+GXonyNEWpm/RLC8vS9gvnk34
z2Woj9hkaxu8KIvdQn5y4hs4NQmr/SJoeHAs/BH7XqX2BkRupW69vDgYo6MAoohdIWf5RYQz3PpD
x/zkTLtN114jaNyGHxeh2idv2s5P3tSEbIR4f+YHD2s08LsV50jh0kFEKakXD7xuO/cfUGtwUrWi
L6SLf5LLJP795gOzISq2ix/73Gh8hZwBIT2gI237Oa/Gihb5djYLRoMuZpALvZ8cjzkB45MYE5mS
MlssJa8LFNaq5+jU7rFSqw3lKBnpf2NuOCbLAxkN61hECZgZNCXG71Qd1zwmZLnLKP0gMEfmSf3t
ag1pCS1G0RLePWZvYVeca3sFOwyCaK6QoCffvFilhDgFE0JjX3aLGV+xivl3ZF4sRAtFFhN7FTC0
XcYbzeYVJNaO2ZO4OWGlAcR2kh5BoNaWGSOxzjbSUCqmnpjmk71/s7saSw70tf4B41toyW3pJk5D
3NfnIvHWKPTq72ytDoFvm/FH97/120RoVXUKIc0Y4oe3vkA0l3JSJ4vpi9Kmdkmm3Fr+x1dHRL3r
BfcuqeENTkN+MxmX1caMsbdvtZ2HthcRnRKKPFB6YpcduYf7QWmkuUgp5zprU6upe9Ii0dgb1dr0
bd1/ULnFOVDHk9QvA/OiNqjUsGWYnAMsMQ6+XV/oOMxM/B9g4PQcf1/wJFsuMYNWAh78FmmiNdJ2
3Y8b5KCr4kldcDJGEVEws+EOkuC0Snpei7wxkquIVHoDztRaW7hT1uesiYy737doPwC4WA9V+9OX
caPAo/BjhrS/cFqoKowIgU6iBuX2hI85WeioyDBtvSbXogX3Di2OgGBlQCz3x+Md77mVkamFKOd9
rDWf4YG0g1oZ5DCqvq4V/x0ibgF79oe6ZLoSQ7vM5CgDeBpU61JIx6l961n9F8risVkiW8KGcaIj
sA6u6r9ElsTsBoXMu/MyA0u+Nh7y78EL9pdMBWAl8eY21dig+4gL6zPRDzL7t9wGhS2TMNPQ4mSD
R1Zww/DoUBwQ5iUfpcl8H2MPnOOjUpidsHWFp/ZgyXwMDLvKsAlFCKq9yUOB8rn34Ul5xJXzir+j
Ai56PwqO7JJZgHFzai+KHfCz3j60YKGohUjgkHbgKVkRG/BZJyJQBGJ2IEa+mQwQh7xTU5bbEXPk
TDNLYOFB3xR3s2lQG8TOZCU0mOrYG4Qey7idS1isMaPFVmk6Qn60S80ZOaZNE9TiNC661mq5aLvd
JeENvBDYaTR6cqrZP6sjSnarsZWC78kyur1EeRUiupI+eQicqzi1hm47DEPnEN1OOoJW1fmrzVco
9jTCfWuUTTCSFbr4wnXvpHyaMCBVBfYuo1qY+7ehtN/j9C7VPMxAf1pdQ9X9UR90xKYFsXbhNK/l
ujQeGzBYbbn8JL1MWfob+TtEET9QCvWdo4uUwAackiHtBAfT3HT/oP0nfLhjFm26MKR02P+NcbkB
VMXZrfjFKZU/4XQy8umjWsuXrNmHfWNFl/rGDVEN3OeCE41ucX7Asq5Nn2Du2P3XX6oCykg+68PM
KHKdP7V9/etwqUYIoqQlSVqT0RBNxjdayARW47eKc/IhjYIfcOeM0xyHaKjI3QWaduTUF8H//7ua
MdnBb/2coKVP33KWsQspiTOWrnnvYGeeaqd3qSx6dfd4ekWcCD9MBEoo5a2/LwcZsmMeRX9Xw5MQ
P2c+r+XiwNl5uXJvkp/auwxbN2V9IfeJs2w6dEIwFMhQpxD4IBceAx2CW7TnByETeXXDvr2qR6wU
+BOpQ2zYjIl+XoJIp9eBVzZ2wSKYlwzCxtUtE5H3l9ck3igRNG5Yp4Sfcnq0XuXpxJe4l7B/GxuT
0dQBDzPueDPZFfmdS9bcsC000b1NE6uDzH2749X/iJDXs2plpSURopodRIdewsvjImhmHy4gVsb7
Z7DeF1KU/BAjzDqBbSiFOnLdZg/075tKnsUKvUlfWe+/A9jgKVrr+UDRiFR/9Aw2mgXmBbwPS1V0
W4V+rVceNcbOgFpLWaDDcT5MWsZMYCs+6nOGShjpvVCJqyBjpo1HE6YcXC3xInY+iFsiISMBLDv+
68/aaT9mawoS+hr//4qxfuZMJpywveXyjo2bzaTsj0Bh3b2Kg1mY+Xa4rEjYI5w8kMu9K1KLy5Ji
iC0i2cpzrl8JCOixGZtypM2vK5ESng8z7gZFvdPl+0H3fMdeQ4WBhWQWijhxvx9jD+eb6gkk5MUU
MokEfrw/dpW9TWCbkW1y/XRjJKZdNn8JuLFYq0K9to5AS2If/UQlG76Jjck/bhHOtL7CF/mHj7OW
m7yzIyt3B4b5T2Re+yFRm9z7X4yYl0sJ2C+Lrr2QjbTI+36ZD2Sho7qulroadIu2FRxw+2PJJhan
StA4zeg5mhwGymzwyuKz977wXn1O35cTdACHLuR9c5Lm3XlUmBVdlC7X2h4A5jpAxqexuqDc3/Ey
HwVQ26UnQ8+rX8zpOOdRTWh4keIo74LGseZyAEkod/sW4fQw+SFs7H2euBdk7zKkWXQNNjo5n4WD
iwDYKaD+UdXudmvqhqrYMmDB8TDbY4eH8HIc4PbSWrpC8pxfVGmOole818+F2NSohIYEFUOq0WsT
qHyE1BM/++GL+mFmjUk1e1bn/loPPlZ9cpG0rUziX10jAnHyhP5rqdkmjpPGKwv7efdo6w/WxUTu
R4JBH2ES5CIbsx5y4zJ/ErQjzxfoNRvjeVU/zTlv/dq+LQj9Q/K/X/8uvSqEsMm5fvhkDozvwtDZ
NtWiWowqMi/XkIJASqlIJBGzL8xfP4baLpgsbxZZtY/Wng8RmRcUfv0EX/tJwr3UxJO4RQ0PkuOO
hPKUAqGNlc9qaWaywC5SiJ+tLieAeNn4BXKO+fE3Yb7yUo/YXWfwBRrBSTVSdx4Y3j95Uxxvai46
z0w6y9lu8Mgzzgxy4yR4gxXhvjUyRf9vaIX3RgOpN9pFKu9iKcxg34U8lWK3Dm8XQ8WbHjirJ5Ja
Jzo9jfY+9LHroaHOCdh4xRfw7Fe2zwvo1WiiR29OndV2LXvlYGlZAM9DTHbGX9GmDmkL2b8eEgzF
Gx2fW0fA19k+MPY8tcq9QJxzUQnJVohvs1hqOoeEAKM926XC4d5WwR3li5dOv4jwDEOVCEHkkivJ
uewDUOlX5aYpvIibdCnUrxb7G5LXKHRGyNQhtBHIbrdyPrRB+kOx3w/gmTBOluwJdCcgWrJtPDcz
9foPb218Eg+EJPkUM3DM6uPQU3P3FBiPuDVimHG2/aItjH39fzLXmTOqCOt+G1GokhxrtmxhcKYh
trMBPQ+YG74kev79u28HgNLZb8vWKxUmAtrrhkn+dYAssNlI3JBWuspsRL0XHJ8K7ARZn4r9ifhU
/O3URsDG9CeX5+VPn6XoAZw2jBEF9IRCrVvFRdu0CgFIhPEH1w6Pew+UQVsHCFHK0j+AQcruQRWL
m1BoNUghBeOFOyeQ/U/tlpHUL0sWZIjj69WE94vjiUOytS/xSGk+gtcAzfYmymgDS9Nw3N4xrUcI
SJO2EQawWOJBxQRaSopzbs3MWe38hFUwufeuzMmz6bktrpVC5F0ztZmFcjoDTrGAH7G8+u1Jze24
WZ/ErNTD/ra/Ee+n7FInZDDY4ZTIzdF2za1FrkWC8VfhT6+8rJ6T6it5sX3e4lAmFwIpI8mJKdb+
ZPfKs/yw98EPnc2B4ZPKSt7iAFJT8yi6+O7y8nzaM2Cxb2/HSOYmRpGHh/z57A34+ERqwI6g6TW/
ozIIf2tTN6YR5n2LH0ViJ2o4v8v8gKV+SBhsp+bhI8Mfv3A32nN5yYyOm9lQBd5e87eb5PV19KQ8
+tsGv6mafMIHE0kHdJuq3tTzVCJZY+prFrsRD29MSWoT6IyRCjzTwv0NX8YGnpyKKB+C3mFPu0er
hzIo+F8ovAjwWiyU4YJiJGIFjbJdvrHp9NChZU9diZimo/dpxcxnlZwf8t4i4BucKXWHEb7gKBhr
tICcxbWHxyHOXoHzGaToReCu5TOp+ur7iSfQT5QvhtimfYO7VljPgoL20VFaTTmox6Te570Orgk9
zOJVhi7517SrkQnrZmU5NI3eQxfZg0OLmwLHwOkk1dUMKvhltEhcRCa3M6y+6AHijtUt7sqISPHv
fsW8i5ae4oGxSglRfU75XuCqWH14+sqFjEUv60Ew37a14ShFEI8W6pdgxfSzCl+YCweCkPltzGbj
WDlM9ExH85j1By6T/VlBsLvoYCgu4qcN75i1t1Zu7lS6Dc8mEMYoSy5GQ2v6wIumcAzd2JYemOID
UFdDwErYB8NLM4Hn/IzCMnWcbmSmXFynC5KkFoPJP1Wqv5heoK5VPvsst0TdzPBJjh7wSYmnvdhx
5+5nG7bXEdTU+GSn7VNT3jTv/3zSP7PLiOvvZvb3g76uDvYGTklT8bn5oNI/yMZNpr/Rx3Sjkm1Q
CMOpriEMNQ5TfKZnCO0WtxykOrVQWJuhHEWcMs7Pd/YuL+Ri5pFMdwuEImkCAVXI6clEC4o5a895
wVroSLmhytG1ixZfyTovyZxizMb0EYkm2/l6TOBirs1XXBJb4tFDBJriydLpFTw6kxGJ3bxIexEN
GRexvddo+aNh2rGj9eQjhhY85iHHPZQhcE9vOnC1yOJXEmnGD35huNeonDPncxyIbSmLIfYUraTt
47z76KcxSxmFNTr43PkY3/Pnx6bxeBy0CBI+1TG/4QbUK0iVyQfKvPnwrrB86rt2lB4JcyJubagB
oCIW15RbP3/JCN9d/DOIDiQ/dbs4lkCBY5S5fk9Vi/IasVvuHoZsa9jX6u2xKC7UR38RFhpXuz1t
pkUFnk7AZAV6imHB9HqCTATZxSQfWfbwgbUiFl2TSg8qTM0h767icBltLvfyFkGQpa+WZ9Y4aDaV
McpGKU6z9OiLh85UCRVEN462YNlJI0pXOFkjUvn8TKeztjHnivtKAYSOjWkjF4K4xw182+1DJJEj
ZepUNOVGqGdBV5sn4iZnyxgdovKsUh4fIm/ag/fMTwfUSzcNdCDKByTgQ74Eg6OMpEhZw8iwsaeo
B5xa4Gjh+hMX9278jIiWvI+BJfTZrciU+56GqKlgWw1UFUqS/sDn9WheoL8Bx8uDSq3E0ap0+Vjc
aCGv2GUmOAMURsY4wfuhTGsr6dVxFBTsYq2Meq896aSMz0l1VJGZ6382qj03nPRYUbMQgr+ERjSp
Pg6Z3Iv5aWf/xI97M9o4AWwHdJMy6saI4zR87NJJ8gKuUoCgn6bEjJNQ8q68keXg/HGE8rgB98ur
HOWNOAs7lb9nroKzrvRKWZ638jUoIfxooHqGfiZL+Bfx8YOu/5iGy/mpF/pp1sQrPqbulncsciYA
eKlaDqhcA1eFJhp1NjXct6FFE44o3qvaZNwQ5cdlRrvdH3gJZLlaLwIK37sxoDUWLGE+hlrhP+LF
5ZE/QHyLlSFI2rPQbol4I9pM8pFXxrwb56ZhTNt0QpNC7G2r1YcqmEBOGWttJ6hOL6sL+abfSz/1
xSqOGuhrvoopgbkJpSb7kaSdLS36HpOyZJxjklVbPDYy7NOHfHJxpJS6vJaxfUdKz5yb7JUyF8Uy
m0khngdkbc5CiLgi2zGnKDcEtU8+dd7R0I0TSI5b3dwF1DZ5j5cI0++SBbJluWnEPhO09t2aX3OW
eMT399wP86C/DfkjlbM3YBUwiKvN0zEeNiukWLxNPjHzQEriE8akMjMUy+FhAx0HTBfQEN+pqzKR
E9Y7MQ6jngoWvILd4Y9QXetTSTAO9ISjwGbfI9p0WUUUqzP8JkbBxCNVhg4o6c8VGEPrGZ/K1Rp5
pIvQlKDC9FLrjtMI6a8ZB9T6r5MSDZZpR2x6l3H6Se8Sa+WSZA5lGCZy3MXKmjCNAEst/Emkvq2O
+weWhW+YJMC7iYDm4sDTM36JwzQ89Yx6y0UD3xBvuSwwbbAFrBUg5pCzgamVRVXERAB19sva7Cpn
dmaZp+qdh4MK3qRTzx8ZWqrCd9tapmC5aC/+OOBH1WYjKKsSEZmP4H7aMXeSJHPD7RYpu7n5UjIq
64R2lPBY1eYy35srfhKdcKeNymJpDmGLjP5Qc3crfb0YJ1GzFMY8fW2n7AfxN+TjJDsOGI0Ccg6h
t1ugumFDcAMvt0lVrmtgeNtGzYDDXxvaYWvkFX1O7JrNIQY5rmAybjKphizromvWwnJHGssP6gaV
zYEuEVO6xoc3u2W1hvaL3cOkvoGIZL8FqpAowUYygePbBr7GcSlNXch6PfBbuSYyKzGQu8UBdvEw
F4UOr+weYd85GhwIzh6a3OohC1dk9PYxQRKx0s+YxE1U4L5gWpAJR5khZGdX3K9bKFAKABxn+J1d
ltRxh1tRjQNW/s2RcziK5bZS9m1cVowHAkH1ncSC5HU97hplu9dhbUhjjitLrQzZ1TclPy0eOjwh
n+m02GQr6KfF2D01W0Q0DdKSzY6JEO/4ZbORi8IukGrhvCLd1xu7+2BMWRP82pQPIupmuaWmXXri
iWi1fgco0ZVrHhKD/kDp3DBSNGlZ0uRTN89zy6RbXZctV9LQjzALrHwfiOXfeqsppQ2oKwJtsoJG
E87QGdqOKcWEr9MUS+QRlQw1NAi0ysCJENai+IaMqbdQcfaHVrgaWiJP23SyS8w6L7E5+p6cg7Bi
IjRrLf03TpZf2suh8y8kWop7tCo1Y50EzKAdM7GW5LJ9WPNcTKydWIUTn1kxOUnMOfCqllfRA9fh
G9QPc4CpQKAKyUSSZkFQqcqmcfuDs/bnqTqJuF5VyWBeU06ZdRFwDBohh7NTyBhvPdTskOXdHsct
MH3BCnvGoFLtCFrLplYE9ACfKsTRY6Q+MQ04yOiCbP0RfkbqV5637Gfye1v57JE6/LV1Jv00oDu2
yedbr5xxcxGRlot3/eK65zTm+IjtxZNZK1hezugIXSVlGjNChu0zdZwOn/dM99BIeiSe1B5kiH63
Xf+6Cz+LJDt0RAAJSQvHYpsfuXxKyyrlBkays9/HAwjKB09k//kTX/DPqkApk8giO/dMHD7LLleu
V4AWXk0z4AEAXhH8ZcLj52Gqe124XzcEZD913rY4vsVtw73H53AjlN/P7ugG+G3gcgbBcd+U6YS5
/dcLtNC3xB8RclJIGvdcHKm1XU8X6vpZtoINJWiDFU/GqTHamxXlT7VlDXAWV8zDzE4SpafyF6r6
AJ+/jrMa7e2HtW38yb+2qWekTCQ8uZbVpzYi7d1w1hQDk/zS70R40EUBuUNPXGxGFOp90r3bVkyk
FiSviuuSg7XcPw7+y/FypQn6psChecLkKvJ2epcTf5jcEyvMxlxlUPTJC5kySGoBNcvYcVlOnOd6
45U6LaDIbr/BvgI5CnuQ/aFwb9pQoFuErcrKMs+qQxGewwNF4DZhXRQazSlwl8DAM/GFXte7C6wW
bEacFSOdOwG3TYwXZ6PrNT/+5sra+HGsG1Qiq6kPz+KtS502BxcuIouV+i5R7zjxRTTYsxEDDE1A
OpBZVGxd6+uf7hpCir9IETVXmCDBOXUZ/iyxNyEUW29bpv9mbwNwkuRBxxcnHQr9UD+CaZ7fuSU+
2cYwe6gjXcxMAsMUcseszk2AYaMOtZ5OCKEVwilMwJp2jnKBuC3sZGcqfEnNuak4EZKtt6y0XoJT
rIz4IKkAZTRsyOs0+rGA5rfMd4pyaydN+mdx6V2tV5CF69TIL3xE6vI8//t5x85xR1YiM/OwL/uU
EZSXAYTMiMeDHzLw+tOUBY8ZgKe+ebWtI49jeJbWFcp8DMNKwnAc0Fwuw0O6Y1G2oZhpJ434MjSK
m+Pq4RfSiAaXARhdTt82sJbS6cdPXN3VMRUV4O5Ja2ZdNCjIOMyeBXFcHDPw+hdwtFY+j7mp4xU1
Z8cZHQenwD31sxxJjHzFBqIf6jlNt1oBc635Vwi38Saai3chG3QV95GyDGb/00rgLG60BqR1JojL
IGQOlMbQCZUTzJONhlykVOLjAAxkcsLdm+QZHnQyMEwSsSEDuJsKyc9uFFR0CNt7LPRIg3jtLCuJ
dJo7LZ177m3iqyeJqEuNmpIY8roREXuLtEgvXkdq2BVugiwH/5iFel2wgb1iYJYdAThzLWCglJwu
lUYNn1W3g0hrwbMIDcTP/PtoA4pacTMAUf3NxUvyzNbTbOfuvSf/DpqGdC1ERJOjfbT1yotmUUUV
aftZd4H/RzB5wgXv9Z4bYOtVjmvxmZlX7gh9VWtTthPnDwRVACDkfzWa6rG3gkfiUVe2nAS2JH2F
/A99AO27mRZ9HFEXtflVRVRMkzjsornOZ8TjmUzNZ6PnMh6qKylx/h93JkwQ7wCIYvD7y67MtKeF
2VIH0YD7xl1lYiHwOSUyw+frPU7Yv9eaOlOIcidjHXzFakikp4q/rQal/gzMfvjcQnt7ZAPE91kR
JcBrrualZMJD7x7zEQ02UjkWVmU9H94OYxm3/NSe1CC+36HcToMI5e79YNkrqVK/DWVf/uqyg4Y2
/We9WYxmiU/uraMjgDJT8Bs1zNBwwcOREaoOUFUQkXlc66HBDLwIKSMf48w3v/En7y09eHULdwPn
XAJDJ5xlY9SBYKk9UA+jLhfk0gRSjWKO7cnYN4Yhg+HlGeJNQPRweX21Ucjl4aumrDGzJC0OCgAG
w9DlVTQBEGXL/SkzfCmIDojJII8tSYozGJG5/pVWhxQ+T57DdoK3LGVv66JQdZR4/P/CowqYtHCj
kren9468pAQDL9qw4J0CxS8/92yzCoYG+/o0Mqo+avtCbkemITpvof6R+QluqEZkCX48SvG1FFCo
eB+AQ1UR9bnveFLwTaSDQ8XV4EsVXRu5l85OOouynkOZbx6rwqPsuEqq0HCwhHLUeoo75sLzwLUb
2QmsSv9+sZgcJ+D/VIIT900yI/lQ6GUhBG/uPZ86s0VdvSvfcusePdnQRq+eKLCXNFTAuGw5fPUv
71pqMVo4gGk2wibzkZdbHU+RR1AcFmQo4i92tKcmGdL2i2hidfFkBrfYAdq5TlT0cqYeIf5haFsh
oPx0RgLM0ZH84AoOJfsQaTlyxTwVGRQcIX0WxnbbbYEmm+bq7R7+vkZjxp9TldWYTt/ANILLBLoL
OHSiSB52n0hCOJGe6pOXc9g94vOtUEtUCBA9VNof66UDDM0eEmOAQ4EJLT3tPHFLD2vcLc1UWNqn
d2yHcYywlxWg0jJtEdXuZqLDDQCk+DhIAwMJFG87HOY6FLxq/64E/JbSQLf0x6wftH1jDLpEVZEh
frJq5fPzyGnthtBgDY/JHsqkdc684c5NlbejtsIX8gCgsImE9qOS81dhBlPPsCT+pyOSGlVuz8OW
1VLQiRTtYaIkmwFWrABsimEf1jzIq2/HtknKK2HYZ7LAKHhgSmXkSWkfSwlP5EWg8CLZUxIO00fN
ZLAdXEJatOoYklYJP7URY3HaxCZkBl+Gmf4HBkPFBYS1zqavgWCsiEftyLk9ToYQx/mgIc/8CK3W
u0WtH6CRvdMSPL2Jq4uRPpslDoh8AIIoZm8gvRO6r01j3imKKGCfhpvfuowuYbBU7HGCNdOvbVrq
nd5GfpxFH/73zfed/mfHkAnUcuAtPSWbpiUTFBwAql/WnU8IMxMxxu7USSyvTdoed4pwEGAsAnxU
2S/Hgj5tIGMdcU8TnLdLOehuslJQHTLV2v2a3MMS/tSJFzSZsWrp+Lc52GdgYf+9pg5838ViYusM
0A9BHrNh59NclTf5uOU160WuWIlI+ifdBSVloqVa3rkXPQaDlLlwSHKfLIqbB0DEc5CczDPr3t+c
U7rK/x1p8yt9lowpB4wPCKyTggV6pErxQgqOL6XLprqcKxjG6xdptscrzZ1DX6P71mzYNQ3M4zeO
5DcwMkIPv6px2XYqBzU2D38wUm4Efm0adItct9LIBz3Izjqe8RacGb6SPH5ZrZaLPju5323viz9C
czgiO7Sy52gUrzKTXKloGQ4oOyrQSqO0+YdDFmsF+eYSHbm7anDBHuVMqOqVBjHDFj2dFnghpssz
bxaR3azjOlioUv7a/MP+0ECPTWK6yEnIKMBUxeNxTsHgckS5JrGkRNlkkOH0M/IdoXUFH3YXgRIk
rzAi4qVsPnm2UZvwjbWIT0aFob23sY0V+IajyPvRe6YYC3Y7bYGpKvZ6F6i/frPYT3BeaNhrs9T5
ZmpIekRG+yWW7pu3p8tIlUHwBeoRP3rxgTx7SMoBcWB5iQi6U+BXwXjt4Dp/x9FjJyjMlrUjpFOf
Y81BjwHq+JlClcEjJva0PfxWxvKMpsoZP/LffU76zeB6Thj8PcoFFxcf7P0Gy2fEX2Z+tFlNg9i1
OUehTvsR9+ju1/iG3raFMmOX548xm130YOwkIXaSeoDd6I1s2goAHbMXU/bDcfbCW+hmGI00jT7j
bM0mRtyc2SFX73+XvQImD+w1mqFrvrDYz//jMaLDEPJQGQ4HF0/Pc39kNBdkiAnF+Pwk4pk9QLi5
nbZFqdxzhkl/weE1TPPTln1na7k9y2NppQyhp5c4oUFfTHINC0IObP/B2bMhezPT21PS7JwTyod4
FvvVrFlxxCy6k6R5uwZ/6vj0LjNCIleTZ2hVuqqg9biETbl37yTGq6lWikiXKYOvgLKib134rDqf
3JGfBzdcANDOdEzBo0aLHOIkfpYqWf3qDb2VU4Vs1jAkYmPaZXznPPK8W0XWam0XkQNCpAuL+qCx
JrAc5RZbrjCxNG7Md7uMt847CD6ngAJVI695BB2nSmIv1CdMmJVesiOa4aVFUSoYr1sLKunu8Jpi
57O3H8KgWMVl+qT4fUVHcpXnbSd6aWJIw4MgWgnBeRYi/yUWuNPohhBG9KjAuNdIltDvAKYQn/0A
x+kyGv3ehWU3WCrZT2Wk7QvKTqTxrAFvTc+QRZBKHmv19rjl7kH1MIVKO5jokHuabc5bvH+K8JWh
4tlkSo47CX6nLoZIJm6whxg9mCp0M8InY5ggXZfCp+HdK+4wzwCDfkzwVvN7eE/RWMLTFIQsqY/p
87aDJyTJLhb8mUeEqW1PDDLuNmWSzh1vWR4K1QUqgwlzmlyEiXlq4aJMJedQdRnrOwDE/dBquKwy
3WtQ3QSpRejGBFqpsvZQzzJ7miazW7psiPlrGEzGWuW0jT7hfKBOuhOF4PsXpvwdTHbKyRuiqd1b
5+CVAq07R7mAsJ+dmFZkKby0+uc8rRnd38KVgFkPUGlJ4jj3Mg6DxsJQRl8zIftaepkBbgnaUBE7
0B2VHUYRPmLq4SpkS7UsGI62PFx8+xtbbiJFGAlIXx4NUc3kozK8YF3sLFddfZjqLlahIqgQbLbj
f/L4i6xwQZY3xxvYfUVvsrmbfXxVPYHFhVsVQDxO+oF47LYUUHAc5GUc737lyVUwPPEIZeIsKs3O
Okd6kWTIMr/yv5/qivpFgQkT4HWFZKniWGO3rR0KOeNzr5k63bP6zyEBFGoyk9O1sL4Cojcv4dR0
dxNoqnEILf3K/CUq8R8OpUkrl/8slZpgcY4DjTgXILQ2EJhqH0+n7c9wbl0o9KKQ5T68eL4tN0is
0Bh0v3TGYdNDvoH9tCHnwrjl4Wkl3nTukVK0nmzuyrLoNag5t17lusq9KivOJ5ARlybiU3KlmzZG
WZlybkYfyozo+AZCKUzZf6HP2WHqz6ptCn6SdLpddML4ZEFgZa/U02rw1pP1EZlOXXxrr87yj2mI
/2V29UG3c4eFeYaVwFgjx+MxbeGtmhe846eGrWX3r47lSYKhUjH0zY5e02A5Fbcqbd9ihIcq+OtC
155O6Gqp/6Xn17Lv2pHuG9nYNVF6N4iOqdnfRW5uZEU1E/AbWWor4/0e2O8eDQt1a5HstwSczg3R
5jquNdvKclyKTg1AMOlf2BO2axv3IPgduGATO8SH8XdfKxVSxwVAxdlKQ3YBj0iM8s+TLAXpX333
5HZ0/NoVGZ1YuQrLYGxIJkvKAB/+ZWr033VoYXoWpO4hWQ2Ls2SonMyBL6LZC+8vTYpI42HTrmsm
pWniXeET3+SKMb3B4HDU/Fxynmm77FZxafbQS8F9CYdIswkQkuKY+HR2wlfdQVqZcyk/SzO734u5
zvK291zITWxl8EZuNbuzcuUPCSLScokyegJbPGjthFdvTyDd4p0QE52rhY6EBpfJEqbAW2TBWBaX
NlQFiwayfiRkIvGq/fc5djzz8TYBCFDGkov+skBcp1ZNNmpz/2COAaY9tLjI+iJC7ZDshrs+KkpV
gNs4mLyq19LpXs/vfop3XA6i45YjCcKSDBmD5ZeRJGk5SBCYOXf78P/WXP/Os83Bs60PNCp1nfMi
O3PljvmtbhqgTeApTQcJnGIoAjdW6dd2mJ62clBefmjdZ5vO94dVwGtYKdttwnrB0obcfLz4isHi
NBtLIXJBp+agKTrCLDYXzETq7q/T+L2YgNxbhxdRyc+l++GE8VAu9l6PD//9ao1BxJt0AlMGXna+
+pkA/4kx87PTVhRzp95nxEPtMOLwKQzmh7ZjK6+7Mz3j+mRpyzZIyr3CcDciogRHg+KgT0PBW5lQ
UMTeW4SRS0MK3dyFNDlm261r2LE1VqNbn8GfcDD4Yqg8M78SjRWCY0XawFe7gk0nUc/ay++6QMXR
K6lRdtH/rXbUKaR5cGiI/at1h9sAceNQyX8uYNCujMQmxPgb3+/lXZhqH/8LCa4xz2MGz3tDCv5p
ZOnuY65gWmSS8qgGsEd+x5dWCdN+owmCpMlA/G7W+flAamj1IYbutqpWDFqnyFcEGfGv8BmAYNoq
XRzKdH3v65TkaObPsmfzDTuYoBySVaUXu2bKCux7rvkDmmKnaE4cj9TjcJotWwQU5pofTHsTGDLI
pmrKnn5DQfbqMaNCkbaESA6KynP4NxOWIOoPmqjxfcy3TnUScg2IGjpYvJZmuMopilOks4+4690u
jI+/8fJjm06JU+hZhUtbzUp1UvSsnRtEd9BEJjiSfwDI4zcdP1sUI5eU8T8zQwUmfUPlGOTj76jY
Dd3u61xTU3W0E1AoA7nDbggiShDh0dCinPBdla9QIjXcpJZsDFJW2J9YvEsPBeLH5QSIY0IOrdGp
iPfXFU4g22A81Bjkrfubi9aFR2JJBjl86kWf0yTU1xo1ARYAUBc+pGOYPOT3zCUCFx75hUCeVrli
6w5mybisE0gtCeVp1pDfkjrLWZE9RNfZQBRqOiWRFORuyb1+4ZhcX1CfC5AcMQdxDt+O72Uj7x5Z
dg6XbxYSx0MXnS2s2dSS/TsZEX4Antj39JiuZwq9kvE6HEBGQj58uy4VeQJ6cR99l7j7t/CjqLoy
548mgraxWXMaNq1zquEwtPQZFViIP+WbVufFvNZ+62NzFEj09BSojsXPqh+dRahpXG5+bc2J8tJh
86O10qGCZjBLh4sTM8kntPortseV24RwQpqCFs6Sp1dgXPL8pg+KbRdNPIAEVEOIeDeUnbMGFwqP
3yayogvq6dl4tPk0IWRdRARWM/3LbmXI3f5hVdN0aMjnXQxydWfJMMj/BFrYEZevUQ/hoGw91nX8
Qls6eQUBnR764wW2XiwU6wTHJOKGdWmCb0CocuEKgBFP3LtE2a6tjV182AhApsSLT+6/vHuT3/pn
CETNWpmwJrt0jW3dLpgw6iNCmEaCZwBcibCAgKz1rrzjMAnLbCCzfbYZ69SFix5zDSe1Oq0woxBa
xkXeWUgzgM+LyHto5hVnv6em7SJewwwNJEqbeNBrzK9jV8DI1xnUpYwRbS40Y5FI1OZtI6VNuzNh
ThAPsKjDPYqIpKKRcjgZYfmwZIMc4EMaUQH/V+xfyBSrFemFOKM9WdPQAObiYhAUu3mgsbSd4j4N
//heyZc3rjV9YcUeo+kyohYUvWl2rZrhOSGgDQlXxyMiKva8yOMTjcMQNnjSZmO21G4SBu2fpO3t
b1dbF2dSJPDoUuhRM05RQHLYUlGeHHovszqbtbNAwLE92JHeuvy/kUda+8Gq2OnxZ/KDwDcjjoZv
7vcEOg3zvlh5qBLCN8z1ViDjN5FJZ2mw0KRJgCdpxu1T4P7aJ8YCpPNJdxJV5ffBdGZXHuI8WemP
lRX2URHut62+PeA27WV8r+J42h1Ox2dz8pwClG8fMzxC0iOZCYDA9uVnC51++/enCpTT7+zINqvs
uc3ADE4issai/sKghFb3t4pwaOsfiGZY4KQgPEent8GsRqovDv0lA4Akh3gT5uW/yLX4xOuNu7UW
jjM120c527wAn7ACM6sbz2tcWifcm06DT+I7IIAzHisYKzJPUqcUQGTE658uVEZDWoUi8+dKI53b
3HhuHdBSk+xE8Qfq/E67NpU48KEN5KcGRCS6wU/3Ma3rGNxRTS+jGqdDtxOiSU0f9XpDf8IuLVoz
Y5OuAU8nnrpnGqG28dK+iEvsmpa37e+C6qLdTyvJ509R/bPOSo+MJhDP7jxa3jGnPrzQTfRnL6TL
5xRjXqYum8gAhwvqga0sAWrvFEEnr6UMCciVCDRM5AC7CQP69KoSv48gQrp4+IEhsgq61RhSUfQE
tRj4s+aFOUovmIFrNOSjyJzDhNbBBIc7LsdR20RGJrRulPVpkCDrm64eW1g5mjJIJ7/5plwvq3lX
9O72nRlz4PfeV0XiBce1H7FfTyzKvDGgSCl7naRgkkG6H/5i7IfnipeIvqN+bzoSC1ThHY5ofGbV
HGbN/t7yJnkSnCeIcf1e3O/2RtD80azj6thmyHrdHBHWM2vbF3edWw3QWnsPn99nFKA/vvbgSXKr
JeIzhZcIOuPwHjWadIjp64F+NvlGehqyGA0uzRjnqQPLrc+kiir890kWuv354fvIZNtFuSiv9YAl
CrNKJILGnT2qpsDIfUC2992Xo6YwdUGfNehWasYKUfxBx1YeLpkgsX3Sa6xXmSkxqdEbxGmVN+GH
OJWrDgpe1ypmNiAbZRXZ+4zHsstwDfXfbr1dhnPgWhtMn1fPd8gfYxYkXO9GChLu1rVSLViCFk21
IugdmAfmy9X0fJRvvnwiPWLpRhGPYfYRw6K5i7N2IvCZ5OG74H1th6zC+W/GFS1Mk9ZhxKdXT5XG
8+TQtvS9jTG/OGKlxRsZlKLcX3ExuUXQUkBSueg/r0v6fE9eHLxidiAxgWko/LBZFGrXCj6fXRzm
dIIZE0kkTWdfQrIv75en17GNzwK2NwaYx9TIGU12OpSPOlcOw8t3XhTfviDZ5uYWrBQHZaRu04N2
1BdqgC0vrjoxQfV7skcgOykP+0RKwm2pmmRUJ25cNiHLPPivb28p/jD7A8FYLNZrxljngbIeF1eo
zdgU536CbxjjySg9/LPhXRgjBZUyyyM/3QvTWIPbqWfj2eAfvA7V7yLURbF3JbR1kOak+fmeVDXP
WNws9dfyCcwfiyofno2+zvsTg7LqA4HZTeT7pp04uWrU4Z0aGcK3eJxBp/BvY9vJBZGLf1IVU4eG
tDi0+Ji2HIy4o2bjjb/viQqbTVDUNsJueRqvFQid6OpKWz16atCQMSA8BUk7taF2vdw6Mp//xKnc
ilSMvyth4MJDZBmZwBkzt1xMAVYl/MHyV8nxF6R5ykg2uV9kAl7u/5jPQArOlpCUW0qBSlClzgql
nD2nC3MZWX5wnYTojbQco4gxOOMnwxHN+ifhi5yqLgDUYx7AukL8SIJ0/kKKMBsgHO7O8mL0PyJN
1YBAwoZztHKo91sseo+7wTNxhROG5lT5mroxGf+gbr/QIzg+P7IWPyHD+tA3JMbvWg+0gvpDJl8W
n2iMgTt9hi2U/6azaoTLhqX5WTv+T6Qv1a4FlwrcvS0eQWyHlW4WJJROqpxB/f31BHDTu51QyljA
lE+yEbSxuvHNFIc05PvIHJUVCE/7f0GXfIF7pb8105QumXL9sRTX6o7Ay74ST8cR3HkUXZalf4IK
rDLKVhNM7eqjmfGQuHK9/Dr9GMZ/iPPu4Jmv30q23maa67dIoqvrioheVT236KPnMGRtAXnVLBcZ
WpRLhQvczPsCpUycXUjU56tvXGxU7wZDRnT+b/vtyPmZafYEYkWAuXfyIn26Fayb8Du7qAnv7izc
2tXa1mqp0i+91Mw7nAqmYXO7Poclm2KaDLoCrb/McJ3g49XOplkgpqDEpbky7Q+gYd+W1kLoeGtD
l08UoUdV4X8mny+vzwqMMrnOwGSGxvF0U9F762L4EGdephHRmbb6wf1CHoGEOoe8zF3V52S2zpJL
g2StoyzcwUSp0Ezty4ntnG4FVdzN0QmMavaqc7Lh62jIpFZnAOcqj4r4rgY7S9UV4PTpFdI8IN88
/tUmCH1xaAh5eF5rIbpqliYN+5e7vJiesyzo0Fk8uTKYbPFb7arUkZz+A6xCClR6cmAHUgk+Yua/
8vUpFAO9CVMDeAKo5SyiRmuj0I1gaUcKIePPwH1SenAQ46QD6tQkfJ/CFmvnYXiu7unOKxPHJ2L/
fmTRBhYccE2hd9T6ZyZMkn1VIHcA1EpTqWB5E8nK+Hk9hR9mYxP4l9rBEVzfY4RU9njlyKmaNNT0
IaGLT2zW6mF72t8V1WBvltX1jgf7Z1E9l4aORvLAzEH+xEY/Oo/MQgMwitDNL2w0NtK7/KZlNPp2
n1sdpQ1zYsMfVoraSoz3WqCPRsp7QLYGoFSyZs4GK9rL6NYhAHKXk/OeVnqtkUxdA6gMy0feMPL4
0mBxd/nwKmJ5Ia0bA7eJoBpFPQzlzw7Cdl+APIxpZTQHJCwCw6KzoxuaeU5wo6cFGtvVxf9fozJe
+crzmJbRcQzMKcHhHL6+G3K2J+/b0fyxKZovY9ZLsEdGcdI42GEAgKjIiGA15jnFgpuZN0qPNwlQ
/2tfx0mcUJqho6oGWw+glHJ4a0+AzwJ9nWBMbasSL/7tLvqDuPMb1bQJvrefjGXNRqyf7SvomzQx
RiDKE3UB4qDyazzXIVyJKdo/A0jrU+1qYOI03om/bqWR6Igrm0vgoHpESpld1QUCXfMqkktnD/5L
OyT4yjrWNTuFjCbsQScnwB8kZhbxpjuG9bB/xR3UhJwL3B/y0HuCxentbnzRsfyY/JJKqeUP0WYg
lz+N/K6S7eYuhdlgs8iN4sewhOIvdDh00EaR8EX+SyN4maPkbOH8PDo6nLvWJH5K7zbaKkIWruVY
BPo4/MQUGKcqrO+gdhzQiIJnQtxpvvPaGdK2wBEOrVy02CZtFTnf68M/trj8iBp5c82lMKratKsI
BEK+s8h00NIoz2I1eIqCK1KAjxCVa3aZQfnp2Pm/IlKAxWoTz3llFLJs0P1BA5h4Tb/dgIeb7Or6
GDU6P+x+1aMGXkRmueOHb0K5+9XIQRF92uBX1EQZKKb3Wqj5RSR4EZBrfZ2xsBxW1nELxb9NrEd6
cCxNn+KkQO5oBNnR1q5X1yZq5Y3cmG4tbiEPmRVDeq+F00EVf0jxD8gWSTjEftFtqfDWNMPdbxMh
VN9rDivUCmk60oql6Mncm1bplB08cAmyGR6e+QkDr/OEgip+WnjdknLGXUCJUgcfk5poH9PA7BDT
nRVg+lKazIP4PqhtbJf5A+jeOD7D1X24UbPOIbI6t1czCf1wv65aRzW7IwJWaeJw4sAlCB+acBQP
K2BNP1qSeH33grfG3ZWp1T3xU6TI8xpjgkP6awoqEyHbbn/jkqleYLzWlMVDWi1+ng46q2Udfsd4
ADzG5+s5ebQlimi4MFkbEiCMxC3qgdQQkqbj6sv9eTDyFzFme61VXx3XGPO2wcHAcBMVhgbuVDv3
hGhE3x5Zsd6o+x5FCajH9UxBUCD7uZkCBwwh/3IrSu7oJTLz83JtXRXPvCu9zAp1yAu81W+IT0KC
+30yUOdrQOepeFkFeX7vqRMjOhSgJUAf3M5T0KQ43Z115XL+F2StM1FQccKY0/kAXZA68fHvTwMB
vjTN9cJ2YmED2x20xSWzZ/cFzvl/l1zFf6l/SsmdKPeOwj3SkMIWUMNoGiqgg5qDvhJYEpO8pwSB
EveWkDeMQO9omItN4RrcFAKyuj9CThZosoX2pV98zHSF/X8z77u6SKAteUGiIlLsx0CbBOJQ85eP
OZdMg1LPDXbP3KV5qqBDtRf4l+OMczvuHWZRMmJ9KfKxu1WNUsRxdIQnKON0y3X3Ux7r4XuDZJc/
Gico29RP2rOEcXYQ478+Q6a5kG45A/2PW7rQ+fH50PqMp9MjkyiNeV2Xz4qUgroFcZf9hJiVJdQL
rl+Jk4lFPjGgM63WjZzw/nOXgkCbt+hEYBu7tNhrjwFnZCdhzrDYFCrC2cCVwTozgBFTw6Yuigj7
D8peXpMSBfT5/f7Awuikzbf8HNpfO/Zu+5hCi3+MdDAeP6K/lE70pDzKBjXdzLr7sb2k0Vw5hTUS
OdCFNV0DbIKVQ9C3cmQNCQ8H7+mu2Tse9Mqj/h14idNe/e3dWpXviEK+pqWqWDvneia+QXxEaz9m
rPmyO7Y1YMwoUiPoPu9CZ+lV1UGintbEPls4uu2Y0uHektxZ2jqOzsP/jzWt5fLVsxSaWdKEVUtD
0UDPZTo3w8jLqcoxFE0ZMiFqHCvRSH7ekQpE5NVwW+Livq5m/KsLSVA8mMwc4OE4qsNMF9SNjAVl
vswrHE1k5tu+8fTBC5wERXJAD60yq+uh3ftlUc9pJ4pnUpRAv6vm+06IYG8AxnQn1AVXg+F26Umv
NQvJFU8ztx9vSrL4C/V6jmZG1wn4LtBMCSKKDkUTstseKgu0q+fZZVEWMuACOIPcv3lAkGTy1bGr
7xhi6EHQwZfdQm0jn1YzRXl+xfPhd5x7F4oLjiudkO3AZa+B8M9eo68tGbKWDM1gKH9bKo4SOKX9
h0GWrmC601MXV9Q1AfvVapernjNGO3eGb2wldVPkElZZxwzUUzgOXfIYjK0EQ8fFnwGHdFtX4REy
sRmuWmEmhqMKY/ew60d5XkMoSmxCbrIOW5MNqRdi1GQzal4GQKtL4OatRKR/Oq/RNIAbhHWHrp6/
Pi4MrAcL4EwD+2lHl48pmKVPaXwh056D36pJvqzmwOfEr7Fn+NVT3p9GOXzVjOfLo5TtPbdN/fwB
qSvrMK87CNBINdivDKBXfW/1zymCWC1QdMeLB8t+RnLPYwsJMPkwEyOou8ttyZZBa4bgV5llWj9v
GMB/BXiu66mz3x03oBsy3OpG0MULShPuKeLCDRETkR2jrHExZeiECLim6+dET8Haam9M5MZFJkWr
povIJ2LWyK+P1LrTuhAajOaNyKx9I7R+8qqVdlNNON0Llufl1yQM2UYc8fIILFyd2vbd+gfGU2zY
4U5r7H5YN47TnhszR3h7eeCRGrJVderXZuPRdhtN36TakowY0mW7xQ1Ly1BqFgZgcxm1e586Pfzf
VSX14mJegi9YCJ1x4/VvptSMhOH713egFyh/nLnLsgsuzSFDNBvybLoZnK0ybD5F2N8g1cwaScod
PV9H2b4bdYxR41vHQD2KkD3fMwNiAVwXpiMTqJ+WqRvJL24C9h+pTHx0TtqDlimtKHzD7S/D/lPl
nle0giE8CgJAlYTUA8uWywV1FzhHIldLtuZxM13BrLq4EmN2Z54/ZnlVonDsEbySF6ME49K60C6e
UD/rds7JUAbTAL8Q6+PQq/lPKITArE7Bh1jBk90x8dvJn39uaB6g/aViWzIieFfjHwOGfHqxVJQ8
3i1FB5DSlfHR0wDhg8XenWBn7ASwjGHrEYL7LiLF1He5IqM8xXm+VYOxG40TJd8QCJXqcn3W03EC
4JbF3oAeY2TFud+ZAqQCoPX4+kPvCfHuG1QpEBloVfIUcc1Jdfa0+LDZisPQKGsI3NCRSED9cds8
zLzWODJkDMLni0ZqDyLS3T9YB9pL9+GS5pa83mPM8bN0D7sqN8tCsQlOnKj8BK++nXSa5vNMj3sw
SZcmBRbCPFhO3dw9HaepnuRjtFj3pJUBMegblu0Fz78tL76H3+1pkak/vTKOu3+RNlIB+EsEjTpy
/NXolf2EKLG3arHbSUDC9T+whpFHxVa1Xhh3XKP+vi/pBDYYOdqgIgFdwiZdyqzuHrO1w9/WAhfg
UBQNqsjSvbLW2hioqMLt7RrfHOmpcCeFT8DxUgL8grJVEAoda93tqCRFfPV4XVtkuGcbyvJCsraJ
H2DEP8x/IQgU1vNl1R9jn8zlW6GgcJS2Tk1FZzL/n2RiQAWI+dBmmDCA6r3bzins6XOnBmoHgzD4
WPE8sQrJsvzBennkezV9SeibZpzvBbMWjRa74NvAF0lH2gpkXkOgVazQMfvK6hNHf0yH1d/1Ebxy
wqICUp28mQQrlEvgGyfFlNsbuo9Cx3JXreAkV2oOiGwb4QPxte98gRNwIiUXxbtSW/Avh1VLBprH
2oAs3RL4lN8l3HotuCNnFHWOzJMxEdJil1xEGqx6Hmin1/vi5nBPIsSvXQQY2YEXWCUEntGWWpr0
0Q+OkqrmmlS+1aey2Ts8EMpGUg8h8+rezzdhYR7aDQmLjQkrrHx85lt0FmDmZyMq1a+vBli34La0
qjXcwEN9aMMbs9TSTeW+cghjykZMIEx7dJ+QTFY/jgM1Qmx1puUVuPEWx0m5boUodG1kF9mY+7PQ
0XMmHNag+rJ3EDGReq0PKjs7QT3NxFeyn9uG8Lac9qpWaX06+wNZ1Yuef6ePn+sE0AX/VFiIGiw1
OB6tPNVhxwbGemV0LxFgZG7JubCmNLQC/GM2eUsHnlI06baxjIK5Ckw7Jeg8Hxxk/voQT4plwwao
lMoIcENkt8SuRppj4oZ/urJscDdLSyO3SUisqLIJ7pjf57bnNs/V12B+Bdv4SiagZu5Lc67d34TQ
NziFgH3wdm3VRsQzdtBmbcPYjoQL9w3nn9pd8rPPP7l6Ghks+zYnFZzuyHuSKktENuGF8Fqav2x9
16LvbhvkeV9lMD8P+VNUUrmNwhO/O6oLksYnhRE2KUfWculUq8ueJDwXMyqg1tDZPRYNPc6Rq5/N
hkkIBY3VwvCONITv72mBHDeHCmLGEEPqSNkQ9MfCbNlLF8yeL+ZBF3TFheVIHH6azPEdiGmbtixT
n1NTgBXK7hPMsU+1XtiI3ILlsDJc0+veSku7vAWyfKvCiq4YfGpWzpdjf+IosEc0IY577YlzB8r9
alg6Pa5zIs9UzQfUe2IN/0v0taKF/7uW003D9RSRZkiHIaEM7dXr7zyn+GGcS3naLKGSG54FvqkZ
Pw+eGZGFDRkGdF001z5LuyRi8BNRTMxeotGtYeOhX5g3+iABQCqPmmg14VjmuHbMuVNowmYdon31
YWRPDgP6iztpN0H+TklpZZ4dKvhjjt5t0E2FSs3ieGgrgBefgPVGdzj218hAivQeMvGxv2b5ar2N
GPbEJJc9lUH0WYz+b1zFMX+lXGSQc4+ZYEeuxnMx6+OjcPjciGDghadRCQR7O0Ac5E5F72OJcXk5
BnW0oPJ+amNNh9lkooU1ipvBZ1OSJ9V4K06P+ApqFjYpq2JlJO7auY0hJ3JbPEiVR2N8NJUP38gS
AjDhYzMipx/YfOb1AnaAIxBd2NS7c0dUgRm1kiJ4bhroQ+UCaCX1+90pvy5oQOt/R+4XmvrXeZuL
Mb3+ALFyhI5Sbv9SotUO92mwzouZVF4DQwmfusaWy10GOhSDv3mktNVj4bOyxaUV0ZOy0TMarYkE
+e3QU5scnJN6GHkL4Ke5/2GptCSGzETxVyRFjNaL3oD9D/L0NqQB63eMOVu3T6QU9A3jNwWLKl8g
xdeuastkybPFNp+UAzZDlhnJAgbwJyX9FN5WKsS71KM0kfQXmH8XJWu604hmTanzGip0Ec5O7LOY
ckHiCI0AeawBVaZYHQIRJeYvsDueVP4h+KLk3z4smaOOxN/uGvbbk4wzaq8aWQkKOIoOM7XFGO8q
5scWeIRYM0jFAK+g2iN1cUfHO0QvkGJb5ZhOUr/vQ28gRuOp93C7wwUiME6KgOpcwUmwy+kjkkvp
g1RAcWCMkW5Cjyxl1gxdLrXOdb1kMzfqNyJ1LwFTAmZ7ilX87yDmOt0YWVCIdRxISUmlfFEFYtNp
g5JOrQcVTH6uyII04CHS8eh5nlOSgnNnEvsh0Hm+PFhXYK7ppvzCxLli904gknD6MzkmcgYAEeOX
EZcQuYLbTiZ/Uz+22fbIsJBJmFg7QSum1Z0MpCPzmXIIB2S4zdd+awKrIIHtMmgvWq8DN6dNZees
nRpLlimwOiU7wjKyaVEezQ78Sp4HaW0Dl2V1Jf32I02zdxfa5OJPwCeUlKftWReLlEvGtM+jjI8B
1zcVfd7KdebB+bS4DD0ZSHrykmTagbUn5t7Pgafns2DJeXskKmhLJH1Z3j00NEZMXSYv59pn6FkW
Ccp68MPGVWpvOcubEc00DkTipNwkoWazO+ARaXcpnqaed1g1L4fMY72L6i2OeHorYznojBFig6wQ
dal/VWKWcShVz1iEJy/0ZvFINRx1aRLzRtq+xOTp5eEeEavhOkWvba4VXEl8d3JktoSB3YKH72hw
vSEBVIChT+iC1N3r/h3bZ00teZbSpUymOmOhoj1CIsCuP7r1gpZ5ZQnWSu3pDOGIgPAzSrcmLxBm
h0ctIGl16xU3dPlpMpR7k/LLhB2MjJay145rfQ+DcmJzJoyyOvQYbUIhA4vT4QeV67zE9Deabp02
D3KfS6sl+i3kwFEIA3bCdUustE5UlIChHzWvUFactQr+kzksJ8ydaQLZj1idGBkC3K0M0xUfhUNr
TxCXue3cNtxc0aBT2XFl/HYNrTJUyHkez9KjpVTr1kZ9AwoAz52tny/Dsne3lhrJrxs7/lhryx46
AB5bGJsLx6QitxhKVbuI3NepVu5ddXS5C2eRKuKvP/t6auoqadX8xyx19sQ0IzGDgZSdrIBro57k
j19nBPAD72kRQwkMjLE3wXGvh+ImrmjnIMjVZoxpf+IpWvM+Y0k9EzNjbpc7TU3hEZ/aFgwE4a/d
fXVNCAxxecPWwZ4EQ6sGY5eZ0IuKdTucWg/Qngp6rI6oDCSunmp83Wo32RiuFEHt9ia2rIAfc8ME
1I+uJ2/0OsnNJJ9hd6TWR0GuCMbpNxzZv4v1qLL2L573FGyrmu5qBkrABP05JhFVFtVj5kgg8oj6
cNl3kcU4ETU2GfVAI46LsMMqhGNRDJiZhCzMEab/NL5Q/U4uviod/RWlj1htQ+QaCSl3cOINgd58
no8wYEZGY7aUaBrnhzV+QR8POOar9UHazRHs9XEcErxyykbrxWPDcN0T1I17Hppl8PGbDCjL42wM
85j25CKzUu76apCn0rERys97EZOq35kAu8tJRLZ2lZj70ogH73OihJ3zERQUTQiiy5Af6mKzCp4N
qYedg3gKEw2EM2EgnEt+RIcE4dWoMLvzaC33/bwA4jsS3xec1cjJc5su04aXzZDDq0rk3rwGD+Bp
OnTX+j1JCp/g+eqQNOF6DMHRH7fNom/OdvOrGsFcrIMaLMrmalAZuQhZY+AxnB532rImyWQ/7HOr
43cBlpQmovVu1Cv/9ghnJk4lTRSdaqA9y+SD17rm3400Jiu3BfoHGxCci3jcHFoE5mbvO1fSwRnh
nI9Ha3qTiatB53wBgiLSzkdyMM2tjkmbnA5qnlBpmxO4bK5nJjchfIF3h14aCfonxtUaDWVSM6Dw
yY5fow4lJX48aj0mpNnn2xJ1PZcwy6mQeq8shBUxawTs5/H6DwyoUeJgCewbrzXBrLLFCE8fA/dl
jmdzKf5umBMbDatWpTRpmcojBce1I9XflIl2X4DzXjyUDU1gIb8oPRsx/rQjQVDHwDD/erdn/bK6
XvFs/0eCE+mrGrMYvb0P9cWq/vkHgrbUfUIENBwqGUSVxX/lCmSxWaraFc2BjxtIrX6oBsVqWMRb
tqBYw8JKPxNpi9YS5VOB9kUjgL0DczAGnPTEIfwECtxVVb8ZRDpNtO5bXe39WhZwyEbs3amGKr0L
rLuDRMjj537Rk/74QrIprNWfXHegS+xeMlG/hDKJzXCzcrvEJxN9ssvhAZgWRjZ3Grd/wfTxnKmm
ZzfC1WUKo1+0AP0uGB9oj4LOp10V/AKi+6KJX1BRgU0RL3b1EkJrML7632Zg9tQePKjenBcFRqV9
lMX7QZc9GBWrkmGUiFYVIhW3vZtDmihTgaFs7VMWod7on0qeJ0FjehWFuzJbWksUTfP1U39B+iiE
R9trFTKrlXFqkd1aRAQ8BOoqxcS/aC5eLvxQ1lBoaQ1GWkjr+vKFhEnBy/67Rxqgasr2Yucspx2d
qqGq6SuDx0xjeT5WQZBEdXQ+5cTlwZyHpolj4gcrcimmSg42wgwqEehh61s3nhtK47oqTwFfV/gs
F4Qo0wL2VAM4LuIXZbJ+uTVfY1B9BTctSvFN+/DT2GMtmYQCdXRpSvsr7rDcd0LSHFx2DUQNfzRn
lXDesuzisB2mLvJeh/4sg0UkkpYpCCuo0YksDoFxEZuob878w6odXx/ZfzLnDFvRexz0RI0DRFyK
1ZkOaVLITMPrxO8CJkeKktaZEwqyJxy+JSYZRcQ2V8KyAEGmvjDxQcp9PVJeb2UkBb1yHU8sSt9T
09j61Ez2gtznzUWJaB58/LUbnOlk9olr7nTznLqZXjKFC3hY3JRT+/4ZL02bpGS2r/9UZE5YpsMw
xOkWjmhCq11+tz0Gyizkyr9cjUzTtFX/8vjWX7EcfdrV7THOglPjwLrsEnJYaigBaU7TgGjrGiep
Hk/tDTkx+T26Xhy3eGdEx8+D+GUD2l34/jPfbLQdFgd3vRuVpf1CwIpPOd2/arlQdYSlL0kA3lSV
cPLaRnq87UT3BVFdgN+ylJAIgEsvyd3IUQv7qzyM6y2KoAOV0TucJ4J3FIUBM41A9UsHXX72jlmu
Cmoc0j4i+mpfKanqAcFnVcg8RczwKuQ6dXDlLTs7VtQ2EEb5EhxPONxvlLpwdGiJ1+tC79UCbcuV
/i80dYybzHOjHUlqoNplCK3nbyTYFQhdLPRY0FLcaJE9Qj8zpamjlDHkeS2NWdgAidzvAZ80qrmo
Hkno6THtT/EhLBOd82+3LEI69e/12xm5Wn/5hj6O52T+u5ECYnZGxrdM7c2/2oaxi8McIK4cv4sY
UdxdyUStu50EROngZ4RTfR7Ox39S3rqVV4ITHrO0KDvs9GKP/qK+2iLSUveUgkdESvljITjU7FMF
Rpo9Ma4midi8u4FQjqNpFnk+0JMfadQwIk2IrEdCM++2aKjCXZWJ5ejvVGKqLYWdcMlxq6LG17Ps
7DtOTkTTPFNWXtqdWkVsVytcXoHh1mGe1FQ/GyN83NWgb93xm0Qoh/M0CKAexjlqK2s5CP/IbHpA
D4l3uW3GL7gj7xvi8g43vEctSL+8Xpd0NNPXPU7I6nnKTH2ex+WC6H5zvw8dkl2QUhPfj+/1M05W
CBBu4Y4RtvJnNIRXUsXIXE+x/rOLV9yRICJkTHXvHbSSNrNDVl4cR9umgTScn6vPosXO+cCfQR9h
SIPC9Hje86qcrnhtzknnXPsyk3mHSTRsUuL1FO+Q2XmO+LtlOE0rwa91QGw9Ne6aJK9vZO4LJkLI
AZmZgURXuD6fym3c1qtV0fCNOR0K78OyplS/58laa5pDg323YuclfZIHTIyV4+fUBFsZcCiujWx/
CAJytk2RslN+y1kNQnVhfBZZhnVx+4i9jGE3Ox3TzQIFrlLMXyQoClYjO3ZnQUKcpaY1FMj/LnWx
tBtqUoSaTYFGVMUTMzDwWX356vfrQCMyH/W0BvEy7yCgOEknoVweSiyGFO+qJp5gNSbN07lnhDXD
/gsWarEPykOR5GSnGLH4Gk7QSZmFpxiE9E+23WzzK0XTzaibkjzZHoZx+TOS3i5HTwjaT4lVy+HL
fE4bdRtgALCs/QDWkvngMsa16JkGwZfgIvx/xBUjT+T0WlFzgIQ/xoeoIGRITVjfWMI9gcPrConq
gzJNT6OxkyIYhMGSPweKw6sgfN2sI1KMC/vpHSKqVB+eDiFiU9OaJB/6NXhNV9WPb4oJ19Y2xv/f
+1nXeL0lxyfGSWViAmVEYHUZihWpmSxjnHB4hrjNjienVIQ6/yiX1igvzo/F3/xDxtf7tAd0BW0t
1JnxqkAVrIljZI0IdfG88cGzvtviyAiUNfCMDHmldXJgMGQZLUUAHxcDzHBHI6eNyO/9m9gRVX5Z
XjHXK53hPwxr7LKGvsSw4EGSRuE4qIxZwmDTuSbvDlWBVRbF+M442y70gSvO27JTsXuBaO2wPVnO
B/6XkRcprM3shZkmNq9hUoCmk+/qrLh6S1PGmGxNR/jAmdOtx/JBYXrcwOVXR2f5/TytQBLmWX0e
uMrKOLRRnRnA81hNZupsouhh3ONW2rSwT0jHjj8nhNi3hrhWBsSIh9XHpjyuVgN6rNKg4x/+wEUg
wbBJ3oPuC7jH0l+6nvy/0+dpsGfg4ue2gy2hxPTmVuVFhgN7asnrYWi3LgHx/lGR/ioaEkfaGYTd
K9aNVTmH69Vdc2zo3m8PVjYhu4AMLBqgr6RDSSmFtVSygGi3kRedC6h72TuselHLYwv57BSz/TWT
O3nkB89BCOtLX/FvoEcTAzGON5rYbqXlzhwQu9CraJMV0UKuBj80KZqIWZOZSkFXX61uNHdr+3KV
EbIl8DFDGWh/MJ59C2nqoXppiD6FaYuPGv1GGSLxNZJdsuZ0lLNmqOpWwkk0b5pYUOW7UT/P0jD5
TPejPIrOMjV/bdiLi1quOPWki/N8sPBmm3Ut/xR4RVHyhrxW5JdNstlmwhYBjxSruRNB+EoLkvXm
MqXUZg/YLXKTA8IQ3UMZOaBH0N0iEVKwncex/xLivqM1B5hTHVpNDwut8bMXQgoMtFs1h72lKHdT
qw0RNveNTtKgZtQriECRxUmkmx+uCFNI29FSsWyOCfnKjB2u9w3Avqc6gAPlFjafATnakEEE62MK
aWUaGrfaDXwMdNs37txXHadNqUcaba/0kg726gZn5VI1PCWiIqu3IkV4RQ3QkvGegmmn/y1Q7C0d
V+LxJ/g6g9z3EwYSqVugztSVWXzw1I1UKpQ9jM1K0kf5ieUHQmUbEZZWxqourQcSsF2wfatQmceh
4rlkARvmaam+EHpyIB1/Y+4Wjuezhccy26X2rEJCgK6Vy7tAfjrzAbvOb6q6K2mxKInO7hvFvvGf
4Jf40fMt8oRYKL/BRhvfkD96MEj5VkNirzQ/l+Tv5AUAJxUEhtka4PP+0am99u/fpKQXZuqsYzNU
/iJ1N+ojc2F7tmDsu2awo/pCNsCBKvkakKVkHLpFmcmbz6ueFEf4Tkro1Svuv1IbdBX8o0bIihFX
DoolUiZNWyy1/n7Oyn3mFqj1pVKiFCRNifNKOfGiLDCPDQPuHbsRwuI/xzYNsRL45NGCX5kaFOId
L2q7sCzyhNdibom8FO2TyMp/NTwr4LpKJfmncW8+hyvItVUWnqi2SHf3BYXr0EKjkZkYQBsHqOV2
E6EPgA1NBXWmQcDeGWX2N/zRx1lVx6PlwkKGmThqKmb6G2EMfDmt0P23FYq/GzoIELXQ2pRQKZUp
zuJ0cAH5iLiuNggLHhiHeNA+lI+KyYLDrYKDa8Krwo0ZcuEyT0vwoPLbaNmUx1SijHE7kIKbyo/2
/yUBoaESnHHUOvmkSxBSfFR5RS2JnB8Ph9AcJiy6G01PX5gpLoktk1EfxXqUee1o5/0bZetSM5Q9
zs0eZ+35QLJADEuPwAewfCAzhNyh+ZO2pV9UYo0fNNvDtO3fzwMlh3wWsB7Noo/01+WLFFZ1OQmp
lCYX51G6QAgtdHCKfEtYCNMo/Pbj15rBp2viezEjEXZDloaLJD+EjpelgfzjI7fKOO3iDIyYq8Qg
t/8q3bAA06P5AkV3bI3Xu26DvC2yelYxUxPa/ohrrpJw1ZntxdrPC/Tx0AQ6Zfm0i0+AtRm72nyj
PFoXWQ/ZLbAWbNe1A5mb5yEDCniWpAMdxDMmR8qwclGGF3S+MhDEMFBHn9d9JW3EdRI6jLoGvOkd
n1VDbYD4AhytzbtrekbPCeaIgi2yD/hYBwvixX9MxR3OIZNx1rSyP5edhDIC9JbFm2YgG59p4KLC
VEQn98uI7Ylsr8d354W7cvaXg8PGo6atWqFLyn/aVBeU4IbQFXZzeoMUCD666Ron5Ie7RUgkbdf8
wQYl8HdupbtVzxjZuAsIqZYvZ8T+oFdCJO0+P314vNq8LjabUmsYcwYwzM73CyGFyDpA1B3GopCr
62sLpYF9kcgDvO5pguUg6yiaGIa+I9hOlE31N9eihm4IA8QCoX/HihoIbOvJyrlF8B/r7ScjWSVB
gtyjMBWNSWRQ+XYeoCwR3jSsDqkGaGGyMHdC9QCZzwnavo5Wn9GhqaKRcdxhCHpw6AFXNEBiW4AZ
DuxJSSuaJxfYduob8sYYR/1jxNhKDo3PRRZtJg6wT3wy4T8vtNhCI/6ZH4aekS1w5gFQUo/umyMU
kafezW7GZYn4z4FaQQt3UdW6/TJ62pgC9bcMtqBoyE3WB9GWNXW43oE2L3J8p/QFwpjnhLxjH/G1
TNsg2syJ2olrOZsFbDxaraHV+MKpEPZYUMxnJV6nYTe9earNmzfgxHfDBpeJhDIHhZRv6S6EV1qx
78/S25R9LO81aixnk9B07IoEjZOw7bZ9pLKFJ7+rTJeBkUysEoch8UJxWYqxhZ0OIad2q/k+efiP
EXLzMSuz3Fi/AFKimd1ZcTyHntGccriscEDXtJ+grfTE02DKfhUW12FRYYbpI3tEdl0lQ3QDNqUP
5uleA+hfj9AL1aecah7p3SgtZ3rSYEx2to7VbioGCsp/qsDONlxnN6cpzFW27sdzZ3UsSo3/RPDt
SOWgNWacnq/4AgLwfMMIN4K4qSm5H3D8FL4+AOK/somNNn+KTyuuOwx1Pm4Feuw8F2fN/0P2LPfR
nFdhUkZZvb+xSlkeFF9jAr36xyPVFcgz0qqazMPG3pxDgOhLnvyTEI+YhpNSom6D/gSeN6sD9AgC
npBR387KkwSTQVJPyrOZo8UH+yXnyBAkrkXcgLPhKJlE5jejv4Qwk4p47ZfNm4DavTuJOltM2eIU
N5Kge8sAgMJDjQI6HMIOlcYFnAUwOUjGjMINdxgZROiHex6Ueh2Ftimd5cU3nVa3x6RX4nDc8f2s
phhqVhl2l3a37WhmHtTdW6W2hCmXfKGOpHCkvMTZisOg6K3FrPNg2eGRWhpIqovQYuK8ZHWVLkU7
BihZRbIeJe/c+dgaQX1dVeBu/5hzs1R4RT+gYJhw1lJMmowoPccPScLdqxVKhJcKrwvWpK4zzZDR
MqCPLvl6svoJ3TczQ4qN4e/VAD150H0iSoCvOt0GouEU/CVDolnyZLatC5v8y/1jT8DOH5oQcbXL
41LwoJ8G3h6c6ftQUcO9avHOkRx+h0rEk0kbU6VXFmD4Oz1s4/DdoxUA7cfGulEOZyPVNXxL2zLG
1qedLR12M57hqhbLrL/kUZ1IN9dbdXJqnYA3NJpoBYWKpTYPvbvMHPZYNbjHtuMn+U4kLKhNybJe
WvHgOJncIlPKj8VYJJYdMTRJQMRClD2UEDlx/TW5Y9edJnx6ti98kgmZD4CDH1+1iTJCoBM1Djac
HHLfe+M5BkxSORTvtXM80QcLmLN/s8MKBBrE3tzwlhXN6cbTjA8xun6RZww/kBiDSOS4qJq0A7XI
xvWbsBmNKOi9FLRrMjAszE7OW8TdF273LU4aFvCB6vzHBtg4DGyylceRwnqCTpmtny7O+BRFU/Ra
dgYbLvxoFe2qZ70z5lQTaxqkotLZ7O5PgZrg4KSi63Mi2zhRoGMj4gId0pFeHadflckMEosLOcX+
vr0Ad7KwAFgNlLfC02+d/3/Em9jZj4DaU+FnVdvjZOYRwU2LpVHrUUZ/wVNvR8V5IPpRUVMQA563
1fYPTAhkRvdd0YSz0UQ293cUoEqCtvI5ieNw39AEi2ePDK7E2zib0urIM4yeDRxDxt9FaUqqfGq4
D3DnPAThDgxaandAFH0TCyT7Q2yrJFdGbgowtwwt6AYtMsUWXnwjhMAobWz6lGYaQnEN2KjJy/sq
OJT5LQfuNTsEsaN++fPdnWC7hnv8MM12NJX0kfNejlHVACMB9g9+BkBJqhu5vyzOn2QlIf1GYVwZ
yE3wC9R9NfAjwFCtsNRsaF/Iing7xN9a/ShRawtHbOkBlgzV1+8phyasbaISko/2AdFshnBCtMkt
h8mqBUNfO1OD3Y6GUOb1bUGH4HitLC9E4w7D6spSTlNg4F0uaZYAHCG0cBZ71l0RBt+JkGtYXofC
H/X72Xnk2TpntUy66h1hLhVpawyq1RZmhRtUmTMW4s3/m7a9pIvXx0DtTrroJdCsyYFKL59DJMCt
nyMgPAhJ2efYN0o0d7BCv6+eXuYb6YFl6I8ulZFEz698hDLGJ2o/44YeRq9AYJV14JIKZ57oKJli
mR2KkDXOrU+xt37mfWFnWX0IUbKoOIxswRceadn0G6w5KBptxnrl/rz/LsecoFgGcEUO+U9rez8K
L87Vt9CDHalzvdIvDkIUDH8Z6bmVoDS26G7diZh95R+geybV2ADAtLGGpIZzhh/VZUNoo6HQ9OAf
6DukO7F2kbbQULvjudjEuCzqxD2jew7A7DheCp+0Z2aOYkNY7NJRhyFTIUT6HtR2jThmk4Obs1Uz
ydRDdkpY40zjOLQCEX81j9rgxKxHhT/wsUVOlerMj/mCc/RdvePQZwRvQHAKUwAX10IoTHNQnbOF
9RFDpdIdTtx8sJ8aUGfwUWWkNieuNDuhRZ4zyaRsVe2Ef/xnRssEu5D2OVu0++GU6+IbGtmWhN/h
kIuRipzcR+B+QrxI8MfkiYMTR28tejHz1LB8sR+7RYY+/R2Z262jIcjw4VaAzJaaqwb37aWvDfrM
WuN0BVFasbMiTsQwvoeLUrqOsHAF2MLAjcuppCkOYDhvnAlmu9hobWHQaxI6aLrO5ERYaswLXudJ
byZTK+RvJapenVqzqpAj46gOv4Mn+syRsqLKJEzxPn/n8T1mtoHmcMo/on01D+36WMe1ZtEM9phZ
neThS4G/vvPQ5QTu3wZlkU79n+uALoVK0tdjyLF+8BcfcROzjvg3+kbonQFQ3hUyB49BG+97f2Xg
unEETwEtYSN5LD8q8g6n/zyTATvUdBbrlm5IcQ7SI3QNtuFqvLhkSjMgu002yGgIgMVIxLMPb7Xn
RYbhuqt4QDvNmTH6mg72v2b0S/g2FjnMU8ZRpxJhvrDTD4qMlBPmShAX7I8Y3avwYwgACJPX/nmr
OuvX7HUcByWgtayxHT40K7FXC8SSDTSluqCWH1SghlVQqfXFoCDxKJSRHnZyTNq6/Mgp8GMSsNK3
SGRy+Y7RD2beYqavy2bMXQQj+gTEH3N66pf2nNLEia3XZdokzfg3RtikdBbydn6l+0N26+3ZPlzb
1mWQo4dQ3cSn/B2TlvO/HotrpbCjjotiSl4vU3IJlymFXjtDpZM7uYoXYRAhJBDvuH/9/XJVf0D0
cUJCPjMtwXFQVySHcfCmKcij8tAaagEoOmg6mf6ASq+QZWLfwUcB/z1XIZV8VbhYB+NZjBRowh3K
zXO4hsFi+aWZWyN5i5YJ0R5JUo1B+98+LTkLQ6TBETcC4sukRsRsyZyf31qqe5LUFXt+BCBQSjHL
QMcNxxmS4ribFTvw5D/RpFGHVqDqslMHHe2DcXvnW3GrgOwteMYZTXmfz7GM/QloEHH0mQnxlGFX
dwYEocVHT7jY0UgozqaJswh9Fm/N5n9GLPutwqBcmBZjJzw7cwUTj3SY6bPh9O/dQvBHMG0F7yvM
Mi4cVpC3qh7ENHqEtqLkp584D2JUYQHuQC728FBfiizVIwgn0XH5DOxvlq5GsTJAxGlwjM0Yk9Xf
yfRi7Ehqs1h+i0EBB20GlPNSpOUVetmNZ4NsiI9p0reM2L91mULvE1kgglx38h4LtBKp0jZmfxNA
M7bPENuDB5uoOAj0ii1rBryNlS6EheZne3grfy3YWncS3xBbcx+p372FZuTRoDX+Nj4jJFiL9V6I
D15miIElbugrC6L5rZti9kTQeLfs+o/VxseWU/3/4N6KcEVMJEIK9oxdiWEM9dz8JiazJ/VjaSjb
19YdwtdLDdXkfxFAQDDzqETqs5xOIuGdkZKGjT0ptPOzVXRc1TPG4EMyGxavyAB3CzXn2wlBv0cr
SVptijO0JlbFWSgS0j4lVJlIiklPP2kRzDNh9E8JWXN2QJwQYNZBeKd6Au72wRxvhK3d5Vsp4DZK
k289ZsESA1GGN2ulu/tRkWBtvndpH0TQtAvrkhhQcbeYMFQ5JaKozHPMqV2EWlUzjIG1zs2OYpBe
a9O4qbPwY6GXn6MhsYq8xzwDwLF12M1lffZBnQy5nmW8SMu1+IGKK+GtnDUpLcmbRVsOSZPd8Ro0
NCHmXYaEw874M9p7sYIsTM+1f7Yp6CQEB6vaDgRC7sJ7FLFcB7ULF1y7bL+QXeLL86AeZRrnLoCn
xz9r5t2k65i9ijd7LyB+7rCWEKGte5oX592xhXATjjEviAm1FoRUyzFYPhjx4QqHR1OyICZShaZE
Jp/kYtcV++jhVtk7LELTFOUPOFjv1kgOvKY8CqZRROPBF5nse4QlZGqtNhXGqxZstAfl79ZxOCU8
HkcGyu1O/KU0WN2YP+lujoRDfuHszoVWacbcJs2ikM9hGcdIr31axICarhEjiv9oIB7esmLAT6vv
/msNO4nC5HH4UpmE3moKDC+Tt2LtSgzKWCLcMGURfbVwRGn2Jh2jddmOVz4S+PONRmGIHWEYys2L
ABaCnKwuLs7AG4Hp0mK1NWDK7NR3W/nJh8xRhscK3IbmzckIFxnpeaw7vmzd+u3CkBE6ijtGkpDN
vuVzUeq5drOi+Rat7Xh5Hl7dDvx7NnKDjk04dpgKLlwoJDbKQ8jMKbVj69wVQiqYyHvp/w7hw23v
OJPJs2EOq0nR0tkx2w6UuALDcuMV+Ejh7Q/sJUSqlnEr8g0tytFvwdyqJg2an/JSvuXwRlNkTynu
wXO8nzS9FeSCi0hGtjtRS3GFao9vnkZWf/vWsS4aR3tGbyauGMlNUlUP35JNbSXH1ufQaBl0TO4y
i/z84F5F1hGHoYEaWHoBgPXNlIUSQuq5bFtDM7Tx2b/Se7VRzT5xI514aes26WTi2GcK5Rnaupla
cE/Pv1lJqXq17S15QGC8fiFqyK2Uno82+zgVfbiQQRsOGObZbQvmQEdmYRV0Fx50ag+Zdyzgmwvq
t6GeSORW0/iJc4gebJQfEgTi9NyfZJJuZJzGflbPYUqCkFaEymUvywcHuaGmQw4YpTq+nhgihaFz
9CaCeqtJK7HgOiSeSeTVUeN9jDs/5M8OtKygDWBl/46oLT1Rqb6JJKuyMy5bQIZkvWi/44vyjXbw
RtV60WYjwno55glif6IpN4ZvH71w6BIFuU6iWv4th+4oi9Th0W3yVUGUB2L8gJY0l9BseQV3Sbb1
u1Thlnp1T6aujuM+vgYeR5ZtDv/suS5XvjYqZ8RKg1VYOvzZBgw+H2M85X8j5y0AD+WVBgmnOMXu
Eaa6/wRx+0f/vj2+u4BGMGi6IaBtY/ZgDrAUv01eIB+LzA1R6vyp5opum7ua9jLsLYwAEpP9bmwE
WMK0egxFI6yU1UVMAh5cocYF8vbWwvb8K8VGoDAYMEUeICtkNYu+KZPQNX81U/jI+v2ebExUjRO7
xkiyJ9403pzcqfTGjbBUo+LX4Qe5zDjcHyi+kk5k7Ef42jgc1cDYPpKWqwN8yuHq0F9eMyYFKru3
X11v1YoDMlpeLKobI0cmVVt0pcF+6BCXVcbMCkNQSSoptYrxLJt3Q2DEFFPvWvjF2mZAmzEfSSQZ
QyyhQRgWrk+YK4fEENCxRz2koyLv9KClRsd0vGPdMRobVf5MYNbasYYC67eOrCXZsElzX1gCqEpq
xXBPFgxAszbdBZwr2rfq9S29gELNU8sVH2SIzE/RTc+i4L/CLE0gI2l8L974753ELsswNoaZD94X
S8L6d9xYmalE3yq/2QXe5zjmizSQIHgtS9loeviTgPs32DM12Fhi7dL+i3rCnREVo1QgDIl1+3UI
y9jTr10K4TmeG072DcYMUcaBgZn/+X/5gKaRrzojOtisLTTJLHJJbf8DytYtSKQjZm+T+NFzM2dR
mW5A7mSxctbq00XhVuPq5euQj2wWijnad9X805MS+dTzyiR5OHp5jOnW3fPx/1wd0W9yEMY+lyVi
hciyrOFwB30Iq2H4yhyQyzvFzRIfSOCf5gExv7gJtIwte6CfJ+9f4Ooetd9zeutG/BLXcuefodcg
p3bFoDyriHwAkrzSDU3wIYz6kZwwzUG85kICBm5rPkX1X2mk4HhjKRjOvdtv5fDJsiDzbYSiTSoi
icfGS/qRfbG/8DsGbTlE8d9JeWDwDlnGRDWTAxbMP0Ya8w8891W4zn8bGS73XyyhWCFuQacivW6h
GQdvbBCKCTfq0frE1GAheo3xbhiWNdSM7icPbWyGvIALJwMgrsgNJP75MX/Q8HFahqCrJrqsQup+
iu64fTKy0xWAdFFP17bFMHDoZDTysrJ/XaoQ0DPt/6/co6DYAZ/5WLMFPpew7/SYxwSYmfnrOq5U
1/Lm8bAjB0SHrfpVpHsscUPXC4acvgxKeB9EUWwNs7iqNmSDu3wQfmajUllgGFtCy0+zfjkEF39D
Ypb2iBQ5G3M8Ky+DrpM/78eAPb84jtlZtEfJD92kUlIq9KFC19bmk9Kum7QXfSc9JmFoRC4lT8fh
Q5NhK7OgQAedJf/zFRNfAHg6bg2XocoUcA/X8ewGiDLPoAZ1FqocAteHyxJx/WEvV1AthrcdGVL1
eZmFSGsRcV5I9k1fwvPTgll0eaR3SY63B6+IuqUzkMUalg/llGSwBQ3JvugQUKUj5xiR47SYJtnI
SxWbd8dFxqnT34DJkS1VyDx6YMnCJYqJhGuMM39cNEOQ5XptN9pqIkQA31mKL7XNI/Hp9GqTkRVB
vwajCJjxt2XwV+THRBsXjiTFLcC1NOrmrcmSVZANzi9eDISmrPmP8EMZrnqnaMDahC4NdMsudeP0
DzSVv5e357zTRCOcEp+bVbKsZGn4HhD80cDof8N0i1qzjvNYl2f+vZYE0eEDCoHMLXaUto/bT4sX
LlIK1lHD4zqlBdCDOyjJeV1N/rJGHtmQ2plQvIra0lc92zxydnerTpauDqd07lIWpmhbFU/Eo7pK
d6YN8jjMmg5Hr/p0GDDOy8Dv+iuhzNlc/SvBdX0RS35k+j7ZIx5HyOext8SJDXLaMlJW+jOTHyo7
H9I2Pdv3uCbP5jnM6hShqcis+P2S8iNhJqIlOCwpq0xKIDcsaTJcznYhelK7LYcgVbdpNIB7j2bS
fRKIgtKbUJ7IS2oSytdUl/to7n9d65Hqm22lAa8gtAIBIss/klCVdmWwZ571kP5CKiH/ZGecZZ0B
XxRhonRhvxFuLZUFOA8DA8JDO45/kBUmpmrqONQeZFgbvQxMegKUqxCphJeHCwhtN6T4tPoC+/RI
4vUYi4CVOE/hleR8fJU1aOcQ/dRsxUvWjOVT7rW4ryYtSJvnPhzELOuJZ6ucWcMY4U5mnqIOQezr
sFl9cM7c5rs6FPKoH9/57Z2e18QXdVq5k4VF/05zdNivaVga9v1m+4XbazRVdFvWSG76cFZw4lBZ
cFPJoFrPpndReHKVKht1MEFYXd2vqZrC6zdI+HO5Rpk3jLGMBTFZtS9UvdXufgVR2F+Oo1MJbNTx
ywfbQHUrnyfenQSwaaQl1tftmqRLnFfx76/KJYXyjarcXhYK8KZTAvjrY5qGizRDlQx8FbGSqFA9
8GxaVCC7euldi7Ib1BC3PmAVd3U0r4jNMBCYAGsQ0ShuYY2f7NAgW9I6uTkG3dycQf84ARaW0/9/
j0RWZJgC9yEUVnizW6l94uPWBRPQJw375d4rD3XLVvTtay3aL6NQVmC2q/mMaShbyRA/EcStwGwL
wowxQMIY2TBmBA01wxeg+vNdLpPxb+V1M7nmWp+uUMG7Nbqi5dJOGVQQrlbr3iIseUJJ68ICt8b2
9eZ4z1iYQ8qrMmO5ClA1H8qjTatb38iJd4QC9BSWGQAriwRqwRfNXZHX8Rm0MWqgUIe/wHZIqPdi
xLvJG0z3bG7E0Dshm30+d1FwGhs/hNL2skIrXoxyZWrIXVkgw+aFA5nCNnNeXgfB3rYj+BtFAZlr
VmYFlicH2eDLoF0cWl84hnKPOwsREpINMVoK4Sgg5teTr4KB4dD9rlKSmVfgFNcuDbouq9MSYnqK
9m9yDNIAxqHh6De586GQv3qZ15h672QPtg4wZTRcG77q5PU1KXO1QwibFlDhQ7Yvhau0cTcVBn2p
fK8h8+0kyxWqR8f8T4isOENPMgAUCQU96PFVIVe0sX3xsMmIFmvJveQhj6gpobvqdJLvFGyXh6wg
8FZ6Y2tWyU2MtD0eQINJRjm9Y7++2pgRRoha62axoKpVreY7b2EsCu78r8xX+9LoPzA5iurlP6sI
13aplT1zOD50cm8M2fB8KrNUUzqcVKWcRhU5Dx2zzPc/PP6xj4xXbpHYDB3lJSDENCswlj4grSBP
PSZrKwfaA3FIg27AVkWMUr9LWwuB4lKlyTqKkS2KO8VpXis2LlVTK61H2jUEBxUDHU6RB7kRWrCR
vtk4iIoSXOO2zsJS9xHgYJaNkKBWWKh6WcU9ZcT8fxuuvmxlqyt6BtWau807g+FSSkEzNllXGzMO
6pei/V0qm3BxH3SQypHLH0Q0pHqmLoHZRtxjeF27I3ESdvT2Azu85tI/jhnTFAgTK4yXP7grntcG
2tVYKpGxRHgincAdBQ7eAUP9LuQSWrAVAntS4waA5bQ1YAkkdh5e8/DEAW2m+/TwBU6Rn5kfn7w3
4SXhNCs5FYKB5R2wUC3zS6dn8+qqxfUfRcG+2cha82VkJV71kL1QZrCUBDdiueAAQAbQGPtA9Lf6
0LO/zbVXfeQTJXOQxh29C54gM3F7yycNBhAHHL9Os4QZzreKtwOLi5HQdyqb+XChszviUYSawwbe
UJiljo2Nz6wc8ppiZjF40McUo2cYdBXEJobuB6pJA0L24qI+ZGpwdRbtg/7iKNy1qrwpXEs9Cv9W
Iw90M6EBy8JZ3jpjgwn+FB2bgVQ98rAFheI9mNdTppcvv0tkXgfNDyvpJTF6F5gYLJJZZBykqme9
oteWDBiZx42BLqVH+G1/ZSfYDklha/IIbqnQJTpPPhYB/Lve9bQuXJgtkqO3w26WCkpUfcX2vy8n
ggvE71IgJZ9jNxGqX00jNYtU9+JHBp4FKIxHZohVYgkUXuzBy//adjPweUaKjwARIJgHkd0qnOqi
5P6Xh8hRtylWwBxE+zk/AFSIE6QxI/GqM7FFtuJiGP4OuLJqgfjutwTTAL1rwx/mPw5bVWXwlhsl
H9WgkPff0VwStQh77fWZTVeTMoGfI9GtSqNl29h35q69vNuQ1UBUackEtl3VNYP+Xcimnpu2GF5/
RYl4UxSaYhrRjOYT07MWjLxYN08oVEu8XFzitQ8sRW4CEnnP7v6mmb8JskRZE2xxXQk1WHEqRST9
y19LFmjvUXRWWTU6FCK2gqJ+CMWaBHhDiSJIWZF9yOU1e+3wXv1UTmhabHElFfrYo/tkucXUHHzK
GRnaP4+tT1hcHpR469ohShvCRXsjIhNVFEhrobok+Sonmh/QFbMnb2F75ZTb+fYM1T2rUKpwvdsa
TeGhPlXnByP7IrnEolu7EbsVsEbSt6SjmKFxl+i+K8rQfdgCe5sDRGQ6uVrETkUQubNjuHkkXQfa
k6EWprwHe6nESumLvi7auXMw2NXbKoIM0YpUdmOly2k/e4EVv/htB2iOcm/RyuyRZpIxbpC4ZK6f
T+09SFpErbxaGoI1cFi+v20L5m6xZEZ6i5hYwlQTaaFd7p0F16wIvTbRQ40LYbmDLXfpxfD6S9MO
6xAPq5Vy+zndqWjErrNkhk0+4DrQI4whm91EYACV6QdYBapUtj2/RZTmkz1n+nhOA/IJLzf6Dfvp
A1nLWVZ1dnNoPKnGaoEhtnd+peepnJzLfOymntFIScNREucv/Qba8ulpclZSERuW8NrWU8q7zXND
MurtQZLgso4G3i65jpFG3eQ7TngPZKNhOrAnhTic75ICV/qD7gVSOsHxYk1ZyxatWuBpBUIUgFOR
aE9d+JaqNXvTU8Yr+wQ7G9Vzhdc01j6UgJI/n1Vq7WPNyKwPoneQGDGS96t0Ak7/vyWCuDLXJxD+
UD1nYglXuzElr5CcCHxEPnKI5yrimsFlybfAd68m3VqH1ZB/SsCZCRNqB3iavRtwzzk1RB31gjIJ
JO/y02OPPAzrgppF8kucAGhmBLz4R8cxZKf7b+Hj7ToWN9tpmWxUjpvcHfwOJqph4tvKQwpIHvT7
Dov2ssUYus9+iRrrKHRIddpdiFc6vjIax7OoY+9rxW8HdBVrgyc05RMeH44V5cWp1YzR6jtETG1S
vfnYEaa0q2oJN2YuFg4/UX5OTasJPZB6j7rIQKe+qC9kyYo8thsnXD3J51P1bMeV17I07tbQ4/Xx
6/umbxBMhT3HYqxMXEXEQx9lNQSLhJCmbE/PkOEak5LQN3tEkWtns1i3cCn/EjOBtaoRDuwDngbC
R6zm33lNdEmI5BuEsJagupVbQkurVgSZwNHsEXY67yWqtyEGwzld1vkN5rPm+Ndl3GbOViQuXvFP
c/+9HSa/sgBDHK7LxC0F3wTQDetlE0thjCF4kcXt3WgmpIRXEiT7SX1N4qiooKCqCjsPLNwlaut7
vU/0e+3kjEiNAdNPGcxjy2UIBTv/94h8lmFSvzeQbXf+GVcE7SQcM9nyF/BMV0TFo2NBYGIIuGqW
+Jg+3VtkXMrwej2obIpjliCykZLnCIopNXk9KY4Endn3FZOUt2SMmdL0nMZtqeqUOYQb9HaKcXxK
wG1J+x7hs36O9xbHM3WpUj+yNdprKldwtPeBuRN9meraTMV/1gwXqVH3/ul1RCDt6fNfUqM4Coy7
ThuZ0ZkckL18Ogpm+EXhfIw2JPkq5YSze8I19DRbgo1N94VDyxfB2evyDNdaYE0bHnT+GuxGxd/M
JBv/bA806Dh1ol6R2yWxboxFi7b2gHh9mR1K9zHQyf2NaG/PkPYlj7UNp5a01T3qMAJFfLbBu6hB
tLZ9w+QIetRJreBV0Td29ch8I1K1RT/GYyFGJYw+gYTiTnUAbGtrgPuPWrM6tCUFC6T2uqj8ev0R
bq45MSdkP7QV2zUYJGr/pp06pv9/TVVICap5M8QWxD0xSHP83LSdrzP9f8sFc6sTSZX7Umu505Po
9Ov4H+3mO+Elv6oHKB6saiSNE2O7yvv6MWxd6TZ7tKKNfKx+xzDSOGeyZjhmXjZB5dqsWe7/koQs
/EZls1gJynAChHtI8ENRzmgVHG/32luJK+SFxRyJNSJ7N43x0L8ATqAIURLpOyjyJ3VcBBEKrlte
FqO6/VeVUGnH59WRydre/tRs85hfSqR299xcTj4DW+qd/MfnvbDekAZjXrVL7WvN21z+Ew6VTriw
QlBaJnkHX6kuzH9MpB4le6pm2HZ9dxdCS5QRhPlxglzWknyrxsIa4SgUtx9m9/jqBYU6HkK2O5ty
XbS9WtGPoiuE0RDunTDJ0U8Zv09gk0e+CU1YSVZQdiWqZ7G0OkKiA0UaiWxcMR8+0WWTiV9JW098
sdB+T1UYQJYfKRn3HYg/BIOn/s928LodbZdSKoLR4Q6ybCUSp7IGjc6MZGgT9TH9C6nU7e0lqZd7
MscCWeLFFT5s8ZEltvvO0kzvbuKB5vKdQdXFcOIpxEQFeniJbtj8I0Z6HMqgrCHbINxvMuLcaDX4
gS6t8OxPaYW+Ot8eGI4+k56bpEEr4gERndX38GQCpXAwoHp0wHcU4QjyW7u0fZgtYPBqJgXUUiEV
h8xycJ0IdP8SsxzEad/Wocuv3l5p399rUuwWjeQ++6zjLgKBHs+qVBBLI1dISsyHmSrjekCuRGUo
oGAPMMXhKo+ERRNfPlXIjHKAJXAJTlTX3i23c+beyh+M5oUKSI0ScRkZ5cGLWPmn6Il1C91GKVeR
auYD09bJu529ahHvBO3QN96r0fjGq5rmxhiUe6grahIzN4c5ny9mCjD6HUcWpoHBtbKAao7o3JzS
OmHzQga9w9ikWAxV/akeFtt3X6s4Prxy4IHuX80bvR2+tsEsfxWhEW2qUkmwR1t3kmhZshBMwKBV
mMuYZseN6AyRJOLqe3XUMfNito1xQkpvGJOIWPoOXrBwev+1ARHFRnuwkrcYOj7RN96PCtpQ1xpN
IU96GGN7clhXV183Uom+2HPk6V5g9LdSXq39aWcajZdst/6Tu1BH6xon+wqPE9VE2bZO3Xo0dGa7
C2UlxOOsz5t1wAKJDzI6TEnZfJU5Xz9d9HEN7EyZGba3sUnIyRNjgC5uubkyyUeyvFAWmBB+Xxuw
uh2/iy0FaBcfLu4gAS0b9u4UqMf5drviwQsQDJQ6Unx+oUUaV+MRhbllZIAdOby+/oYM1lkhGFXl
R+j3MAaapohbqMkejtKrLWYMbZF0GGAqiKDROmfO7MCp9/KIzhjnoXVpntXU9SRglaJ989OiO6vn
lmEapTs085Fx5ROhj1EzusLEkEN/v0rEruM2fGeOL/khtCEG3sukC5orvBpqb85KXyDQsGxY0Mcr
yGh9F+oevGhmbtG+oIe9OS7gZ/stICiuEcgEUdNCfewsYO2RIhvhHQBtSGRG2vSHS3nxti4o7Vzm
zCCAtOwAf/txrooTBwRgUqZ/rAsnOHdk912brVPRR2LK8FwC+9cXmTpD6EEB4s0mkl0spDtSwnlL
BBOdyMEV4wZU8wOSGq4n1xwEtpRLzD4RnFSizzQNVeo84dlMI+lpDS0drWJ9VaAPcH9/vEpXeGr2
SxSQ9WZ3FFUjN3t5kM0CjSx1o0JBiay/6vCVE9jHjopwAO7A+YMX5Tk3bl1dzqg4jVtBVFKyZbJr
qUXd89U7DOmnTxIlz33zrcJFIWewLImCeumZGgdhfKKu6j8bVa/vAdvXATs2o2W0zTvcMe2BSu+F
32xOe38ARvqOyHBHtFMV1NrGCW1O2iLD+bmnIgmRhrfDDdimSiA0/prI9WDpwWmb61L/bc/EWdqa
mpasO1XQof8RgevmKqqDhc5IdSPdtKSPd+HjdDzXSdjIq12Oux6GLF9qZUMGkYczK1c1xo1v0yQk
80yC1bK4dctbvMluvgIzjf4Aj8z9zDDwWIFPiknGIBuVJWpTi5YlM1XPmXhQnrK9HBv1wfYR1TTU
mrftU/crPwHdY+jHJYDpkSHDoXMJB9GN0PN7IuhVVFvBbpr0KElPq74yguO5IR8xv8vitWsay3fB
Png5o5Zzll4UEZGAyN1k1f+Urhfy/zztQ4O58AyU5jecaEs/lJVUBwCigkSV045t8q7jzMpMP/So
2ACQ3nj+8XH3K/O9eF5Bw1YEsmJM1zDKlbJvQk8XilZ7uninv60DNoIhCI8hWBNB1pm5Tzf9rA82
I7bYzGIvK7ez0TapX/z2pwDX6Csh1YHngk1ftqdw9eEDp7kFoaIQ10CEEgYnPwMj2lWVdITEyAjV
gOebvP6iqMrcymq7l1V2o4w6ort3jHtFH5vfQQTK/TUEIDuXUWKgqJ7lBJe2R1RM47OkXqglOksl
E8gjz1TuRAZmId4LKIL6UkIKfBBqx+zZsj7QEdCvTlVkP7CKnNZd+Dkxkaz8doWvzeEykRdEsF9z
BCd2cvRKBxgaWfRUKkrAIq0PDUjfGHj/8JawlDORTE8OmkuttqYRPuKmTFoboVIxBZVtTuQWu4cz
JUfo91U33O2O78sErfUPMmIKM9dXUTSaextelDSem24o3JK/weQ5sOh2j26UbgmSV4K/pTeDe6R0
c01Ez3zN8g32P7uMcpGVDKS0gnJOFtI0yAxCA7IBIFsiv3meXk2VMCj3UabSmgQ6mDZrXwVY62yL
BatFeR5TruqeyioN0/YXOuIDh5pZDDHpNeqXu35hRo5AdP5F6D7CA5B6oMDh53lecapuBvUMcdl2
jOa2oVClR4koOh5LY1JFm6YPQeTLyi8rhsty1AmOuFL4amqg8g96YTeESnBHW9uASHawM9WiJbta
j2CmIx+WHoW2KRlgxJkGfp/xIdKKWu6fsBKjYRVbxtjPCh4SM/XqJqgU4GE+9AQ7gMjhVlMVbqKc
/zUBEY1XziuTtPIHsv8L7GWNkVDcUonm9I6IKln9tcxD/rPyv9hZ5FrCidP1Z8DcoenVcas0G5Uq
frucA9fXnqbgZ86JFNl3Fez3963yPuBFctxJCZ8WpYR1Wp9alEAckFJe6bIib7KjInuq/bDeLrE+
/vMJauXsx/DP+tiYo6YWCQgzJArU9ekF49uor5UD+Sz5wWrG6cHI67GKdNBtNgyhlZl0E3er0C6f
meD12O4Hyb/TZzEatVnyKWtLa28PGlFF2d+0MLz/FlxIpY6SBQnFx6dY0nPMUw02jrS6jVouwQge
oNRWFydiABz8YAu6peg+dEg06+/iKw+ok7y5QMqqaAfrmRuAKDdIOsN52I55L99m4SJCq2Opk1iE
WisdZxSLTz71TZdALnpU6W97F88bENuiBrY8fvgnEQrVsVzLBhMhFlCUDH6JzHGtgZZLfHAui+bq
Wyigz9YYaeSPcDqkPDdnnAZ4xvJQj4rU6AeQrC9FX2esQVUeSWtxGKDGRNsVP8gglZeQFxDp9t0V
3fzwqSMbAjJ0Z3QL7JA7mU1CDgRhLkl4kdCxwFiMgEImGTDKFh78smwCUvZhvT6NLzc4kq+IyRLO
oTamou9vw3HbvRGuGB11MJ5BuLV2vU/ZHUbFLL8z/k/g9z3UscDCMZz6lp10y1EjvQwSfSgf1rQ7
yQm/ZeORC8EFm8sri6PMZ1pAjWax1/NUrwY95HBLBvr9bRh7w1WNwnVa0KRFxorHI4A9ni10yRxZ
fky48uPMVrRyIoeZJbvtCz+fucc5dxiQvJNAp+TE2dx/24BQBbAaZACgWgmp49wCXYfx3oMA6WnX
sGUVE+1gC8Zf/fS00jSZ6+rccpkDMuZkhpSMoelj0PD41lS/y2aXAajD44//M1JI4PSNDBurQE9E
54AOCAKSZofrI6/T+qvFVqtA9YEjJFUYtUnHHAQtR27KJdBVVUVD5v078tAkZT3UO5lEQ94I6tbr
ZEIFHLNCSgaticWELTye3gfGjDQUR1EirZYEGh1Pk0CXyXGErpQZ2CWsZvxFb8QmWycfyS7CGWcL
/K67AvzMqCTng8iAoc4VzaFbdCXpJEYmSl7J5PxBpmqgUopdsI7RCAaPOz8dCZiLFIG0LSpmJlUY
OdUNCMkMC2dX67y/8uXevcHaYMZ7TqoLR+GkbyASsTM5zJRrShI6lJFdWHKMDCc7VBbmjTHDe7h1
2sgJPOh1WrZxCA6IWXw5hrBi+oL7+KCe/CYTimKr/5hAl612o2M7ctev4UVCXbMBB8F0v5BK/H+l
7MVnXe/g3Br5Sa2usNwQqjkK54dRwbqi5XtaxgtbFOgka/efLWakNeU1/bEVWS0YCn+a9ZjG/1mD
Ptxxq4ZZn1W7z6w4nLukV4hj09Nk3SjIQd20GBigWg5C7lSthe3QRmVsR2TxKhtFdCBYgTGpggju
4onEp6mgCyb0VVVy694ALwmPI7HlsIkZ0baAKrGRXYZ7HbtzojuLzbzB29Mrkpi5n8AFTKN+1sQA
w4HQyz7iC6jeUFP05AWOgophcpLlylfmvd5rT45yCIxNBoj/rhMNOhzbC035MUZXe8/NZliFNUSu
MQXaMyT6XyuroZu9BpqhSxJapzFFueTh91VSe94fNqGwq87y6nWv2uJfBBnjjSZr3Ob4JuKSWAvO
td5+27NBTX9lGa2ESr2s6ZGVgjMaqTg0EXhi33KSS/X9BXU8DUv6ICOTi3nv4MEGXwUyAkdeE/vn
lM0datEo7zoI3fl6xkKn2D/kruN+Gz9Q+AxYRnHzY4AfUEny0dlCJC/rIShWz+UYa4GweIYauB31
sGyvw1HeaWMxNogvPdM/hyFm/MH1Nb6YQp06CGW145C4jM1cF4mZ/IBb1PuV+xJtmmqNAgIyhaM6
Gr3kHmyF5AYm14duME3LZeafeKeCOEj6RMJAAu/GNoggshWZi5Ocoz//fCdMbP4Sbwh1RADh8ia4
ODwsRGXkQACrNDuq3yMYy4KT9P7AutWMkXUrxa9CxiPasvGZbWAz7pAkbwMdvi/7brgfC3Kz+LJO
Sc1E52Pz+XopZZ5wBygBNiOb5kk2Z2srDFCZ+l418uQdmc7e4YPo6FcbK7PEp8bhoUjVvUQ/mZFC
m/SRQQLpAe5fELeeDJaBCqBGgdFa+giC225U1RDfA7HPdS+NZBqbHXK7fQT2NVCVArLfGYdfA3MT
0HrPzWr3wEupbzW8Ykw2uxXSohxv+B4q8R5Z0CMYB5HU1DNEPf/iSKKGslm2vmML4ZR1GBncNr/F
slm0pNGVdaYYHvCR0EXFc2T51G6DJsHzNuZtgrMY0C1vNvHaviwKr6kZJQrKMcVvn82SD7rmhPlF
hJsGKHbnj+a8Zvky42+FoLkFTSuswAm+/QNR0nL+HZ19yIW05UCcMhrsTjtyFqbfTQkYAu6IbnEy
v6OiUuxWXlfuYf2W8MHa5vcpQ8tnd4SNvCY1Pe5Tzu8Nrj7d4UU1ELP4E9TrHbKOWHNeC22s796u
Ce7lu4K6rzp0mTzhfjGexqERUMho47iyGzp9JNyA5oEi/MS/bkCr7q6dnMsgh74EfDJDVls5XdOg
lF6mRW6da0zFaoqS25J0Kj6x3Gop/LE8ZFFMFJxNEWhAGHUTH1fFcrteUoEvi2nrxc2f9qPd34ur
tD9G7elLj0Y4z2BJjqd7UiCc6q0VCrrJo3qCpwxgRPf2sA3JbwWrP+Nhtru59ZxDoGKm8sxyhTeN
RDl7htXdQM5qMMORNcEcGfYxhYsM9MbKAeOCc+rX+KETAnJlngQwUWq1EQ24ZXQ3kNTq1iuvdDP1
han+YGLl+vpWxabU+BxLUwzHvAGuzTSTL2SKaJQ7HAcqh1xoO/i7r2UXRhpGiH20fg8a8lIXcB+M
oP3EIiBchlVj/9iv8ORWiimUZ/g3VAYbp7AcabkY4/NzpCAcIF2gHthEQJJNHT6TPM2NGUzye/2r
U1Rw512ZAjn5HsvUEb2LNFhqZ6LtxIzhvE9sUYa+ihB63TzBxtcxWAEh2rLojfXYvq67KwQO+1Ui
dYQbYXG59hlNcJWkAgQp0SYklBRUBndzr3sSklOXWO4SZircqU2OA/8N+tGOcRa6Zh7NzQZG02sS
ihcQmOPHvG5f2ZKUnYmlMtO5CAMWucRuee1aNdkwDZsckfJdMRyUZdfxTOfS6ZFTzuVcvsQuXYcy
Vn4Pd2MHq+jzOmM4ZsGicvmhIQUkNxWmcFaa7FrIdHgrvi7z+7Z7de9/Gp/dQL6TuBBC838w01MU
4Isi7X7ZMgnqG1CwydG1VoicYNVtrCxNrAa8zi9jn3Ut/aBAuy7+tx0RC9kkZz6oPj4Sur0dkdMs
Bmq2/XKQOW2NMEwBKkcTHvQvKX+Y/C+wdy5Xy2zn6ZJPyu6HPHpA5Iyp2+x2IHMWRWAdBXnuYZ0g
ieFYLJ1yZqYYFVnxq1twFsKUo+kvvWzq7xHex7DrJZkLmZ0byvDE8i3FuDDsQ57Ge7T8nUxFBx73
H3ZpiK/u+xLkDaWRL1yoJnGXi6TINU4dFY64BsPmCgx1sioSWa/Zt1mNew0kRNuH+ZjJisEp4DQM
MoPTgM5Jjz/VBKjyOwN4ZFD+pMXl9CBBnqLSjReBlJXBlEUX9Dto8Z3+QFfgqrsDPB7RT+/3Dqap
4dzpFjCg3MpLDdcgdVwyFCWHW6hXHUbygHZ+lpJnnBOGPIYzWTQu8NLuZUfhBE3xooB/aQceNRKC
9ZQV4y7HUcLACOxIzF/lmMtQezfdl/1XAsKhuaUthCWaqnfT7eU2066zDz0cvAo1krWTihyQb33h
Z8ceBZcDeehujKMUbAZl4e/6O8/QjP4JVenxx8CKyFfQI58JqryA5MxrCng+ssZ9blZwK4CIHsZA
X1jyIaR+sI4Gp1cfGDrtfQ+sRbsNa9H7JAOuNLUsCDnf/izJKJ8H49OHwknYlDUE7ZVjaXbD0wLj
f6CFxS/n/7cqX5+KtH8y/y4/S+WX+xWEk1MlHa6FB4Uar6SB5TDagi+ot+dMat7fvCWhChO3wrLu
qJjRUxG1F1by8hfqtBXR9nbuDGM5M8dxrNTpMWMYkBKY4wuJ1Cn5nKJ3WLRxQsDnB4gLAnLTAcsO
JWioQtO4YwnlfIjXblpidWRNZVWu5DljKbzSmKY/yRCyqfY+h7GL66sfGt8MSYK+KQCk55H8ypqy
D/Ak43LCtJz3WtUvqL7r9NKUJbqhxOJjymnfgCQulQXHqEP6/LV0UmwQxPdTvtFAmvVXFoLqKPbL
nJB3bOw+3bSKppebjD2t7+g3qUARQA48oiQ1HCTg68ssX47MwzrKdyrDkbEcSJfJdZrzgYhA7gA/
l9ou0TDnK9FV0NSaPnsqFyO0FwDSVSI8oFIYSKDcOF5/UDQrunj51dfB1iRY8RHZJb21vTqNvIsB
vRwxUh9gbmqRYCPrleg4d9Wty9xZHSy6PJgVgWu2HVyGjs0NeRIls4hsDLfthqn99+YQPv2FtJdS
xGdD58+gsFcbwP/ViD93u+Zr2WXxjQvUMkHqHiTIXXWMFh5LmLKGWsqgavhvUrs46Gui3/YlQGmr
KlK2+zkCIMFJ3r9gnKB/3sIWaJSgztfhq77p2z49vyNeDe7m7N0Fwdcs/RwoD+eE1Ck6rTRqf9LU
yzoq0oTIrlFyfwW4xUn08laugBOQg6Cd2VHLeGfkx1Sgj1rIUr19sFmdj7A+m5fr3xabCLWYxo2V
tAnJXN+c97KvRRai/bW+h06mPUZBowPO0VZFcXp+oK3jDQVK8xMw0smgwmGNX5pvy1KdxrcCe1eJ
ptaBy/AlgCaO+WoxRhUbwobv01IqJbltuKHeYrFtCNS45SLmv5i9hn4oBtXC8LtXTI+s5dv9Z4TF
EY+AZvnv1QbH5lMHaR5AoGR/4osDb68hLZcdl8qUQ+4EEJ/6E21/m8dVktlxD6c7v/UI+2IftNpA
7Q8YHp6gljDoRw0/FrHHywE1fWerKQjRKvIStbzOPz70Tt0KgCUmlap4FZYBAoFunP5hTyo4WMMP
csqtP6ZatRk1JOHK0pzp/zwJLdnXot8gBVoi6bKnUvTXPE8TVbexrnUXHrzi+s1Q9WZmGOgFyeBV
EImbYs6tMWyhIHOAtPRNI5RA8vhvtHQYo7RfD6XEESEdzN4ELfFfIubmBQFZZEwjV1JZSSN9+ReU
TXkxzBgOsn31lDF2ujmzaRQKudxsbEHCib2qcx1NjFPZCGyt9unLwyI/Fqc5li5M/5gPiwTymFuX
C+KgK2eBxIrnbMm9gHxUxdEmS/PSjm9Iw24pPEmp/BSw2mvNYTy7ocnN5QTswmpQ3qmdpGcRtttd
zho6jSYN8sNWf+t+CPCMJpJbFbJGjLeyHZPXQDdLLVotqsSzAQEEDCf7/YCZ9WEslrk2b5HDHM3X
BZgAd1eoDm9jbnbM9YRC8csYQJh6XVq0pKHx1aGntTUHDA2dOU4DQ0nr0k2yGUUT0XD2UrgIYum7
M4XSeeIizH/j56dxkoTr40YvSEQsqBLDc0wg5HlTOd/qSRxWxxrlVbVR52V7wZ7HZ7t5qG+ND9CP
f8Zw6ggEoBDp0W0SMB9xKWuipEjqUO/oujfm4GtGq1fx6/Z8zBzpQk2iKBXNbJNN6UTwYJ7hDrTr
R8ZCELPA1FHX9xRMxWkhhHZrAJkgF0h2RK2Frc7aATuZmgQmRQsA87XsxgRhPUTkDDH39mCHzC1r
NIhGedVQq//fd6Mxtx1lNcLA5bgIzeEigMKpcRbhLSGkZuL/Lwj/3UpZVZoMhWTWw/ZZ469RZ6wO
WtYEuF2oMU8/luLIEbIZrkeRIceNSuDqA8OPWUE+eBJZc4RtdHACEcQePgZQNUcTzlDn90VgtDvo
X9AYv5eAkGFA0L/s1gYCKqRlyhXq51c7Y+DlDZZAxiRoi4d1fcFh1XmkcCJgQkp+uvVluKsUNwlN
kH7AYZ8hNbzvzpxLHDnV0qeTcOzsHWW5YDyNucuotnS3uD29SmvyARLOzwR8JODzGAjgHaLQE+Z5
gVRKnBgFkjA83sC03SnBYbYeK1jzijpX3N+81+sTh18NtayVTY6ej1j7EeiJdGfJSCE5P22/ZE0m
I9it5Wtxli6F7P+vRkFm//8FEnt2Lu286qj9iQZf83C2ttWdT3hvgLC9ivARuUdQOPf0td4muNVW
loORNuVygp0YQvLMHAfXhwopSaWfozJ9eAFS+Z/J8xVIBOIRWJAaxGojuK9gz9NA9c+DF5UG6fyt
oP1MIAjB9eUM3upOuTqyjkUNWEEp7EL9JusvgmfcYlHvt0h9jRsvbSdTrSR7eL8d/bNgVXQjx9lc
7a9I3iWa+v4AmB2VTSDW355SDOUqwyzKYCZxU+CjcecKDG+en77EBqoeCI+XOU6U4sDyby/tZBA+
4TJ1t/ewgZHE2yawpAqvCsDFMQvybY9KQOXPJYTkAMVsPxCu/eR38NZyfgAjrk7gxC5dFOqwdooQ
2XVop2XTj7qqbHbd1KI5yV4Ah4cV96jenMxW5QS4rc4P9CceR3YjJoN8WaHU7S+1mkDPtXdnpn3J
WAzP67BgBMKqBGHsQDMotI+ikvYIKV0DZX9mQGN0rXoeLEfjcophYllmKD9uaFcLpCjiNL55TxU3
ThqjzXChocgxOc0XxUgrddgo1MypR5CllLnKYmwbAXrakTMghDphbA0XjrlZELnX4nTWv8xf1rfm
2k0rF61FuYEJWkEfZOkkuRVjjjRbuUDsNsgLJRlddLQRIhGpPdFuGrdnsccH9mYd6gzJcMPYZ7Hz
7U9YAtNBZgcJshcvR8PQL/9N23q2NRvLmdyeyXa7aAm+QJwKNzsbyUrV2cjw9UshzSOpjhsIxAco
vsXcfdjuGRJ9KeFqPO8GtYLIFkkCtXn4Td0dmcWdbZcYozVDz+Lr+CVVoQZ5QalVOmMqUCEAHzFg
exbQ6oDZv0hceJaIVK8Vpnhh1BNiPqMy46ME8iez/V1Z7ZBCwbIaAxmgLs5K6z72m1/c1vzkzRSt
rqv5m0wekQ61PrFgQ14F5mgYAKbWMbCcuviR4X4qeD4L0H1D+jJqMILC22IMK/Q2AQQPKGFyC1wZ
O5nMr0SYIEdPAJYc0ze4o8k9J6pEzMd5Wutdyo9aRzKx2cOI4Y6d93jjdocLe5Fs6rF+Au2pYwB1
5qaPB1lsUVI3inOqS8YwuOaLMrMFi4RN/J++oPTuknPvZKD19pFFRnRbTdBnkCx+1K3YHPtPEWkq
ISA9FvKkWzMZo6gbMp1ZTXlHURugbMeyDNVYepmGdmClgBv4rPyspSnRr606nbrOoBn/ZmVgJQI0
Uo/0/c7RgSeySvi/pY7NfeL0N3vFrXBqqklHTuWQvhp9fW2zb+Ox43R4wmTR88jlzkWZmtzNeGci
6qT7+yAnKaOZMGyQdqHcq3Zuekl4XKId1pl47yMxPiK8RNwMJjY/DfHKKLt3y5QZ85gcHBsilqJx
872tgQb+hDQu1LmYNOrUndPnkFXzTGyg+UKpHw15ZzGyGSSeXEUqpRvbfRHGV/0nBZFB0jWauvFI
wKaLLMF1jiAmuiulCzi1ssAVWtn8CAhLVYRDJ99x+sRUId6azIlsLG6uVGKSZZJZZ3S95ew0uliw
FJAbIQNEFsMSTEC3/7sa0p/X4Amcp16EWeElT98mo8Eb/dN2iRpAfpGH8yQUw4LEtqgKX8aPXgkG
gRkRTqSpymSG33HlY6iv7oZAe2iI3Y49Sg2vmeStVeGYujNpaDgkdw9Mqq29dANley65jzzDLlwS
KOrD/TV784DrOGNBSUd6yA7iQUMstgGZoLQC2z7I1T4asvjYO9wFNeeVxy0u+/OZMnQgyhO36gT5
DTfwxQiKc6TZu2wpv2T5gfHYBlWkB9BA7wt7GnHqsOZfWyxA7+gyRFQ6axk2UuxQrJnBEnJL/ovE
/QPTdBZf82h78VR5jXwPCzp/9l0SJesYUluZ//6ExwymPtu4vil1CMhmix0AGwsyXuFwmg/lDzFO
sN0yZrcjoQN2zY+hgQM9wZHQpYlW42YaU8H21tJYRsGsh2jjMFhnYZV8HZEPq4xxTG+YuLRaE8NN
xmyBiu2lFJ3xkOYVnf/OysVtrAkdoQPKyEaW2szlVr3755ovCAZPX7fHw/smg9gla17GDovSh1xj
5fqxZ02JO816+VfWUTMPvPF3xen0wWOp7cG9kmdJr9pwtHpJm+7SLgB/92rsUWyqYjUQQEbsFF34
N4H2Vqr1S/UYNHOKEoeDOVDNlPpktLRm+EfTDgB0pFGYHQ2GV5xiRZucQnOCFhEgfnWCJJvnus66
MTaCFSSO3+rgytxp9X0LCOg8MDDgklqPouk/+rSRWoESL4fcXrxOJDTAioYiKKLGy17PkXt2vBCj
4PRVxBqZNb+JDeseKr3BwCGzYImQ1TBfe8V3gkuru5J149y/suY406veTXc34jDPCsVOwYMXO7XL
ytjobqVo/yETvP6Luqv/nRgzb3EAbLTVhK8939hHRbWtR3SeAcFpA35YZrtF4wbtKq5N92qe0kCE
3kOlhBgCAwLAcfLc26v2fB+N75UCxXmcUP7P/FQ3XR8xMx/JDviTzhrxKkPFn3eiQvZDfqxqGqPh
hS3kXuL1NO5StnJbAEYdWCIYGrxl4Ao2XrQVc+XDnk3DcgFRCacyQpWhW077xzk+tCCBsqEYUdSL
foVGQLUkY0xFQ0AZcPdy/kejUFXJ4/+WTim9q0I1NrFu9XV8OY7IamoNT6ExYtXJHojSOsGhgBVS
hxxivYHvLIQoj/dvbTTJaFH/jNhB2p5SwC8sPg5vddxmiJ622eIU5EWDK66p5kfsYuw+edOML1KI
Bb90O4STpSaew47ub1G8FYMOryvkbIKLjhACsuecbGzGbhSt1MEQvAImtm/vj/OXQ9N28JMu2168
kkRKnIO5ewHtNrlcXJhZEKfNnztF3n5drEb/4lTACyBzgEyYejYwy2bkk1GXY2rOuPmTJA2doF/O
nMkLm3puaDcvbPt+osYkRdiqqy1TfATAAJMjPIalODBXXt2QErMZlNJwSgR0lrYThuKiun4jjzLu
vVUtyyF0sAyyEo0JnijKygLJnmaFYsSigYTAxmyLlEWxPsXPQwGIvJfZgSvSA+DQYvslNSUdXu+v
vmZxCoTkeQoC+5cWnvTasIG0WDH0maDXeAXRVH/pfPL8D4YPmlfSeehheRapNh83OqwwyLUfG+1l
ykJrozanzR9q8d4ZqqUI03kSfgYILgohrAOeDW1aNAkJDIHl77siz2BQwnpj/LlmbAKdx+feEoBj
NqGXn04wWQs39hW1XgCjrdjuYGZjXXmeqZhNHcucW8+n9Ih0afotciTvUrx1IFjwHtF3RxRCuEyR
HGOtx9Fg4q3uoCqt3IFLp9NgIEbNvudHGsKIwM2Uuqjv638iy+Gl6gMUeAERt0QGqQqT0RUpoEc9
Pipj5XHEbOVmPlY8fAeuyUuJaxAHwXnpxrpdLdm1jDEuHU6x99u1T4TdkBuJ42t9sC5RKMablNiD
PSa6s+jqDTn4gvoyFeHmYLqTNdEXpAuWO4y7afrg1mCJGjA0WQxfTdVUo21R35agSbwIqWmdKX9e
MKHlXdjIvPj+ZjpwFb7tPky6gRkikpkTSG7nrJaW99w/NW7x/uB+3GJeSJdC9mPL4SeAmg3De4vg
icxytgnGaje5YyojPG7FdJHAYSpUqihIDF70YxKSID2WW/LVsCuY1RS5T3SmncpDJO93zMQoXtNY
q1Ihle2qous90Y1nQYnUuGMLeXXPRnb0KIPa5Rk8bm926cywyUyDc9Vi+F5AHHbAXT6VbERAAQme
FDSM42SXktiOGyFr954IfTvPOcFQlTV3f1ktizOew5L3mrIH0kl+ApVQ5bPCA5FFsQqDLc+gHLwA
jojo9/UifE1HrvhPn33To0u7MqhyxZwFTt9w8c0YQH1CBjvfRfRQQWAVS7LjOcTmhELFCINQ5cbB
K+xHB7y8Oqred6r0cmzF4zp3YuZ/EdTbrOSqygCSCaFauC3UEqovZhL6gGM8wT5K58R/Z/uClqvl
M0rdf2om7OVk/70KieQky/cJktcASkvpGH7onjqIfd6T3pJ+XOKUv7dlLpbiaScHtaa1ZmlX2OhL
g3t17iPy3eiteKRacS3l1rAVNuD8k/u5cQImPZ05009NzI4IgDqm7IJAFlHbeZNNwJI3ZmP6FSTY
faDnri/cAi/ZKctib0pQZT4CrZg3xKzZmmjLJRJo9OR+S7JSipa98OCwu7A16+lHOGW1uNKZsdv3
nUqQpDQldIB8ibk7dm8lYc8heK4Sww6lZ6M2LgU5LO1gx4H9kiqJEFoHP76mDjK+nMrm79KJyGTh
izHT8EAAn36aGWOQnvzqq+gwDpo4iQDd1nTD5DWUDrvSjplguQexZEBVNZJLFCkOpr7rD7hc8Ugv
14lLm/PWeorYq8srV/dEt4ZRxUH/8L9qw8CctBIxkK8jKluo6AaIz56GBFt9n0FJF62+ykMtwOY5
dTNypBN05qKQEtYYtEwp/apGzf5Is9hUX/97EXExuGDK/mDFYOlhIytTvvuR1CRWP/XiadBQNdIV
wQMzlFKglsFexJ3gHgpaRxmClGz3+gOlnJQbl1C9/uzxss2rPQGRVuAhds2cbgrTInvC/jwb+qOF
RYujb0pyoGamW5rTopafFTtge3bu4FcGfWorT7iQiq+qmYnROgHvL8jQ7sfyHEvfa0Vg7jtoSa4S
uou87zKn4UyGfH4dFh474QtP1xE32Q8TPn7JS8EMjmHc8gfDT0WJhxZvLqcysMqXcDpSr2sR8HQK
oAEGJg76pEXhQahTkV3SlbWR5x5B3GcQTdk9s2xnsaOHiham0vtKEHIE7CEUoyRJ8MN+l9Oh/n8H
9/EBPGDDIq/LeicWjln+sVPLjebUBJviTYtPtMV4Fpl79H2dhvwujjoaFGm+vZh3nWEHbVTDBFiX
oUmeuQlC3Yg6yJpQJVF5klKK/UUm6LXbhvO6NIXiKHjdapNi9LpX/TA1ZdVBmHsotyDj3HeyY4zZ
iEbSh5CExlj406U4aePKJKgMcX2GKVRkcOSUi0icHh10Ff9JiBi8f7Uo5hgcqifqMU5n42qxNEgJ
NSmyjivJOXBJ/eA1FI0sQekYb7VmeCP3zTAqZr50wroMDbWEs1q9Og1fOqgJ7qsGN1agE6i+ZpBz
c846guzcImWkb5RAiftp6iy8ZZyPyAnQwxH3ozCAIFgzkGN5QcIEn7djYjsVBRZfnNtPOZy1EWc9
vKNSsRXEg7r4/ui1QG/qlZPqN+KmfEvjFaV4W2WjzB8rjBmKb4FzYBQHKFH7FAcplu/9/qPfCoaK
KSaAgmpa5XsTEsqmKwivkBP9QsnVbIJZwss03tyI4KzL0b6veluik5IKtrx50bPsdDVliuyZZMFq
us2zML78B7VIEbNy2gbJ+jUaHHgDmV5e5m8N8BEtK+XRGNtw69k5E4BQgt/8UKzq3mgSxJrPOns4
YSg3KnZ2HrmGIFK4qpAvs/TWQue5XIloLU3kaQrV5va9Yx86Qgtq3G2hqBWVCqd2wgtCc6ho9waN
uth0WXzpEJWmqD57UKEtTqzJo8lwr7dEcOL7NrCKZ50X5mNP5+8YwuSQci7PxI8DQu6gF5vRIxuq
QcebhqjkINn/CF9Z4czVniQGCXLCUz0dH1hW36sAZhUmYDxvz8V8BWFDKysOyZSGt4Tg8wPtZsK+
ECkptCYeyM8Wb0BYL+hj80n5QJzOJb8WDS/cWQcJR2TgPc29vV+Xzn/Qqs9Y7EXXXxvJ18gtDve/
t0dWs17GlV1buz1S5zP8Yp7D/fJ+vBuBN/pmrWLPm43HwnwvLqsJGCH891zy3m8PTvSEbOibLJdL
MC3RNTi0/6L/g7uCE8W5PoxZmapMigOUgwwgAHV/xVAEcf7he0Wa6Z0V3ivkL+/QsfTKf//yYcmn
YqGLayXV9js4MW6uG1KAIwKvWd/7T9n7/8fWlRmwTGEkASe3NSpTSmxf8TD8wP8fpI+brf+zDSn5
PPfCBDWPNTQ9D2Bv8anTsMcrfqvJOez4ze2RVsPDmF2fokBRR8XenCd3Y2ySuel18z1/Wv0lST+g
Lq31+ce/gDFaRLBeX9YRh+mmJ56E3ggJhubOuBgMXyRQewpzo1QvsMo3Yn8BIA9wHa5fdqFY6s5w
UmG1Q4dYfwkhlsjEYEC+tKXpWg58D5dTeQRpSCFbAxPgOYmgbHSk7KAChORUWIB3FwYM/hq1iyRG
/6r83W8QlkscqI1dwDz2b/ksZYw/BBlSqi+dpGU5ryt8dDu9YWhUjm0Hgd834R7AQK+dnyf6+P6E
jyhAs4b8Jo+xc/Wv11RpueO26lWhTHmwv85PRfcjuKh/4PdzjBwaF+VPob7HsxAOnfvuGDMwDKpm
5jtfczT2c1X+DaXOWN8Dzgn1KYJOrzvVRpjhn4+W2zJHnoLRDsEIFXnbORtWSbq9VKtO5v4SGkeV
l3L0nh9AjZ3bGQK7G3yEIPznZ71Q+YA3w3mgaz64A8wllJ9rdrHTb6BrEhAOz6a3T309SQ+TiR5Y
YxBAcUpOKQT6TuN6hRQVky/d3PA96e47NTXK6BD0kwiLty/5JDedxLFM6eRvWSAVF/hJYTq210aI
IRXo/zDe40HyXPHfPNFJfFYX+9F+mGpnBmBJhCoCGKI37DdVXWj+biNf/adUeWVlq7qXOyo8bjDn
tUFYtkRU345zGlhcCYJJ6/K0uM2AMdeu6IXMzlxzECVfPrwMwUv9QR8fNOBaTXo34eRPhHHGp6dm
7hCH71kCb2xIsoc8+S3wQUFc5N8L2u9M+OCIDGQm5W469CFe75pNOGIgJhK54iQl1IQFkPcQPJ4z
ng1pb6HQBOpErLQXk82hDRvIIf9hP7U5Dy6BR9SF8+UI2RN5VNVQOGhn3z6j7XMC7DOGmHSP0ytJ
85GHswOj+Axvq6J63vkzOrS/7UDPjs1luO8/0lmzjCk1oGIIhAToic2tZE81G8oNSIiEceCLF/xn
mrcktodr0fdYWUagBXaiM/q7LeZIH3xCAtPaJ0c1MQnND2Apg/EeIWi7KwOmBekGNpiR2aIbXOde
oGiPHVt8/eH0hS2wolId2W0Hm4KkdHYO99uzzLjqtEg+v5HkoxUJywJtp1UMkG460OiCssKCZsXA
vXLV6lKY+GYIS6AArf7Q+/m+6YkMICxJ236LJO4y2iIWL3lRIPV5AcaqwszVC6tUjoGBdxSihFTU
rfd9J2+57Zsr3Sue2YH8/IPqLIwhqtfAiq/sUwSFQfHdaJL5APvAiTiXnHrzG9mgd+oNVGlbKbTe
uC1gDvhN1Wul5EkUccwiHOd6ahaH3KyAK8CvACVWf4izQqHOxtSxHMYY+YOGvL9z4GKXtf87yycX
GyGLHpuTzQOMuv7CU9dVr9o2UeqNA6rPnKFCpFh+13Dk40viWhCzkPyl7Kta3mFai0KLSztyI63o
QU+ENQLkUxvxnUhjcOacIUAiSPaO6AGutiUuKIRUwwNyVrlek3OSGvB9K4Q/+nHxRP8gZ+GbkckY
LDm+W5iIvuIjxeV22DuaZuNrR2WSXmHO1fgMjS1O01cSaCWemLEV83cxHhLjPdmGUw0erE2Z9UWZ
4aCCsB9Lv/A8OhzFYCoKAhkuzH+uDodAv+phBjM0AVk2dN74dpmqfPnxPbis8P/D0G1yR7gJxC5i
TRzqQGgvmkqhgnJRKZR9aThjvYFsZd72oJtf0RYB+8/oSlabIlNeknXaqrimpvuAvZFgoAbAVki6
Y9Zx9sKaoGt3QXzPaxXyMpHzZajyqd6h82fxDLKGCmzxrza42AReDU7R6SAK9j4P8p6wCZr7EG36
A7wlD0FXEfSio7ov+mVmoLeiLpdmgeK8Uyw4fqkIsW5cKL9i+ToKKY0Nmd+eoYyKAbX8T5RC2IMb
FNq2o/bxcT35+UkqvxHVVwJyX8XpViWplM+LDK9iruNFYUh5gssFDBoPWrluSRO8ZotWDCvcfFNt
Fs4HnvNSxECzj7vVW/JtwqlD8TOg0zZxl0Ev8AJF7HvsOMnGvPK5G+aXj+ILWkD1MKFm8vZvGfWd
4icqL2iVv7mkXWdw3SiZeKgg2A94e6Y3HxZzR6CZ7wv/hZ6S1GXC0RbNgGMA1eBvYzg05c0sfuQQ
R6fTSE1d6Fhwax0Fwjsjb6ehk8r84mQT2Jpzv/4Hxl803vlgsfGhUFGLPb6GKjVrj5i9JQ+RXVI7
lfhoIXetpKH39iuk4HtQfzs3i/zRr8TpSxQWKihhth0/jwjiUat732gBJqkJl2N2VQltJ8sB09Fn
GvofMfbvFvd4hrfKWURI4VR3Hnuvgg1ZWN89v1POTYoEEEG5lxQZ+0sfXKnD5Pwx4gWd3EMyCLYB
WKr0CcTGrdkvZlfLUi9bHtMRN4aQZ02Rx74iX5x7D4r/hiZwansZ7veSLsV3KhFtGaUj59dg57Bi
Dtc6T5N9V5awrf5c7fwZTYFCP2hb1OQOQyl3hWkJaNLT82RE1kTs8c8ydRHnmwPYKw6eaFd9RdIi
oNmYv4TeX2yC7n7H8YQBLqsy9YsbTJO3Ff+rr84twCNCWTcFJ3tTlkkh261R+ggbAYaPfDscC1re
A6PQl+LbgRqGFmYkGViFuy0aeCxAdpJ+441/soRimS8nXBqdt3EDAWYw7vSwU9b86QkObfW2z023
Jkz0t9/0CZo3fuA5k24Y7ennhjJEcMjdWH27OaEp42D30I9T/UZyTGgpV0qysscuGKcMltqG0LaO
/lrCj+Okg4O2keXJmWY0s3+yXw+HIjDqf/G7wgf+fEH688CvDa9/uwFj/I5oFdcYHaR+SopDXips
flsTxGtvouKxO6IQH/2CFu4HSyZ7AAuRiM+mNWz91XPZd/fm7EruMWYwpv+0TUZdOsVZQIxca3tz
/pfj+RZmekZDO6XEd83N2HQY7+Gz1Z5QxwqT/SHKDgunLsUuQwboyVLEWxnvm46LmNQtny5eXaUj
iO7wgbmgQiRhAqBgwtcKc6YsLLib1dpuS+xoTyif668Dc5BlP4ktXp7oNz3yBkuQW9xFUR/VKhaH
LPPXigp12BE+DxwG0Vttk7XM2CeO3/YCrZrKUll64OQjP8APr+eIIBsdhsy8I4lw+r8e9bQ2Pk9Y
mQpHu9tNzRYyDltiRF4GOvCemrHaacFmnAhJRuMdmkfGxwf6TXTXpW6unS18LHBjymxhjcgL+OvK
pGB3fzxcAzqRBeL2Mfu8dWQzPi12Ub1llmoCnqvgkKjrM1kfNr9o0441v5o9TzTcinAXHmZq06/q
IbqFjsEZxP1h3qYeztbtn0fr1j8bHfyxTAAjgMztoBC3FS3MGwN4gEGUoAOAktsUReoSskcaqzCA
dM6mc3kUOWKm4YwhWYj6RHj4Y6X2TesmtPv9lYWJp7pa8wNPZqCU5+3igYv4YzhiGVFMZeJF/DvL
9irHTxdctr3X+s1GT7IZ07RkeogXF2iu+5PG94lSm2TA82bVjXhpwm6tzO9DEZThdQeDzcMpxYAx
JYqVLV3Q/mX1NmP9bXDOtJskakwfQSHeOApHwnyypOpwcpBTyse/FWX+Yrn1HURFRGVfC6aFOh9u
De1U+h5Kez/qzXe915GHQwc0fB7vAKSwsLFQVMmc8HTwO9wBx7boUBmQePN8nMi7aUKXkU66EaOK
52iWzcsbz7rdkaLxZb9lBovEVVZ8MyossXfcpoTZ66IkQ/EGvi0745NBT2zAMvUZMG/KQjxcbZjR
TB4FMLVUwmM8LkPy1g4JvNVeGtqT10hT/b6tanGqtTtInliQy3jdggCIrWvI99Ar9ActlH15y237
3PeKFizscTwOL4Dv4p7+PSpFsIzDwAR8k36Ot8pTjwElKdoLooiqXdAIRq8IPqf+xYCwXxSrQKch
qnh+APBwH4aPjuF8Q6FmGvYmYgIyD1tPSt0Ze2PfrAjEi/sGHPvTdWcbcEXznp7ZMIIBl/ZINdXk
eEqOcJeBL8YAm1LYmGDU3FKlZXThe0Vo2nFEFSARV5Y3XWbNvqh243BcgbpJR+zc9twFO2TSXuZB
4HSzeYEo2x8My6AK0kUiMVWiyc5wWsxVZifeuCJ69dL14OM/nbU6F9eWG9E2fELw/TXs4d+iiYY0
TtnKvuVk96O5CjxLCjh99Syu0cJZ8LRCSWsJ56u3OzKLKkK6+aL8kJBDSoW6jZDyyNqUEkNHvWbu
87PtGaNEEZEV6s+dN3HKj9CKorez6T1kxeQG2bGM+4RH34FEBAmBqgTWjjBCxdI5a1ZyWaMIcq2z
l2b2qzRotDyDV10xaHSqOtYWRx4b7/d9AiZBhEjRixEj6T+bEmfayb4m5HzDrzqSq4pICY87qzr5
xdGDXNZ25FxAymCQ+I/wWxkJ+YfpP6qTrmIVEvvkGPKSbhfXezUeJq+QRyw6R1dGVHnv3AqHpS+8
Vd0VdFqn+CPOIQCcRzj766Q9cDL+GuKMhaZdzyb7tnKvW4yJt4bX0cvmeqhb1wRmw/7AO63hPRB7
AkEPgbqUBk0kU6Dfkr/5b7ovni/cWRuzUac86X78I94qXKTQm91aojHGcDFfioNREC7p82h0G6E5
ET+YGmHR0/KhkBBXDVSpXJYncS6pTtcuoQMVjWLqswpvk/aUNqC+irMPY//lNo+mLiXxa3u/cxHb
J25a5msQf6mcDaruh5FkTzylSfuN8E4B/3o3+cMAKDHrKzVN4b+AWgprX2tCaMtSWe+0VG5RLGTz
/jnuxqzroL1tQQiZawknZLrs7yyhmKX83kmZSM0t8Q7MCbbQ/XcjlkWTHsv/76v0TP5vMDECcQUC
9t7TVzYCiWduD/Bv8qezPQ6kQ6LEf3azsRufD4NevJ+z/1fiLqmVjloqALVn0dVQyy+gJb8eMhBp
xim2xDSUppuU6GndXfVQ4bWrMkcoCZw2Xem2MSRxUin5q5YenIYCgxL9VWvyX9wgFgHVb6SqOm88
B9hqwQjsnsexcJpdbvqywgqCBGGnF6aR+7PuN2J7EHW4dvmw/mRjDdJvwQKNd0VN+l0ZKSmIO0jp
gf/2WtHwGIylp9FxHn0Hq0R7Kr5kCfh7GTktPo9bSGs/krKJCs6Rw+TzYtzCJcHkgP/9NfGEQvCY
+IGVumq7o9E+/okiYWHSxnJiePPMGVD6sHKJczPPR1VShlXvidfsiL9HgYPpmqL9ZFlYM6U2RU/w
aUryM64auk1rmiSMfkZtjesdYFre/g7sq6wNBzaa0S8VFC6INVetaRvjLv4ZNGLUXQn1sHOXGyDA
5O+W9f3lruzHEHaZssn4dTI9nZnGlwpO+75nMzyu3faNRGovAQTknwUonXfiQ6TQLVwWfgJ0aXqT
tOfxAc2JQX2+eTzLrCGV037IIdNHqMvnD8ujymQsMjbM+L5PFjkK5pG8pSRZ45wpzCT2DPZy+Lez
YyQn+0YiV3o4pCLpXq5Kpzci+PCnkTY0+9TeyNd7MC0pYwerxUxv9jKHzK7iY/xbk/rkY3hxfxDZ
PciXz5eCTaaWBkiBsN4vkWFQefqx0YoyGKkpTB+8vNjjWJzg80lFh9xmRiu4t6D7u6gTNOia+SB4
u8p8gArAMBS6oHvPAb+Z63A4x9CKGcm0PXiHFsNcQTc8m80nMcRe2OCvoC0cb+8bAJBBMT1aXZuO
Rj89hvQMKXG1RtGetqcAruqfDkUg8euc5EMx97/VOQf1WnV1pCmYEokmVh/iFG+MXep45AbPA88G
DXyRWwdqArw53fHbEpTMWcUOkzcdUzjNDpUgUQX/djKeKqqum3catMGhSbd1B2RdKre4Lahpf+BB
Cww7fXucFayO1TJ3KfTEvhvx1UkA09A1VDJMO0m3vRz+HXf3B6DSDHDa6viEvsgFsX6ewvAPZ5Tb
zIkpRAgI+sTjPE54RJVj8Co0C5qfxr0vFseDq70+OY4SRHk9V/07IJ2urnu1SK+dnup9BQfLTlOz
TkhJwXZTOGulR3Tk3rZJJYjlx8KnEHpTmpHXjEEjmzZvQ5bJfURHySRWVUc/v8ThA+FMYtofKRbt
N0RHvav2DgDaqahMKfx74GJo09cc/FQB+80Fd+mNoGlH3nZPWSOprkRXvD2VvBw4WZrsLH4pJDwc
vwKsYKURDjyd4zPEpNtH9KgiLGAldchIyTpy3l2DRwAG69/saZHUbHyTOWAsXX+MfsP2qKjY7Qmm
NxuBiGjBKNd61GmNENP6zQF+QQ38noMn9ngM7h/f16ezwmvJXDDx2eOV5XcR3HEGieAxey9MzbUm
c0KVn+tjc5lW5jvhWPbmlP1dEc6LCPZDQ3KdoIRVY/oHtJHXG8T+KnSP9gJafnY6byKsnsaPqg9H
6DNgvWGO38GeWUk3qM/RXZA/5rt4+ajSDAr2a74zeYjkxlZDOEwWNVF0dQC2S+oXPGs5MZtfkLAB
JaW1XcC+45KtgCDOQXPU9tbgaCkLFwKSUdsywWR5eNHA3oMhzzoo4oDlxvWPRFELA3fmdLY6chjx
zMl3ymxG4dSR2q07g4M/0+16fWNMkGm3p8rLHSYmByQYxWHojLbTuQK8sQ1bRnVbSu2OoKvU7JiM
2zaUeVexi73J3HtW/ds0cxGL0UPNryj/6pJg3j1R6ri7Vpwmn9IA30kVv4Zi97gRfVPgYvR8bDL3
6fj57uMsccSP0Q+hYdYkNU9UWXiB9AkdIM+219d7+LiWlCf9PkjFoRjgy4Qh0FH7yHr+lXZhZ88E
HyUzXOF9J5eWCF7yzZVO5TEhtbgii+590xSFJodEikodlV6MU5XWj8QYICgA4qt/LVtN5DJ0mKIp
w6+pIfo/tj4S7919YNpbb6Ol6iO2RryIdTNvMHtGF7YAv3PEJrWaQeusNipK5JxpxrrQZHR35Xfp
AHL0HWwPLbuLhZD10BfRTOz7TJZECXBtv/gHX7+PdnIkAIoVLrKxfnzltmRAzgPh8+FTZW2DCwqe
SpByPseFy9feEAP/AyYQF9XnSE5VMlPvCsfFKo504qT8nek4Zo1+GzkuMZ1PeX5rIHUF6fUGoTA1
WSgVReF0HC8U30MYCPmw+vXPb9PwTsO3Kmwdk6tnT7g5wmKKxSYJ70rF00a7ucaGRn7dJBWSuZF/
UzP60oIrwwLWbMacuIVAaQezMq1kQ9fylVdBG85abGn8MNAaSC4aLayUX/3R481Fnr4KoVGtcuTS
hwBRGETXm9iTXnd6+vY0308EdR8FG0NR4OZEKiC5+3TthZiW67T53NkoHOnu17WGt921i1UBgc7g
4do8QD+PVf1vtP2T7hl3IqAZQJmV93S/KdkkpzyyQkYJA8uyE9b3/5B7zJ7LHsB/aRoDQFewgCv5
DmOFqABUo2M+jFzpYz/ERiDHc9RlLlNbce0htJQ2ALI84IyUJgNIXEZCJkkfdM/TYdLY6Vye4xUL
x6D8MobLZJk6VW33RzlA40vLE0BYKtHSw5SBQ6ImRZAPVgxtvAluy2jSfH5V8MvR+fTIv2FUKoBU
gQabTyv8k7MMkuY6jT6By9yREKYMzdqqzfoqvVLsOh0Qj/6MI79z5P7zUgd8a6+6xhpFRkirKGw5
5s169rU4AZHRZqMwcomlmHwCrsUWfqVARfrH0TCFOmviKZ8VUQ5/LuNJo4fSrf1PBFZZv2e5J5vA
7EaLBPle5mL9jj0dzKjWMYVCrZrVhaSY9eEhhFNVjnxr9bRMz9XPtt7YWxSTSIXReRnSZC1qQ32X
Y2vIhSN4Pzx4DYGa5CRsmkkTxbuayOYoFZ85LCwWSLIfyZOUM4W+xw4Q3ACamqQWquWHmIB0DIOC
kBqcGPCg7nOfgojq8JEp5RH2TKUUO9fDvTObTTtF/H3KA9asbEpBYyns5rbXJN1lketxk92uo0fw
smsDZeGD4ugrGcsvTa/3uMKKxwkD4yThv6XJhThl/vlYO9FnvGwrrFzBVp/RGLEzSyfFakQuJkz/
eZ6+bG3s3SZdjCI8MMpLi0kYMcVwk/VhLb9PMwF4870qircRQCONdMsJB//63WIJ4dMd6j/qTHUW
/I/7nXvlaxXHSnwl8GJiY9K1wW/e86kZooTOAuC0eW5RISIAWq1pYV4rS37lJc+wuYt3Ey2i511z
qxS8LHOVCWuYVZHyZbLCkewnpfPqLq/vHoFHeAkuDdW0geL/sHkfRr+H3MnG4u6xWtV+OGd61GiI
wUdcxEKCGk+yuW4jSgcDGcW3F2D3fJpOAtVLPES1l1fUMnZsuOLi0w1wPhFMpDuXQ6XFYA1kmtEG
oWzPGjJJciGnp9D74JjjGytTFJ9jCIVpOSsjLSsQFhoCmdjFRNbp3wf3bMdDsYtYAu2Koi8P7DvR
StLuE+2NWnyPpNkKqag1aMYrOZXNkiM64vI2gTMxd7kVGKNdPli0dSrs0FllHWqBl1u8lQp4vA7k
y/QuVXkiN7pgqyJ0+msrJnIixrINMaN0U3cEUSLoYDG0UdWmQXmUF+bujQ0UMqxBj8gwn5DZPJDS
WkI/DaYiohByJ39KWmjG873ngN9Ypp+jrxbcOJYiJ2T6gHBPj3yJ1O+h05dplPVkTnaKltdQvSD3
27SUa/aujGwfHdRJ6mqIKLNYJke2z7IiaAosgSfFJotLVUveKE/ucfWOc/ZMRyu2sLNG1UEIDipH
8wg0N+QdZ6j28T7+UvpD8e/APkrjargl/ghhxugJVHQPHHiWLnr6vIZqN3FPWTebpbxVm72R0JFy
cD+c/6mpzK7jcRACqiP/A2TA1dA7nNnaU7b+wlxSYytFvIZzac7Whrc6rbIUw5J2T+KnSas0Ohi0
4f1yuc+ZEtEFQUNqw7ZyRfRx0zRiziF6xIo4UB90iO3LaEs7CqJHuRmd0XIzGXPsJkdUh7O3Y8g7
YZzJYVo2SmqCt11492GJxEmnY84dK5VEYt52jzCllTJVaXb1nQs/2Af3vV10M4wTK8Isvi/f9vMp
rDbkA4tMRMFfpTgta+FUsV9q+Gen+jE7aB3SoWxH3dByKplKFheACFUmsX15y+c/dKBw8CpmZfLP
cVGqHIH/ulUomMq5Jpr3oXqVkfcD9DmWvKIDhQG0TPnVrtw+lJo/y8OOk0g1+hiPbhcQNj9Ntpby
3KS0yWkAjltdwq/OlPWg0dNmaCI1cn4hiXNGbxi2DvTwgT6AOYLJKofTdmQg5Mr0Glo9GTSOcIye
mDVGejPkuReWNPkdHCfkmLwyjyTX31yP3A6gz5XMdr6NWoT8GO6zyGhvoTbzuDrWxgGmlkyQwOHn
KeujVnFFemODnvSP375W6S9zq0Fg7ay8GJOpdLeV313LPyEIGYaEcao5nKTEsrlSx8GyF8D72SK4
82ErkX0Y79O85OiY0OHzN+CeoP3zrt51j8u7k4UyjHs2kzGmq82KY11E1qPmao14CpuKH0fI381s
l2ZY3vR0BqINkGjBiQnvyPJ8a9663EMtO1cMndnJHOVmFvkNXUQEbqVQo41okgGkdmjFq0sOu6Px
MIIfWXIjKpN4g7fKL3vT3ZgFYrfiUTm17FKCY1GlosPKj8CG+UvOnt+14bPy6qL6m8BIoqmKIYSq
R5dO/PHeKGr8h7Ts7g7Na8u9NQeXeurDa2iJzOhKr9+S9y/Po9s78CUAqwCJvPrAgw9jsg2d2GDA
alt9Lryq6zw0OiqXcB7xvJaZcE5hpfABZHH37GmQ3Fa6JGm8xJTLhTtrhlFK26fqud0NfD5EvCy9
T0h5V0XdpKw6c3CMAhyARY24whDrmG02DEsXONnYVFxB+TJXyATGv5HoXGFVJ6xY9zVYKRmzjT1P
DEqh+4GWScbF7Bmo9jv7bUYmueS9Lp/syeNxab9riCVoaIlB+YnJLRsmYqiIozLf/0BeivXAJ9HS
CFAorVirKnggqYaRAu6kDni/2Lzkb2ubdZmU72xZFP4Tptki/B4pAdsAkVg3mGWkwWsUnaCOgttJ
9z7se/jmQSUfxd/+n79aCtCxBBY+Oz0L1rlYVuzCMdZ/7p6L/WF6eNrob1E1wKSVEeoBAuSc1vDt
yYb5C7i8ArRtqtS0j8ngCWtpXW+XObk9V1pH2Elc5f8v3Wvk2ivNNkbRfj2x+axpQKtOnVPXhVqN
BWXzEFVlDBvX80lIFovKTY+jGD6Esls/5i9GaSkyzhcJITLQQpRAAyWyPi3yfwAfyK1QkKHO0Pu/
c1UyrZaNzRohNH0w+bfkLcC2jjwmIiVnRPz9skVXqJgMtZ7SRrKSpXxBctqTQKP6wUhrqsy/8xdg
JbmOzkl6cpPrLagxXbYfxR4qoGLXTdFKkW4TEDgbu7noy0+88KUQs9YazfpxF1wgV5iL3pCZG6bQ
hNkjcxp1A8oLlNHU/N8tYd5O6sBPGusVXy3YtMp11nIADmbMWYfzwb4+rm3qsURvU+qOVbFpE/qd
ZEiZgdHCyO3njoMRXciQ61SIiAaSj9ctL6oDeTcZAFaYYk7xIswCI8METKuw2D9gJcSir9VKleFO
30BqHhO9b57MUVhrPFrEsba78bxH3rgd499TDwvvo12B/b8O0YwMVEM0J8PR5WxPSjtseDis7mYM
0EKtLbd8NmF/Z3OQbVF/8l/JvFYX5Etd0CifXaXUtkQqlG0Nk6SivLuPAjMqrWagQ0MOegs0jCvS
yUT3KSTIm9492Ar6IZCajjdGPYh8OtKyZUg0bg+B74+9Sr72k1JyHY/jlheL90Iz7Alq2eQ0bZBI
hyj5/BcJtAWz/VmS+0r2OE3byG2XR9+3M9olwVxtywyA2ZaMkqh9usoImhXTpVCWC2UbZYsYaLov
xwBb1qZ8VnBcWx7vpe9+zKlEXqwKDedJOD3Zm7SDxxyKGOXCICnCqg6mYsz+/rkb1GbJ3/POzXZr
CwQxQuI+UgbHbevrKeVTYqRgEtzsDGCgUB4Lj0HAJqarrUv3v9spjziO2GuspaXn4KWnl6cBSRJz
IXqeAqNneywvr1lgaEtAB+5yTcaOobjoMjXBWm3j7kOCWbxTRDCv+TisO8ICqdTIWYm8rDjcsBoa
KZ6omzpKYAWbQ1okNPe0f7xyNt0N6N7NaC+pbfM+9Dtj3jnfWMKKRO9EViF0zILKwyoYPVG4GEj3
75gzf9wXE7T6R1aRQ3+7UOX+hrwWLq7HzayKnQAxnlu8mvbpDWMEqgK7qQoH1ko8HmBfhIm2qQSJ
wTAKQOg22231bMqhv0pDW6dGpt5pky1ZG26wPEpwNUJfMDOZxBpovr0wMXJuRLlU3LurvHyagq34
gtXtW2B1fDdnQaTH7v+QHNigGfNK30K7ymUKQi7JRVpmn/k5EHzcwHoTpC506fIxOSxejxuan4bS
Ft6D9CiDnLMPEpISicde06ZKlP5Ra2QnJXc4E+rmvkluAZp1mg8YUr8zJzi81SSZRFiJXOGgyeS8
fLMeAiqxLWwGgYxpPte3ZBOuenlvYwnii5ZZZvbQI1Qtx/ICVRyDsKJlkC4+FIhLrkOANvxB0NAQ
AF2MbRrgAD+6Wt4y50X44BDH8vEa4iEIyjsVoJazlLs/ZS3Fe4K84YkWTxH6Qgav5ew8L9klWSNg
DzBV22AqhLkxe4DE5gPbkF1ntMJiwDcqNCblyxOlH+gdaykM8KkvXdSPHto04iKF5NHIgAhR6B9Y
lHXWfYkbdIBjvKmqOHgAYPR/rxx4PiVJM6qp17EC36wpcddv8n/fLpbj2zbBAe5f35T86zPXj7AB
IgQPUDcMKk4rMrg+s9jhRM/VfFrvWzS8ywESWUcly9zXESIni/0M+4llc8z8ar5/yv/W5iOgo+23
KJO1fMMtvKcz8R7j+8BUQM0g2KBPE7v4MIQDJvYMEi4NqjFLp9OvZ6fFHBLwqreqliFKE3VA2uz4
tV2brOoczPOCNogIM7xAtRQcKbQzfVf34A7gGFC2yYziB2fPZIwDjezsKVOw5fBrrkIi6szNWtR9
5xI79qc8Op7Vu2kXfJQoBfDL8MrQDSn9t/UNUYUdD/3riHiffFTmQgIy4YXqOtUTNMvH3YGQiHTo
6UpNW8HymDt28AnQn76JCoMRUD9Vqelv+YOcpowXNKnjAB4BG12Oo8N9j/HDyhbpR+FmIQ8eTHax
6ScHYZVz2PIR+repxeLkEiWR/cK4is0UFImNjcrpMBp14SuHr4IagGoOye1bJUSIH9xW/WPk4Ts0
HTmqXxqb7zvB5cn+nsZHqIRLczSj6pXPsnyWr+nXAbSe37UWYyHp9uDZH4NgMWbbnAJ1f4ww7ET3
hwTNDbS1msHnwmoHw6WCAOlVcIHCFw/T2sqHJmAgl0v6NpRgM1kVOzDY8AztgUPaInSoE3n+1Kg0
zLqWXG3EXnamYg6H/wGFsU/ICUHKo+stkQbQV/6IZPrqu5sh3WMb/cmI1aM+aynnRoTlhfhWXy4T
UXXOeP5eOKuEb/8p9Wf01BUGXl5XbaJsDcXiSAYd6eA18uH6HZvBG2+p84qtWvVfL+idYekNNClc
onZ6ooHlnvy571nS4FyxL3Had20GZhzIwj3x0c05UonkZMgn9vBb2IsTWsJFAb05NR9RvG6d6f8u
AcYHBkTdmXSSl78R2ixl7pKei1zso8Sbzdx1Dw09gLjkUIoEfWv3bImvie8I6wBG9KG5LxEaHI2r
HA6iM/K1kB1CyD5Higx9YeQmZ4C/Vt6WZiV+WWYe+AKKJlejQFiyWzTnwpzBWmQnXl86Jxqk8KXn
CiZ9oHbohN1PzxMK2wQyLOpuODnqQnTmn14OxcDltv3vQnVEIOXj4IpaUMnzCspZ+jImvrElEAMO
Vw2uJuiJWJT8iqRw/c7nM59ex0QdBuXSEHMoSlD30y+rDmzC5aFAjxxPNLFrX23cy9GXjpmattu5
3sjx+gzljG2S1zAWmNY9lTsg0RYu5r3FJI47dVmOqci5cOpT6X3rsvhJfban398kC4lQVc//Q9kj
fdI2Yh/6sG5CYK7cUA+RrxXlhCu72zAOwV8ZvkHskZ+eM8nTTepQvFuQYiUlZCiuDH6VfszaPkmI
4gbBV77Cs2jKUFN890IFxGygCkqZFVcf/5bm5JDqTlchao+xcIxCUbSfPYh1PBM6jCzni4lbhWeJ
Lkz+TT+LAJ7jZ4lBUSkSph14MGoTGSa/DhFiL6Pk4foCIp2tMV1JVrUgWMpCLYPipDqxIbJOtKRt
F0HO6H5SHMNOoxN+CzXQZBTexUE74O459Y9bO5c3pGz3f0ty0HV6rR2ZbuvZePF383/o0M9UR6o7
rGYFst0B6s/qw/jmOlMUiWwt0JGzUkackniG33YC1kbUUM49QDUUnXp6gDzH4P4rYqfXs7scABSu
FJVz4CNOpn5YSypUSXVDS3S5wKHGL8vZC4vWLZ3lpie89nDYF/uoJ5b4nG/l53K4nPGaHoLeR7rJ
NJy8VMmF1k5Bc1V8G8dVmSnrhJ8UNgiNCKdYvPZAuGXyY8uELvNLMS8mb+3GkuX86avrhcRGgpRQ
KpBAiOxC3IP1de7H6PqL3nHWULP2vVyLgsR+UT8zXb/2zjxPnDlBZk/LfQeOOtfzLq3dlD8aSoux
ct8qS7qeQIWYFAbA0z9dDVGEbVXCbKd4CtHiMGLATwRBBMfAOKyg6Q4YVrrrGzln7fRyKCjTVbRF
kKfM2pP/k34Ds/Udrii26CGUEsxLWXS6Gq4Ey/7Pdr2zrVxAJz5jVEDEanK6H9tZwxeXP5uXEVvm
/XlhO573dPAaFdeDoCXCp5exIdH+4vH761buC11CRFK28XyCInSAqKHtQWix/TdKGoCemDcbrBIz
vXRZhytbBrbV+vQYRTHFQWmNjBv4933e0UVI/h6cNNDMqCQgGIsEotbh9wzVyRy+katk0MSHbGDT
VIlkK/GgQubgJeroNzLC/fVQlzAsYcE9fe+k/d5I8bZNpvytk5FAL0TUSglElGsyliFhDpH/bZJ/
M2I4RRhPMdjlmZmpnvqrMuv88hJKF/Hutt9VK7MePKKO0s78G6K9/rZnHEyk8aaeFJlQ7ObBz2a9
+b6wrMgcOp2Xux4sFJrU0OLALD/sJLy0jiH9Fb5smNTxpCLj7zSXvBBgJoYTe6PyQW52tNczn+u2
n46q2FRTpEj2DcpN5l3StqJE3j88/sih17g0bXJyx+7tR8QFaFLAWmmo7vGFlv1r9RMHQ/4xEtND
JWIe7d/FqrYOSKM362a9hBBGXNlMT4ey4jJ0RIPX8YX+CAEBBM/qyVTeIUoWCerC66Nu+8LdiC0l
L9NWOCH2W+sZdHGaa9zXgnIc7p3WX/c16Pc95RilW7HDIPzHADVno4J8v7px35XRcpv+y0kXi1sP
ovJuxzVkNtLUVUMgkD2cSLGy69bjWq/bOlBkQZFWpq/Mt2+M0HxfGHPzxEvnIOJ6lUUrFfh+Bmhf
vZmIBe4hmBBhJJz26KTbaFRcxwzwu4f274IftsNE5l7f0pBTxKEA4UPCOeWlYQFgQjwCNxAj9Dj6
7b24MsZmn4YRGGYe+VsQO/jwJv+l0NI7hA9LWmPTnibsIi2pypyOGCfUUrJI69dAROJX1NwBVFPU
rnn2fliCQvmi2hn+kvikZoBVyr3BLYFTLRJYrKrVrju1qcQJKhwtyMB4bf6OEdfLkpkU1tfgR3J3
AIk2oZDLgAfCfOu9J+TynKblEteixwZzwveQYWK5TkWu0fy9gB1H999ptGRRnkiZgZ1Br3wF7ThJ
EnxWEWFTVeB1giYZvxG+G1RMf7X3OEA3CdnltWtNlJ7RLlgJrLaMjAve0ve9c7g0Yjg9L69AcabP
SujGqm9kCED914yt99pwcxDovziRNaZh788oxTZ/9sB2yyR+EAb7E90KVVaHQMk2xIpAtZ6em2zP
OPdVxT2CeEht8BX+OdMaUBkE2lg5kjsgrkuDVguvhwmH5V7K1b4W0sx7rzgz2t1P8PHIP+sDQv5g
Xk+dvl28k7Kc/+kxfH9mTtRBe2yWetjAWJapOrcb3462upTZ5rhPfq27mPRTiFh0F8FPjH9+cU4d
DcPbElw7eAOyKt65xYk7tvEcp4Dt2sqhCHsFCBdUvm0aQjEwzqkhKb60arl3Pt81cpcHzgewZ1Q5
zqm28p8b7TwcGARF+UZNnxepaRUJzvEb9yeDrKGluosuoQWNYHT9+DQLylBZSbtTgcT10Qg0Z2+r
SIOQOYC7pO++lQUxk9ln8L/UMeCRx7DFwl2ELvY1LAJqn1runnnT9tKlR86aAL5R+HVQFTrjVZvd
ABCebIQIPNwK44JiStcQRW4VGqdGxIIEaxNQOniNWrT9OsgNoygajeIjMqq0kfa8Bc3fhYbcTnbA
5H2ud2oR3hgGJwfCbtemYD4qEgCD44vUUmdgyoyRvL753StDU4+J6Rpgm+FLYrwynUn1Bo47+mVm
Tio4nGVGzpMe/5CFfxnO5IN52FRNcbsIllh00/rqZRXKI9Umyio1DLrqp35yK2zAcblxS09OeTbL
UJFKQjE3edbGhfwZ2b133a8mUzXVuVHDRQj2eLxDpYOedj04UjhubAYZJcgi6TQYcHv9wV8VQGov
Dq81Kfc2WdzytR5KfO/+VWbymXbWTFt9zpJgWJbKw2kPh7Qo+5QuCwAq1tOQK2E3xX815INW1p66
wlLhG3jE2GcXpKnchZUc96LjVZKr0LBhCZ/ZxYoAAG2xQcxN+2NN7XjirofNUCNOvDq/FBand6YB
fQmIi8a5ccgji4UYbSaXgzIUFqFqr4TQ4HINcyue276+NfcD98xwu4Z+aPKNlZftOcHd0Ixp/fWb
O1GS2nl9f8oDj5Nb/uZLch9sIqiExUMvrC3htlVQ9JYuM+zzyuKTxB9/U23+y3mU+sUGJ1rzt387
u8m3dNVI4NL3X5QI7CyGCSMSOAo1Fx83JDVCkZv09ZG0S4IbT4e3YQ9zakYbW9eXCdsolNofDKYZ
PQXevPt/7fIqxodBnGHIQwN3cK4FTMRjXDrOZ7qel6Em/NORnVtN+fNzeqtyVieVR0rMrUrYOxCC
/hsTk2+V11TFME1MyRz1lK35nnjkTqM0/Zb2Ls9w9B0ELlKm1y+0JKW1HpmbbE675hzTLJmFcgC2
bdM6XBjtaqFbP5gTCvgkJXiUnN7+olXdBszIP96klFcAlb4HpEQCuYiK/atKZRoNJASdH3Zfxnqk
UfbgN3RKo+4DsxqMCIGygRNQ0QY1K6aE/cPO6VKh3cEJwnjvyKFuhUzYBr3ifAokukRdepeLG347
4g2gHxLsx0rPMzE5+u9cvTtKlO1Oi3KcpsnAMPnhb5T6kt7GRGbJnjk24hfsBTeK/v8NcZQdOgQe
mGSHF62afC5hJj9KK81r/BM4C3YrLU+fCmwcg8o7R6MsOLdb275Nz469AkzP/YPUxoPTMwE1QCY1
g3jzeq0tSQ8XQ8E8kuIxuNf6LwXe6S0M5HDfugVpZek7pqsXz92wHD3tSUxadxHjsjEbNmA1sGPn
poTnEGiQHcHPI/XyonfkXlB5vaEAYv9YvLCyrFfTuekpO3I29QaiMbGlGsn38WBMRkn11lntptNA
hy9EyS+RsvQgcEgKJxCocdddB8fkEnCuo/2XJlbC0MJQQaNfKETaYuR+G1ilEcO5VX/JMtLv3zQL
xdjl9VKbIwdl8489qn+ybvRQPPGcRrNccOh8/0RGgMeajM33yDqYA00g0EEUvA02x8MO8tnSO0Bb
ifA3FbZ9WEYlrTXXiamxtNFbqghgNfDVtC1AyCqEUmTuYD5iXsS7kuD7/HirKnF0gaE4PyOFxJ7n
TLKd1P415YCZmr81D9RvB1R4Bn8zt79mSgDqfj8FF6ZGN/X1canj83gMM0TckiBQ2osWhgWd7/q1
AuVIAZLLFgPpbaQgHqmL5kmsYXKDQxvOh4wXBahnPvsKe1f1hQDHbIh0NCmRR5Bk1S5NihaQjV+L
q0SSZU8IhQWPTstZlw4Uw3tJH5AZHZGsibmmg3j6J6HHXLVeKJwFSIKvWbKrHn83WK25XwuUD6Fi
MVC7iiSI7BhlUzhuWf2LiVrAxl9MGIngIIodncFB7BQnXLdgox5dOQfJgTBEcl00ZMXT3ko1OzPA
aGr6Heofg694qY2SDaUrLSqhpuPJl3i8H52N/l7iP62TK/Gak0f8iYrSQwZU6TVQMc5pRZvPB8vM
fOKif2a92uD7yZzzPq2P84ZH9kgzCN1DqgPari3sSes79sEXoDE4kr+AeQ0D+u0LjmKcLHwRYC6A
z6aPqNujMNmgK+BQ1uGUh35ylOe7QQE2by24FmAx6Pd1yEy9Saqt2KdbjyyF6sZmRDp88C5KZE22
Xj2LIU6Z1s2vTXwdT4oSYY6n98Hud5c88TKTyeZcyBKcGMqQd5FMqd1FAQvQzcTOZPpekdw2Ph6y
1h3X8i6O9DLLisIf/fVxGieTgEe2nj6qzuHVMH0TvjryzcHRX08hm9aouADke3Mi0HOseR1lzU/1
RMN+a85G0lfinqJ22m+xSOCaToZ53Q8ZYg5rmQYr7uyg/ok2WtBTRvp+VWJ8YVvZzYinTc0Snf7n
GVXw2uCRPQ8OeICM08MCQdsXsFG8GymdCzfpMPTjatAkZigutLp1xvrdwKkiSeUkc37i5+dB5Y2i
7F+BbPrbP9JMpm5yIu4T8Rshz6NRpaxoXwZGbcUpqA+EWjHn4JKalr60CQkfbbmG80rOZGIcGYk/
UEguczhxniLBXh+apXVLJJYouEx4POvqO8mUpRFc8x2XUsdlB5I1kLT7aidYK2eWwOVJvprvj0MN
V5SCXqYBLTtttt5BBpHeN2cJloq5dmGfxAmzFZKRI8RnVjmCAS9WJdFISoFFa638bgEG5xUl+DpP
jWESUU9gNEstFnRlWtyLx+ZJ8QdR4zrqX/cVp43Bt2Ge/8dIi52Sj293DU6eb5Dht91LPWO34qZ0
B1xEF98MxFb8DA8aX5ZekxhJCd7Kx8494DOYJhv14nQ9xr+pUsA6p+2KamjIQ1Z5wTwkZ+QJqq9u
PTpFWPJ1ckC2Vdj004IvHQJnUrLFbTbKshzjPH20Vu7zxqX/oE+0LDZl6qSykcUjjPnjdvv4LnKg
Sr0bq0+VnHKNun1xb9cA9P56E8cWp+jSPPjC6Aty0NGy3iMxW/LiIJFpHgcwROL0rpPqJkhC0Hw/
W0FguDXEPDQ73yPlB7xPlz/V8EMBIo/c3Mk1Enwo9epog6sown+ctyHn5HvFDMbou7ZHL+3mMCHO
GqaqQJJOU+4fKso5NzfnYGexNdsRPowgz4MRajG2QCOI5PNEsEIX9hPvfI8CWBfedWp3KvHskaJi
ojGh+pIANHcU8bjcDvQJgEPaSHkLjMMGxvul12ouFNmzCTmqe4g/C8VXXY/4tXTgGog5QxmuGX1M
LlYOXR5yaYuKtYyPeNeAA0SOEz/92twK6GGij/bC/iO27i172S9I7TnqwRQcQ0r7Sbq/JPlFQYxD
LQ4zcb+rVletDd3xuet5OEnHaKhb2DjBovZJmd0mC9ul4ttbb2AYBc3iuD8ddP68nEZEjVOSSB06
AeAKt5Q9dNj4BszqESg4kZodXQqyTtQQvab0a80ergNUSqQZJ3qMJyxj01OUkwZ2u85NyNFCYDfq
5qlV6KxqUhKLFxNIBjyHXlbzsD5mKWN52jsSZIvSCIU4bcvETtTAMI7s7BYYC5C5D3/tapzyzaS8
XOOtBpXWzu2rnRovwz49hv0NViN53V36jVCs5wr4Dbz1cs9mKd6OVfSdS2qgY83h2a7gdorgqEa2
1OcHI+NRiBEKxoB8ffb3i4dU4SPuzg+YfI2Q45cxi0yE0fe3rIaDU+YqUySHpBs7iqNx4XZ9EhTz
JLsFrmegu1xqsxHGPBhCNGsWVbKwsWy0eUPB6dpQ9Zf9aXqPUE6qnOE4pE/sAWxe2rvTM98WfbR9
8q9rqMwOXpLu3FOoSH2acvx4vEaf9RpE1woZQfF6z5hzi/KJ4wgkrsIxT4qKHXL2NjOCoaaZUptZ
GoGbK2yM6sxtjDE95lDSo+/mWnOeJUvQKbx1qo5XirDOpB+S725fSqY6U9153vdrvHeuplz9DzbI
BiQmVGuX2BW7mpDaM8Fx7Fh7zyz3BIc7GWvhStsMxvpYjRZiPU5EZi5R6EDgc31axbUf5SsCeyqN
S06PL18STbBUIwdU9lQwOaF9zxfKDpuPPQjBrykR67rYkB4AbGOuViJjlry3xkUNh6JNHjghO9lh
y6Ud4jeQcNJ0tzBormmAbXCMLBkoGfBwY3kpqw5re9g1IgnA7uYs+sC3Udlh26yLNx1s9TjUoOTt
REQpWYyqztP0d010hsNKwikVUCajhuNiK0WB5oD5m9QJNMALKvLbkRrLZocX5D+QXNure6BB3ydU
nE2sbdt33PI6vfX7iik1sV2jBU7sa53+YtPukbV/Lc7/ZRUekZ5Zd2pEUB+iHUJ777DFti36X6Me
oX6dH0NF2xEryU/P9B2lRFrk2TDPB85Lj+7i/PtA9j5YKswaWnI/w+IoGKlXGwGBabOLMHZGVnLZ
2USfY/la/lK0uwGEbxhAQUJxlrUzYo7tdhjBMYxtGGPI2afuRAzTg9K4Wv2kJlaeYKUqXDd0gJLS
RSkJJe4rfK1QgIX+rEswuMWAw6ard/LmiMiuuTzALGIOZh3CYwunbpjOuhf4VsJLXJw3APSMmSeK
lAx/Jh9A0kiMANbXQocACB+ubzqvJ/MQ69XhAgnltFBVtVhHwn+/vwreLKmADMD8AwS+TRk9Yw5e
opxVTspEw9yFFJSi7u7oMa1i4yWIj+Vfgbx0O8qhGMGKjvWZIpebWwrrawWy3GTjGKIfkpxvJ/3+
fCDyt1z0YYy2TVvSTykW6B5JzHbFMVFkd6qP6++21nWTta2gQJf3FTqgix6cS4M8rlgI+092Q1d7
eRJJwlDjzWjmG9MeBhKzH6MvmLqFGbm4XAmJG0JP5TVZc1xXjfYFRmgx9Tv3iHQYoUv2HRbHud0I
s6z1glLe3jKaLeV+Ua4BuFFbUypv11C+PbkOibjp1gEuQAiHB5C2sKed1OIsZW+qXQYg3Gl8k/ee
bT9KDPwMmGkb2nQpQQdT3xgxYt8E4WtvjwLDJWU2pO99WuPtb1JTtj0ZWUMVNqYT2XW7YkGzqzLJ
vy0EOlcFjL1CetDR9a8XgcphpWr4Mze+gmfCRJEgwOVfvRa2lJDGeQw/2duiu2uHcNFAj9Z9mMJp
EgNx/NHBa9A3VRjeNnWpW1KYSbUukkr/qWiy7kEpXyJSNgh3rX6nlH8p3zKZzrluGyL9YjOF9v5F
5WR2J3xtG62r5F0Q541AJbsC0YeRCKrHv0ixm+VaB3JUdNH0tLRXGLpPAQn41otjkpTyqU32TFKq
aWcKD89FphzJcj7M3nb9b4DNrjcAXmK7YEmH74FSxOV2PpCk//ZsZOXjlMk7w6XRVrmQ4a7mvc38
14u2MXcq/lyl1mnJiRUOmn/RtCXU4jHnkPu743Zn4gj6qvu3SUZn1eCC9I4lOkpJE+pxyrCsZGI3
CfX5A3Xb+cLwr1aYVUmwDDND0xIoz2rudCmnlw6Y9Ld4L3DAX+5jkz4K2VdiuIy0GcJzrfiZqRna
Y4SpA5eucRWelsw5t+zeS8AXvxh8BkoDoZth+9iFLXEguYF0wUFy+4Mk19w43KWLhJpKx9CEGG98
FAkTzWkMCn8Mr1hzSo0D+9fQjgpJ/NMJO6LI7fo4rynE6WT5k+94Uo1/N8DcDUyaYhOdO3yywP9E
IFOsyb7G+JBSaCLMyv+XfswgDmUJJto4Klo+t36Q4buWAnDQy2qOqcek0EpI9pUYlZxAHm+5yNXW
+j0DWzzLv01H2zufCsVza7sKFScOfutyPNd0jb5isdcX0gcQ4VsY2JZSK1lAFFjyQR2M0m1z4Mt7
QqHKv40Ezb+PyEY3UIBVxq4xJcuobuHEq71ac6P7AHzqEdnMD2cyX9G1L9rpf13hyM/9G79Fr6iv
7DvRc1OTPc8thAvI0t+rRVD/HZbrYdXqkS0b/BE8gDCNluESIPg9R5PaSLw3Pml35Zp+OVpwcmVM
HK0/1i4h9MKXWwwN76q8QZIfWpQcaiHK2RnLGGhh+/QBW+OEuAG8fOtw1nbIPVQbDfrRDhsYX44V
EPsGJYkJ2cwGgWt7EH6A5h8jwVGR93/V2/V4josmApKcBfr1NtVe77GkusndPjnnI+/3lDJHJP9m
Krt6IP0qNcpGO9Zrvk6hlCQKAQ0xyiYvO/UoSA5oKyPzzv+sPXWqHv+mNmQLFe9LQjdJ877FKmY1
l1GReZNtmMJOjj6TFn7Y3fLK99bFJyf32S7IyhiL7f+sxNOSlo4iGuonUWS4EP5Zo7IaJjPqKEnJ
gEyNNsm/9tlqR2/J8/EH4QxciPsrKFbdULzCUt5Ge8yoNJAM9b391ULEZaHG+odWuu5lJmNmVJET
IjLiznj2FmwWufnqb0lflEtlVXv35Sw0dn3ugj2rho7FStxyPyU/Cn8j4onLn2/mf3Loy+K8o5/F
SmYuvRdu9DqV45mw+uz2aVq/PHWakY3jiEMIjBuM07bTJS8w1IdWrV4Znyjb4a5xRjAyxFd/aA1X
3SIdUmGcstiycigJ+9WzZp/9sf6og1YbQdhRq+R8W5BSv88w0alJWiSLHGOaq99zeuqUD5w5kf7K
6XImZUAvZZYU9DGowcNgmZR49fg4/m0daOEQBqsw/eghExF2PmvqFkHiQNGBJah3G1RHAx604WDM
FMNBAhFxpX1OpAsFNZHkmpKXsoaNgDFtsmw741bKrWrGlF2XYRH1sWMPB0+4EResOmVZER4npNKS
H4iiNN2FVWbQ4Mew/9uXV46whNsR1nkuqLBAvfig0YApuuYTUo467+Mo3SEbIRcr9s1hUHC+NaS0
TIN6hSm9MXCMTp4JdfncNWYmVElCG1x60MqyenN7L5VyUKUq8mXzDuDPEnA4TguHF1V5nvdmbZQi
ADSCv7w2xDse81/QPmQnkpewJZnYpCDBawIrVtnsl3m2a2+PXca1m5J6LNdIbreuGZyBUbYsXHyL
i8RwHs7aJY8xgwpk4t0eOZbPfClJbNaUsc7xn7EE89yOUOjaiokpugkkPFX8ZBi4DygTbvM27YAu
fbbe+2gSXtdJF9Rd39nKdQUcOBRRhYezrjLHobdj2cWZs0/BO5noBKDKbEeAKxiJfiQC80jjnGMy
2Gzt54bhgGNY7rG5WKoI2Ik+pZQJEGYd1dtVtkJCSLWBGVBeGGJDjkLx2Buc06nXPlla6ebLBHTT
0wJxlocrBJ3Z+y1AKWep155r3UCQWgX8Ir2iqinKuX10Y42GDUe9wRMCANz2S4SKHm8Kzz3WEvmz
5KE0/VuZX4kwkGFgqNNjsR2BWK+gR0SdGYNwOnHzHaSNN0/TD54VWAgx3qy7F7hzz6dp3sBEtjXb
f1VNFnavpBCKClvi3LXjHDlDYoNojaAzSHfF2GqJrmB/5tCuqu7IRs87vHrLaICd09q5iT952OBR
fRPfr2ylv+AOSn4wnA9bQjfQbii0OqhBmsR+QfBIo/xA7xQ0hIBDRgsDPsZuKDnBmPHEWF43ukwE
xnQN6LnmAdfWzM9MFQ8MoKCqu6/qblYER2i6F7IXzrrYYNV9ZVC1KYmMyJbUINDGVLsMgy3BREvP
RLwDT2X/gcdwFYZZKjGyx5qJOGi2zz8PQmiinVuGAn4tbAF0GXmKtZQ1ie2eQlPyGx5kbO+ImMcK
0sITfn6E8yb+27xzi6LtuNCgpGmUFYGE4B2KncP5rPkewFWwFP4xFDib2OqWBazG8Yq5x7d2nfdC
xBWeFKbEnPiKdiPMfnd+gqho834N6Ivl+d4X5A30Ks5R6aoiN5TkbWCNViptkV9bYjeXOnz+CMZU
pLkHGrBJArK6ry+h0cpyekEAbQEtWJpLy+RChxrUv6V3nvl2fQkc81cQdDIfI7WYO0wQl46gCo/e
DjWaeH+JP639lqN+p4ALWSCAGlEDYvaVYlveH1W2m4ZUlypf0CL84K9cvK6pfDcHygTwyYvBFbPA
2ctz7FyQnTCduRn95xBjFLZ5pmISF0Be2crmFZBnJV2oCDlX/00nz1qsg16RppgrnA09dE2pOWGh
4//Q27SlyDeX9PvBkm7xj0Def11cjd8s2wxfja/YXsOt/H4SyWoTQ91hlRyqbtdCK9HtlFzDLMSa
gwHvGJIRJFtsZ8QTTECLsjzmm66xJRTE17tI/GPbt9HmWU5eZ4H9MxIPvi1NKyXavsNkAWSe8OUV
Ycl4pYzj0qvvw/Kl0eaXlzDNwd2xBwU39Oko3dlg+H00krvULOu+boZq00LWUv2YnePi473OPvis
sT7O6Z1J98uGXkIjtaKMfudOEbjy27NX9Ek1J26hYMLhVyGH2D3jZVuYYwzGJluNbfJ+g+XQQK8l
UEECSZdlplNZoTYU5usBcUFzFuAUkyyLFMH8+DHDry3zbWMEF4OlqAl4bDmdcfS++lc/l3d1Lsbb
gZ/JuVaHg5hmxs5ITwv2YkG+Ra8PQf2cjGI+ZnImcRhZoGvocfaReEOPuNZr4RlOLxIwOplqlYyL
LOewZlOxejWMPyz3FUm05lHd6ii1zCaChqzhDr5Pel5SoE6mOd4hgRovoyqpSOKvuF0C2lPIgU+3
cmka331yAPuuKawk+7IA/BdJGoRrj0ixteJZ9B3g+JOrq0kKwPsraJH5rbLgOLDINYj/NP6cOViC
ZBLx1T77CPdwLZSxh5bDQAg9fnIeMWGoGhVNibXaTf05NEQQYxQTFa8xoWK+8L/NumzlTp7EH7Bi
ChILbd+0E5OtLzSD/u9rOJTR/4JAEgcDuy9ba2VZCyXpaE9hvgClK2GWb3AL1rHIzeo53tZwi9r+
xcpri9FMfLbaSXH7bkUmGUJ8HuPyTzmUfAgGVyp854MWg9e9hKOhQL80RK5ERGbVfekVTOoVXcGO
eqUK5L0pK7x+uwSyPcGmLHlgTB51hrYcVoNyjHn7UkJk4QAydJRx+iUeB7lEf7Jn/DjAWLQQ1nqq
BK8+BaDFSkLs0BX7U8y1/Eh5dwlxpLCLwYDSOrORK7GsOgJOFGQm+MN3M49LaPEdwu5Gj3+98s7B
S53pJwo38k61sbSUO0K4TWetb9KDN0PHpbkiGi+5XcUO9367t8JlKJnLynLkbixc20zfh59109Yc
Rw+jbSnuOEMV7wOCgrvluholYJTsoquPGqYWIVs3wwW+CPxUTS+0qJe00k0JveR/fgGO5LPk6LDC
CuuSwahY4sst1llws2vre1h/jxM+bbzJNUYkodv+Glw9luDr7IVRL0G/r/O1z5UOaO6JBo92QXRa
bQ6+0Pehbp0DTU+vkdOyidg2edOHr0j+6aXp1OVWiuWOdhB2Ltfgi3MQVZyDOBbfjqASiyfzMnL3
7U5xTunxMVKMbCBjQzY20uz03vxjBuLLGS4B7eKK5eJ7pduqwbcbZH4FP/kUIUQKMahCAIsMgZ7H
KNs3RrRCgDs/uaJh1QyQnlG1kZ5mgil4xmGAAIIxLF0ujiH0JirFly2P89SjXhJhmXWjbZ40dbdf
l4rPpg6E93iLGx72ZayV3wRnRF6Wonnyo/y1s96Pm/FSlt9PbcvoxDDBY2yBtihk+Bzlb3PtQL0q
+0mKpnDaMqH/2RN1hZNaPsGOzeKwymqMsvZdJY1C/PWoxT6gqYp4f7DvFkKvqr/njAsVGxk1HxXq
Lff2R9glNjPgwmWe10iiMdM4xNnzvdWu0qKPWa+raQrZGHOJ/QGYD0FZsoe0KBK4lMXNKm/CC5V4
aDaOpYk7/7Be4mfF1OyNDN2origJ/1QDGzm7iSvzTKtid78msw9jaiKorNb8uR6+vIz8sxOu0y97
QXXIdcFCEWUPlDiHlMcDz3r+rjn/6ZEhPmBXjSBxHQ3Aw7U8iNqseaAY6MqplrePp+atIFaNuO2l
Aw12l8kbFaV0OQ/Jxlgn3d9L6dge/VboLgXs23PiilYCBL4Ga10uSips6jiKj5XsOaHD2bhFMXdR
xOYLC8J+mmEosw+N9KJvrzypTRwBPFowN//4X5OUx6bH12XHsSnXs2+QLLBjkqEumyTIQe8oaXu8
L5hDj2IbUJB2oc5I0p7eAMWbgogPsJAoFcufmFa6FwLyCpVVlAX3/G2V+jgRwHIJ+pGfKVr+4wM0
3LndnNK0CqI9o/Pg6VFgjXGJcDupxkq3M4ZX93lUe3UQklFLjCqMbYL361DEVAHzj11dOR/I3S5N
xOiiCr6+kzUDQbAnrE2riPZDpAukWAV1f4fSayFHd5WBSoPYgE5Jr38g/GzkS2YRVg8c2iUXDj52
3xoTEVpsJxPiiouCMFTcMUA8seF6mGiIjU+AlZdBpsUB4nJyeg5k8vZv/XSCkgKlCzkhpndy9T0D
mG6aWz0qBQ44ckAFujy/GL+nvXdlARgWRAg7cJPCetwc130t6I96DvJlxyArLNuLy9N8UiEUDo2K
Z8spY+A1mvlzcv1brelKEyx6UoQ9eaBpOpOMrnH4aCXADlVy2Hbhq6qhENH84dBqRB9UNs9iRUaO
3EqmUDKVbnmkXwI4RZog5wQjRxcEMUhXQMB/Fr7Z2nZiL0tIsP0gwX5PBxjCzQNh5WVn+J9t3cJ9
K+j2n9f27BLHLNu2FL5As/f88hjBL8i6Rd8+IKJjlu4qN/+HefozNsR7ViRRkYIJRLghvdQlitrj
V3sA+wgaB2nf+fzNMf2642fsNlJ1GMkAuEVPeUI5u2clv/MmjzmcoaEZk2m98a/QJp9UR5YuiKGT
+M1IntyKfxOcKwtEdLmfh5NIJcxWOmk7tOoh3yo4jQNPRUDOR3gA8m5uwrYGvL41REkspfNJfL38
0Alewb3dVtpYNYcN5F2KZer32lVfGhPgj9M6HaQTGViUahbQ7MyzSMrgRNUUw45RrH4GCPOvAlzG
zqR/PQa0upwouuaIcU9GlZ2TJ57vfYN5GaFPHs2IJq0dP+xRlLIiM+LUdbFNDS5PNT/hc1BmhzhT
+FJFXAOMnwuLFgZr3RQKyZwAwYEOBfVxCWrTGIzo53om26Uygw6x/BqtMKvrQzWOTxr3SlR6Jefd
zOQa75K7KAbIwp4ozhzPXLQQOZgt04XnO/5DvICFWovZRL3FV71zsuuZtPMgWjKqvDHUUDD9JN22
cGqI4junpjTxd5Q/zzq6nHpXySoIC3J4+e2+pF0o4Hsh4gmUAbIEbkjUMErfh5LP4x35poq4jrzu
YsMAnfM5WTx+FS8CqiWW8fU9lOwxTxV650Y3EUmWsCpYKMlqKgH+VxKLpDAQZBXTO7gpA2hP/EpI
K8cDsK7eHvCR8P67MKCMS66oTfGw9vQ1U5hmEVdiiOVwl8c3TlgVc1VfFqVujJjfbZOkRCAzf1xr
ZSdUAUNjPO3n1Dzq/DZKbz8rJXMGB5M83r77vBadSi0CMvUsUg0621jpB7wsktlUYiivkY0v0UQp
zIOehiqo9lUsisvsnqH8VUW83KMdPEziPaN2DInn1+iybaG5TNR1cb06Hv7/P/5u65tVScVr6Nhp
B7WEbcPCdw+fk8tyHZvXS6EI3BtiFOO7jPQv1Jqfu91xL2RBohkvm8/YZEFV+w6O6Wpp8x/M38vc
LCYSFf618ClX8tiEucP0kH9gGB2eNWcp1ANE0fTsbs2ZgTVdEA8yXYyuhHhQ7sXZJTkzr0fg9VP4
9zHPJygdpGQqi1eBNaELAo7pm+kTwE/TiZwniz9MomAgq7uHwp5e2vrqUgBUeGdn4JJYctz6yeKe
Rkckd5oNW/ZCby8FhiCgQbofFgmWQ77iXAG+BFMkje6UPAXEMrLGSIUYVl568oNlsv5itL4alSpy
TzZsoMR8UWTwZZgoPeVjlyySRNI9ueaMymSG1hmBXkZdVJeHPWN/iDOvGyef6fZRb1kfpSwzgNZh
1BYFBt3c36U8ZZ9+vM0x8f5nz5BO9DLZXq9YXypIvpopuhMxrvOGAat/H2UojhSq45YNykeB2SK4
xHCOb2XhQqfUFfEK4WPX63L6jtPVvpz5kM4bYWc148YT2g09iFvWdg46do/Fwn5loKlib7KWRjnR
8FHpvv6UHJZMX0BnpmZIf5gYKFs+sxV7jzqzG5YduDclreJa3tYfhU3sgFR1Q7NOUKJCRmWFFv10
pjBAZ+yajOyls/WOb13UeyiqhrUFxzpaHt2to7Uje/ZArB0oZVuN2EIAcl/fiuoHyj+QDta9T9DS
KvgSXqDJC41tm8b1vG4R8vEd6+y8ZU49VhL7Fzsy89SuYcMcQAh7n9ET2gE2Bed8G06dbUaQslyD
hzYQ3u1dhMOE3Q+ECXc3uWnXqkk/DGPjUBeF3aevdA8N1Xhhk7FAeyyW5JhYJmrhRm2Lf1x12OFg
eYW/ljVbZ6jZgb5kb463ciRsG9Ss2P/ovsH1jo2qTMDLJ93tzk2Dni5eDf5UR9QKTr0Bby2zfVSN
8KH/ur4HKrfmK2hIQSN/M7iaL13F9l/2sW0q2KQl6ZdUtTBITe8O1a0qFYL9aMsuOt9QZK0H5ts6
x/1xeIIHiPf9CtJY0x9stlZ0/nMZfpnMHyzG5YwChvtO7XiBA+IUDAK30jLVGE1FFWptpfXv9CSM
5sHQ/N0lsTvpwFmFFYjacrQ3sKUJ1lyywoL94Gg9sHHJQCPo7UeQX8DK3J5SbCRhQWVYZyOt5mfC
uK4GNPuU2TGEV+LhU8kDyqOOCzOAM83LGpJmw9xGmYIB3ZMAWxzH92HgdEmTcuYUW2oQyZXCRPsg
jjKZkXU5Yv7eXnIY4jIjzUweuMVdFFp9fw+6GMl0UNAcVQeJNkUlzVrzbxDbqH6qftzMOT9DV6gw
cHRSLk4tv0/ImzYTnWJu/xiTN3l8syFLFUzcP9R5Ip0bk9s57iwnxAfkDED8/BzjRUSyPFuL1290
rD9FTrN7KuG3jEdtaCGuq8gaY1uzjEar7p9cXrqdsKZ5fmZUGgFcOuRbHN/SrQ0pkzNZjMBU9emZ
9NS9nQ7/+vIUgfZmUzODp7ygwxKPO7sYELa80m/sLK8DN28mInsN1mKvVXTuWzlGDlspPtflH43O
Marbl5Z11l8bAN4ort0lu8l6XHOE6zfqXZ/Ss32IjQs3dLIOlJ/j6lSEfck4Hjosxx481+zwTY+D
/Vk3HK0gpuHtzO3F+t4EHJ98S9cg2RpjiMHCBn5SMZtyTkdvjSlwP20EUaNPtHnZqlfkAqBxovbQ
+KM2o7VQJblV/G12fklrCHAC6SQ45an9irYbcsHPmGyqjytlQ4YW3XxF8r3681uoluQQMOf55YjA
6JsN13zp1fywPVZ2J4yFAdVY3MnNJQ71o+W2nDwOk4aJFDvPZWtdvGmUKJ1iWeqOujnjrKxWKsB9
SIBs27az0Ese4WifGQjiJuAlS1ezewyHleXZHPKwnTQ/pynnv7znnYtg+yAIf8wZQUNfPSwXm9LU
Ifg5K0yu1DJ+W8pJiSVDVBDyx2PVmndAJ6p55Nqjyh9hW6eHiBV0+TTQzAKO5N73cmp5VAtISXPm
ay6+q1XRy4IhUQW+gSDM21fm69vtl0jin4i09Saga0kMCCReIcER94oOmT6WbmrPvrBMrmLRjFWL
tw445dUPBOwUyRMF0C52L0h5oglld/UYykXs2q9FJYRb71IPSNFNRbug9EiMJh8ruVf8XDMYGlpf
aSlYSDCGH+ZveQVfC0dtWyOJDNciCRTP8fq5F2MG1EhQgoqz+WZx11DlaEu6EK4rHzjpxfaZ3BH+
mpaWE6DW8bvooOq8X+tTxYpaewA8iges7Zmevq5USjEEDAkm9HlsqJEqg/VoTCqWsAUsP24mf6Gp
xW1VKrj1uqeQpvay9ILb7sAKFsE/AGsbu0a1yyBX9jd5BD58zPF7kOZBfjtcdSuDNvU4WYeoeh0m
+BialOyObZ0PmF/zZ5zGJ+uc5sBIs2Cn0SBlv0zeabyDVEWPgku703r5C1XezoxhEzjdcVz6SddD
4xS0x4llo9Un4mpXLPnDCP74B+otmxq3B7qeRGY70Bx3KqXxa/7Yq4uTGFuIVbKp5YjlCiTiIgQA
lFqF4NfJU6Q+H/hLEmKxZWxi/wkqTSGIIbxXJZEHtuT9bIZUgt7iamIUaryL3XG7VG2JNfIY/Huu
xvIwv25PgXgLImwMjxenf9IqcqCa4Ygny7Anj9Kw+MtyiLBwjXDOEdLIqS1+dnp9TIGQ0EiqnO/7
i3kB+hmZzG8tZz67maW9xkNLwgyRodjqDVSoZU+POsJ6hqcGeaSz9D+yyeYv9FFYpYeyL/goQZYU
IEipWmp3EqMYVBl1I3UgXekGaV6hRtnke1tATCAU/V/pLeDVWTZ814HI4cLOkmSz1nfS9LyqhcbL
PbCIvBhvAsGw7VzguQHM/LakuOsLpXDkxd/oq+FdACrd4vfZ3xZS9gA2shHEbSD1RfjKZlxSeb0e
QIZQv1WRJ9MJgAtklIQ7KguBmIiT0gIGNhHK3YYvaGtJlUNrRe0FMkRJAxY51hDjc3KTRtBmwmHF
JgyQTjhmkXT07W929khLYa1i7jzAEa+cjcG4aAnVXs3W2aJVNjgU+Ty21meLDzQjKEqmVsfTmzrD
9hgEwCR+R5r0rTWgLqgFvWd5fHIvyaAYMZqxYrybzDmk5v/+Ud2hAfySW2vjgY0o9hNtGvppeunI
1SQ336A1n4xFPxI6RNC4F5VFOG8dXFMPQ82F9H9XbwBNlX/inugbx2Nd3SmHf2/eI9p8nxUQJcnw
yy0GMI3xTgOqqxPvaaALE1UvsiPdJx5ODC4AmmTdI38qS6IEaL1elF1+fCoq/aeGuRlUY/buQxnY
LjnnLUuIR8Td5IsJRLeOsvXU6o2GmUfNciEICxqTFCPoox/vILMYHhs2kcCPWJlQK0I5UwJZ3KgS
+qHus+3cfcY9ZxWUUUerXZBQxGXdcc0JDI/eP40UD9XNjkLqUg7tu0NWabrqFGIUMV8ao2bqQRl3
cx96YRF/QKI45dBBUVbewYLbiOiLijrBC3SjczxB2HwpD+ErDmmROaiRXNyoTqWNM9LHVI7fmRPO
5GiienwBahl2XPC5QtNYWWoEdIyMWNBvkxEzo2wjlxdwxMQVjNy4v3HxguQQ4ejR1WUsdIape0XZ
PMkhvm/BVsDOVeiqZCmj0x8rnT4LennuAvkTsjjqoYQwK7AEhLua6WNa5Z/Wve2X8saPY0OgAyCU
7T+khPKvXEO2yIBsuNWJgoehjVhbbVzlRkB0zBfXFBWZvc1sxozKltTJHlbi899IOW3resOrPnuk
kstcY+j9wHuh28iN5kxd+3GUpP6iRj7mh0ELN2PaNo9QBKqYrRgSMwJ+JTr3TonuiY1Ep+/bHucx
v7hmashx5/sn4tAvwt61IfuyFBK/MVuQ/V4bLVI8HIyR+slPI3UoF0WkzK7Rl5JiA3b/Sk/raBbT
RSXD9P8szRQQ2TZl29u1QH308H7skQyQ+xLlnuVHZo06DccgHHoSkKkAPc5flQDa4eBC1iBIJlWP
3UU1t14FaEXMzetZ6nB7tse2yJNNboQ6YNf3vSQIKlJgVhG+x30KXMiyImWAaM2HyRWHWjTCA4B7
9/mksRNegXZGbOYdFS5U0oB90AL6fUb4NvOVmlpBfq3q4Le3a1ZPYProjj30OAJeFSUJ7sKBEnrS
hcDdD6tyamTS2RIOv9uUjm64rra4FI44kyj4zJAQ3oLk27ORT8nJEkQAeX05kGl+5yLRItZ8WKq8
yiDNu6lsvr0w8OZVgzzDuCxcGj7UDEJz1jTOHUPjja08V+EAZP/9BoQCQR3aI6uqMEXr9MU0C+ky
3AzwFRG4woX01uN8nXboTx7XACgPYWLeekZVEWFm2WTJlzoO+9FU6Aw1vq9AtGh6BZbQoMfQrMML
5gJbWE6HvdB60rcmwVie2xrVMBH80OnWHTiGmAgPKunAr/b58sIkXgxw4hCbDOqE9Ba6KZ06wL2R
48XfOgbAhk63EXfMS6fKLPSLSHSDIAWRNtg0huKAglaIqeTO3ACcwfzqEX4JqPUkoZbJYG1lM7us
2RVgZsAm9XUnIKbPqHMNlomj/FCGZLyo6sLrheFCiiWuHHh1ZveZJDX2FTUpkkebbFaaGEcTeNKN
tjM1s8llciCppcqaDO/uGdGefvRk8hreKRakJeX75eiOOwFXhPjh0nh/HFxWvPvTfGRErObh4mzf
k2fHDwCxihcss/v1zFh5KvCuwV9b19+jJzuZEf7PVpnO6uT2OBuQ6ypUkTM6YYiYaVggfBrJrdrA
t6SbiHZldyOKE1pqgpY+v6UxynzMeYLNaPaSKOse4gw8HXsItNwz0EN7lfcBOuQDYGbr7lvQ802N
z5PXw5KjUtiZQUE0mNHUe1IwDg14NSWxqXISx5tuI+5MbddR1bDmSV+eaN6Kj9W5dHplBDAFCgU7
0+eV2aAeMNSFyvfXqt+7ycamXyXTXpqBagxOdidJh3d8+p6ScEIHdAXPOO59o6RIYJx7itETq9g8
/R7rbAK9ZeE3gcBuzrbfcenhuDsM97jelNHMqr/gzwQypWOhHthXoaabW3g83k2qhD1/gQlysAky
j20oMN3wC9RQbHIhl1B/fxv9caL7IU3c6gRRa28Wi278Ux7dR/+xjj8JRjQXpivMopkPmCbmp1B4
6uF5VYH5eEFIxNcrPa1W1XG5uuVWzZEj5lib2fxo9RO+05hmpigWJ2iuT1fksZV98hCNno5yWi4q
Njx2RnSImdM15wtK02Iw1qNMo3h57dmtmd1tGZ1Ld8BZoIF0S9qmyrCYJlSTzBfKjhH7Yl02EGCL
NsUtfp743pr/AYx3IKM4Wa/BeooI6VCPkWES9VffpHJooGkqgGN2I+EU3Ae+ZSSBj4B31rzERbo7
AUHxrl+lY64nTOEfplL9Oj4iNiCsXJUIzco4+Tl8ObKuhvyOy87kHej7m011uUuMSFdQtq/OSuA/
fism/f8ejPPBkQAsL1d6yNd+g1WFw56+Uoz4C+n0Fv6osmOWBl8XEtXz/O2VRP4Yp7TDunhb9Hlo
c/qoCTxL3dlISg5MXWuvxfrocjbHeQlz2Rr3eV64BxbNdJxb2IJVYXJuytu7t2+y7K67zM0Y1Yo1
wUEoT6lFHvmv9upqwon4+S8S3f8LoVHUnncl+wRxiUUuMCeYI+9uht6oI5w84qmF+PkyB1tqTPs/
idkFAptmo5V+hVYHjKrmesNYHmWaTZW5Rmcat3lzz9e/Ps2PiFSpU6jWgsVqFpwprz3jq9Dc6Mah
y4TWAzK/qe9xdOcLjC5NCPKHjxKyUNsV4St+FsScP2Kxoo0HZFCpdxTEN20f/zpQ7k/3IKLSvlcO
IZUu+kWioIbsqj4T4vYL70UCClfr6fxrFGbEOB0L1opzeHzij0c5x1L03VTGomswif4IMGCackZd
Kt1T9K9a0E7B3qG1djOjWFa6D1kyr4U1qNrzKu6jqUcR1GwgNQJtEtwgaXRZVv7VMnNj5/u0ne3A
ABNbpHJm8FxvxznGaihte7wgpdDz8yIWCpGoRjRKQocxDeUPuAhejTEDtOj0aK/SfgIuFjKu87pH
eh8NlE9Cm1Xkk2e2F4JIyG5zQhuORaPmF6G01MGXHAJ6H5/YKXjN/tVEHMUu7uJjoEGcfOmKyr+k
POEOj2LHjaEl/i8VK6Tn+nYEYLZjlFTITMlKSKkuSYODRgEho1x2Frh0PHkyw5xN8PumFiqI9vn4
ndg+C4TxQLAS7Twwv4eDOOqFykxCEKU70KMuHFavgp88wnNQuigA+/G2pLYxHbbqRu1emdFQCa2X
FUwJf3yc3Lig9xOb21/+lK0fzqYEg4gnqDNvNuir1YWM4iDIBEfld8oMwMAL+tE1UR58c9l3xvYN
PQQ1bppyXh6aaqXqSgzdFqWk7NHiXhqA8LIHnQFpKUKWBxVawWA6hl6a2BykZft6jPxT34/ZdVHZ
sNgrLfon1qOUEsyJ47NkTzmtWSDKmJM0qa6SXMplTvt7NdjNWKbPW9Gs75RYJFV/tSsZ+fblU53H
emQfro8+sCTYAFKoH10nPkuxyKwWzgTxTgDeCqZNNlTTJ6uOSU8rthT4gbiVXztzyIWZHzR74gtw
QGqFCTm5wtluuLUBBPTTwekX/0d6gRbH2vsat133tcRVwF52w52/7bHTmMMvfiQnxCnKnOKOchkV
3krqQM7n/ygnrrzzsRu8g99oSemZLNJryio8IBKSYKvZGtIFWBzUgCm7dzErdxeNgfgCEivJGz1G
5x1GhU/S1qfyIWOW5J+XscFJ1RXLbJnrQn30HULi9uRXGJYmPrC9iVhvJdcyMnzvuzJofNp6ZiGu
XJiKPrWWxv5gJVQjXSESDvKj6YzI4nuQowLzKMtnIzmvDosHKMnL/pKnVr6bVhDjOYlgPmy0SH2c
K+5loffcstKLKIHBrsBR/JMUosFQmZbkXLPV1OvnDWeupNdO/z37/96MKz2ghB2zZ6gnkREHKQy4
KrzV0A9EEr+i8Kv/nQcuNlWM3G8XZ8prHY6LbXSyWn90CTe/nlUs32g2jc4j3xZAAJ+F0wdTcica
VrBPqFYWVVuiYgfcW1WQeC8xjCLPgTVJTw7ZW6+rmqABcpvKfwhRqz9AL4+XnU+Y6bWasOYRTZao
WzgGXZakaOkS4EeWW4J7s5IJ3ynYRqdDc5Or5IYNztgGlIGzTDmn7gbKX1+ODq8kiMhtaOPtkcxY
ktkHSiMr/+Bo7DHTNdS7qH3D7/QcAxUt+NOtuIgGc/YrndFt1SPPFOqCF+NjIWn/dcGItR7wqxx5
Y2DgJD5idGuxTjuCXMDY7nJXjQAuaAhQvkZ/ng+DdGOKqF6wdz+i6rc0y8mD78+OA0GcVBn3LNMu
SmkL7tBUxjo94jUE6GtykgCi/IPikIeoRb9sFZwGqdJzbmfyNNZ5FqPsDBjkNnqEgc9s4/VGUmY2
y+7GQyGZwyO0pSQ2z7HwXDjFKQOLG6L/9YakCFCd8R/ukcCOb6dAh1ovBIcQksi2+2gVxcWC0JFM
8RXykwKh40CSxuIciQUgMi+P3MzfGSQjuLkVFDMjEWaexe3V6GC9u3ukubKTl9LwNM6uIvR4nfm4
Brg+252255VlMSeVIFCH6W5+uY4ATlgnwHt8tmuxrajIYZovU3TUSMNB5Xdhqh2Y0253VkJOLUx8
v5VwnYyhyjThCrrAhj6NQSdATkrCKeiryGhnpCIgY9TPxlXHJIKZZEDirfZ35b2I0fGqy0+clyBk
FxMw8FZBbCqCaLpG12hrDBPjMvLUZ5BMeixkpHOyH4zHr/Mrw+kNOlWCY/gZtDBu9keKxlvXGDxk
wZ5cPB0iDS6xwzUa5EkTQ4cnkZZCISAy2pYWJeq+ZcOsu7G2VSI2bmT0MiilVE0hbVVPZwbVkBvT
RlubKvxp12vvN7I3OP/nhoqj/OQy/BqOtp0mMDwZLnU2WDFDuERRVAQ7L3x/1Ss63ZdgJbzKixno
st86kwwPLEvkCYmvd3AjJpKl6i/lp8gggGPR5q3tKDNVcLzu8ETZdOFxbH7PbpkGz1y08Q9GVOdZ
F2w8QhzWaad//RmirK/cwlnStkB6E8IsKcsxP/CZZf3BdlPJZvreS808emq5vFZEq7ruPpne1Esd
sE2iZpffS6SHOslaepI6EqPn50/4cX8zCPVlC+jTT84ZW72w3EcN0FumZln2MHOrEACo5tqdASFx
eCxLBgrsMplEsG9KqBdyM1kKKlQY11eF9bIl9sRGbuWsrajqKYNiApNKsCp97z51+bxJVPOBCuqi
1CapzLmiMbbr3U2Hsw8GEilqlREUulkIhdYQTFyVpCZ+dAexzksLlEGB1N4bpWiKgLIqUBgnrph9
zxbVmDeDFFYcQBkHVyeCYfIldgSzdEN6ThQxJq/jM+2TSFMVxFryPxUrgZFHMLH4FjPfmYD0I6Ce
sw7/bpck4CmAHlM+0rnd5fogVlpMmuHxNGPcX8OQ1Stkra7O+gQ5439DbJ8UiOYSyctxEP7PIJZ/
RA8va3CdG8w4rFk3LRTAfl4j26DHvr2gglntBHG5joDTSPOSx7JmNq7Uo2VTQg7IvqkyEBogX6hj
y5f/RXO5gN+RUbLEEwbPP/CWhCT5SdgZa+gN53i85pvlruGIn8xysjMQm3p5D2AE+wmnsbZBEvw3
R+TM5plOY6IkiwkUoDSoYyrFEOQgX1mhTCHyOwYNQY580NpCtaW2NyZkp/uN6BPX2P+vunYIrBPz
tMzkmnYFCJvyLqdI09KNK5k02wGktj4dtdjOr/Capfpg1LiHjzTCeISZqjd0SrT92KOULqUMS5Fi
s1gfEmI3RD+LEsdcjvsIOj6+8FW8m/naACHy0jd9MEk6yrbunGvKfdDmwUQ3QHMs+cwGtkbmkGE4
MujYMje/ScJsqAmhITXE479tHVKUVSEobMs28sUGqDZ+5YOVLXgY4D0HGBXLPRuFmhyVNEA8VcnM
0CBAGsZ8Ben4W5mP4h64RZIITFugLy7D6apK4KjbsaC35DJw94ac3ZL/3ylsiymGKjYueHm+3yeK
ptpPkxHzUseKrAnELZMwyqTGenJTrRLUCW9RVAyUMJv57mWAS4uJBEWjzadfvLI25omOWpdIovJ9
JlfWVGME2m5l6gvf1cylRyGzNAcp92geWY8sKjyd6Kah3myCqvqELYJYm7FCtxAdOT9J/+3MSCic
4T9ke/5hlYVeuvSVSkjof4+ZchGTj6rZZ4kNGhbgeNQWNW95dIRBYwM+eqK+D4Fz0EuxMSfd4n9W
86LT4MHk20rlf90v0xDFXDVUdTbkY9xPAaTcb6uVZsAvqdpeqeaIYTGMtrL/iJ1ZA/aEBZC1Hzl0
lZVxucVgmjJKe6mGsoB6+jG0bjmEZiHEdcGCqouSFc9w45cms5cK7wPtkb9rplxGpL91NRTxeBPl
7g9Ud3Le1vy/RxpGxy8XSWgHNx50D0/TUu+sZjiyxvWXnllDhtfvAQkcdQbS1hGGoy17Yj0enpw3
zBwEDLUpDLHLXPeP9pZBfNOlGf3chJHudQbRVHi7J9TSjcDozCQLWUf7/rfNTRy1Eyi31JPiL0WP
QZeUzEE6wyau7KHnS/V/ClVG7qFjb/oeJZZ9stVOVdn1fEevU1Y3JpKl515T9f8C+nwq0FFu6AtU
QY99TIEC0zSpNE20smC10fd/sDEH0lcL43V0Jw0Ok8oTfIXFdRuQk3Jp/UzQAnJC+8DCklYLaLy3
sZ6IhYds118BDEMSbsxSRpEgEMKcbzMyHY57auMfxPxthC+DOMUieW0zrSc1cXX2LAoGceFPrJiP
F60Ya0irMz+gR4/Lw17V8UAMsw3QKBMsED68zVadZB/ZFcu4Aopj9Q79JaE8oKaHl5MttYDsAwZi
mHQRT2pFgxqDtW6gMMGIMX17Fybb8h9NKM5vNWsvUgQDT2Xi48CFqhxBGOo028CzkOEjsMAFW1WM
EiHanOECYnsl2jnvc/5QMu0DRIt6e31ks4eXTTSnlk8ZrXkiFbjZ6ZhiZy+7H1ndPx825G5rxCYZ
GlvJRJUkVFyyD5jcgJPSAwHqA16xJnS26aNoYOV39slTAY3/h2PIx4C1Zd4Snjw0QzDisUVcEKA/
uLJ5Tf7W+s1S5w1CBwf6EbbeM3trDm+/WRU/cDuws2rujMWNa20/C4cTRqT5IzbKhxDY5+ID8HFZ
9sdBOjSiIgqTstB6SEK+vRlfmTM+AizfHs/oER8nInJ1dq3R3s+slH3wvbmqP+gNfedfTKymRXhF
T1W5lNS9+Y5MO6fGorzeRS7SeUT2962bwCm/dG0TqlD0ShMpVS1S701IHsmKZEYOyxhVvRe6EpsU
CU2ZXya5t9/kHOnwee5Vj/sXKZcPGgIvB8mYK1+9H1Et3Hqh8/u9/lrhYgFJZ1Z3CffNbo6/XmDM
k3VHiT67s1lzDntMCHN47tq1eVFsNA1PQIImehosoEiILPf3dJua/sOzIHQsJZPN/Qb/v+L1TVpt
8Bp4AmIU5LIKgiNTCvr6572wuJ7kOuYNgn3XJ5MLvoLk0k7J7gD+inXiLF5Ts8/QC6uH26i+KeqN
Robz7angs+w4dXRJK9072GiusIBHM7AnhDe3JmOvrK0mQZmXuV430U/mbAYhuxX+S3zwFXe5TpKl
TiuPEewAyCgqVcgFCrf0CuUHhtub4hRXFHKXXBCZpq+/rHwr5gk3RHq3clRAFMRKpcqxuGLQLrsH
BJvu2KcUffhKejnGemmkCGLqN0Dcvgk7JO2LFLgVH9nV4WPZU3to6oalOPfqLYiTJ8SbzeDDWsFw
tYLEIB5S9YHAftmmU00brcGDzR6Hcju03TCliMFDF4imOiSSnozay6WNT6yZL93TA/qaKRupL1ny
ej/7SLnoaL4BuPEp1xNuvECv+PTIg7YAmwSJ2jYIuqYMdkHAvuf5GZcdhRZ9cvBx+GazzJpyMk7Y
djveVF9cYJ23/Ym++F5C6SJlQevBCgigeEcNTtqHrd9E4ehxXM1HaD5xlbLY1AixWRPMK3eF4pcs
ighCoBmXyNdiZUYHN4xxFTSt+93NAquOBvluv4F5TiecIaFMjw9WROC8UwGuepOUooWQNmwb93TN
L0OR4ZaJ3eMd+HXqggkdsUDEy3PlEsaMHC3FClqeRx13F8Olc8UjUYjoeImcpgOFJ5/6K7WiOVvl
MWRZDqb6tc25IKNOyZhdLioVIH66jUg133hpbHnNRsz/jgun9VwxDiNapf8FLDQfWHhQ9VBjm4OJ
ECMzwDylqKAerclXTqfR9Q0UQhg/YMEYNwB/PRaK8mNaPI5QSa0iPgGT5tepFD/75sdd9oYFiQbG
gT3IAtSTjw/hB3F5+D4RCKqEyt286iOucEGw9RWnXNphp9/57l3Api9nsBjOQX0KQTejBaDS1bgg
Tx7wnXacnX7KPc7NxM2aThajRdqyT4Fc3tgczIZiS68HVuZn6rcATnKApYLKeFGL1NCkE7HUJpeH
8VVLzt3Re2Pmq4fWD3JxCoKDXCQS5pkvpZ3NqmTQLF0Pn71yYFaOcweL0GcF2SuZfj3Sw2vBl6Fd
mjPWmcS4spAlS04TxXv/0ZUMJRlDmpZBKM23nfROaf1CN0F4lXfN56kHGy/u49uPjgWiELkGg1uw
xY+Yu1VE5R2InfrStZJt7o545PA52GnfvTU7vpMyyfvnHUUfQfA0w0qKP/411aQwK46vInQFPb4q
DysvqJJjwulrAPMj02Hm5X2BgnuUo9ROPA9EEZZpHPS7+IRXfzbJQrLfJI3zpZN9adTxSEFyZLPU
Nnal3Kn/x05BnOoPT3di4HhvXPp3XAczJB6EeSYyoxk9Y8KDXG3BI8E3zZCkstl10dNh+vL0RpSk
0hTc94VGDNb3KT7e4FsoWpTMukelVpQqLy7DVXIHLz0XJB8E9fK7E+tpCpo7OvYcpBpklVSg/CJS
ODsIw9IDQFcmmDptO07gWI4dE0iaK/DqUp3DAICFm2uHsoIXsfPRNj0JpuuUmVYDiTjNSnAP+wM/
r7D8lmZaEMpe07YHmoBKBjXyE0WU7NztEyW8bYnNtO+gfY3U4YE/+5CjgDka53qtXDSjqFu/x8V2
lug/4sd00dzsvXJENJhq/3FWmr3XnC0o9vgyU+lN0PcTQm5n0DaoLYsw4qgFIviP1U7j0dfrBFln
suYnHdygegk7MIaKNhlObuOPZGJa8suzGaDoVKmbKf3FIj/g4rIIToTJjtzGshg0t/rO821oNjKS
TsQY/qxIERpwKfSJSHxNHAkL3pXuks29X4DE6FRnfBsLHH2/jqDZ2FsDJKs8PPsly/GxuwaIlhlL
2vFJpTWJy2wmQ6V/EXaPHrvryPE8hPXXD+DwZZE/e0aNpj8PojHIGLbr4TqX9mijlL3dENGjO04x
wgRyYvt0bOKhFhIYP7VhVQ/TzWa0i9FSOiSAZ/V20ysq7pbuTTkxldqONh1V1C0OQ8HfMnsscbE0
4PGmqJ1RV/JiJR94D5sopoDIji073NDmrzuO9lrw6DEsHdhoVVAtWuXWQJPSl9Xrk00a3fAiacRL
0cLKTeOhdMFMoYgi8P2h/PD266AfkCyXty5OTiMQnUvelJ/O7Sr8ntf94G4SiCwZmWAKR4iJEZFK
fjVpB51yav9mJ2sr+LCgb0eRY/cE74leMext6d/79cWI4UcZ5uUEEaI2DSP4JEpHM4FZ4zB99v/u
WgT03MzVgjfVi3qyIXvMME6Vva9YDeYOlA4VeYPFXFRL14bHFDz0rsOBLIN/L0BkxQe+OQCp/CS3
dKmB0vFSGUW3+i8i1KtB/bFXSpbRFzt4834b37uLcCKQHupI82MNngIE9zUkqV6ROWm029RDfODa
jlo2PbuLRvdI+uVAc4UWo+NmxJj5NhzxJtO/txCzuX4eoGkLotTVx/7PAAefTWJe2cq5JFWNYjpz
3juljHMe/29L0sXkxUIsu5w+McAXRg+lW+nG3eKnI5HBB5UFzvA1qoAu4a0ZcQHLZdb0OtF6ym9u
3yChh6yFs14BI42Ggl026QXz8RAfDASXVczjGJGtGK3dbTHqDjJav0Ip14OUxB2XNrLMJmgk65KA
LCQSjmIG96mq2IWpMBXJFosbppmMBj/yXHvBCL55rxMKb/BU7v9S7U89Ue/LIJlex30LcqA8pxCH
LXk0Ah8lBnAtlDvuWjraCJMvpQvk3pkmN7ehXE+5hyMxgEUMucWbj8Pej/gv7K5NUk2ZmQuBotLP
ANut2hVZWi/4DNrq/Ay8fdWAp6cn1B78+0VBV6aXYV9K87WTEEbHzfelh7tz1Uwmw8hw3Golyrqa
VAZt2TqYOUqMtVp8uXWllzX8Ip1cVKyuALwia3M6GVCJlqfC1uDpacrvMlImIDWrgOFYrrClFPbq
9dT13dghMpfm643hiEipnoSPflI55EHpBB3SKKcW7wiv40MTR42lPcYNMLx+cYGYJICJBUvGcTFU
P7J03D3Cq0VmqouRxzWryUYM6Y+O3CGSttAPsMNZviU8lICtnKJl+MDrFinTceSZh0Q1IBCWHA0F
uwFfTnezJ2BaW6GxNy/7Wg/T7yi+20fnZf6dwEHXSkwAQwgCum1Mx2mrsGeVM7xRCFvJz+RtT1Gd
ic/Tf3J52y5S0KYqSjuLRelWZ1ywNP6Joh/ITawFv1+4Xp0cXm8ESUMdk0/GigjZLlSDzKlYuQia
vV4WqyXMUeJtW4zb56OSul/8z3EDmIK1n+lNQ3oNPRgeVKYrhMLaU+sh9yUA8Lq9wvnRS2/JPYxt
ByWy+IY3sEqb6LHgUBPSQNCVI2jjP55tRUjL6IM5r8Eta6llAA7PaiuejDrsAup2864icICwtTjS
SRaPjYyZ9cB+eMzi1zuJg5RZVM6bNfURlbncX5yhqaDgSunOmcDQn7LDcGTmRugANn0bJk4CZpar
tifFfcwlLqyez7GxzKKgifjk0bUQ+9DIkG/5rFS3wbPEA0F+Eu97IEVwcJo1ghBW9emZ1UgJ+SXE
4r4sYYB3TAh+lVR8N6ddjTuRSrOy7U4HzxmHtWxhQmz7eWjJIPkyEepnZxeOPcKu8tqVgj5ihuwL
45zpzfGKRCoCr+iZdnP6fAbmAjpJr5dsPSQ6A7TkXCjnD7TkAvUfuxgXaSFx8Wo0OBBc/wiOoiBK
cZV2jJpZFMV1NedxSV+AeVgh/m1eaN+z7n2b1ciYv3qq19TmOqdKUq4wV9XK6Q4W4EoRPVNNWNUz
npY0Xmfsa1pUnIiwQFy74drhaj/av9R7OvM4oFDWvFIcLQB2wYn88shkY6+1X6FXNGSD8IhQ1/92
Mf/zftAb5hdYf1Stp02QWxXaWwXAoGcSnvi+8m5wnqfwNNcWdOzH4rEfRrX7CbIwygg1u+6Ydm5m
O77yyJMgnSO0Sqiotk0Gg7ZMjcG5QgBDQtYubqrfixxtuH9KSCf7qFS2onr7O4sBYMtvzeBqiKMR
uFqq4gZlixPmp5UrStV3E7f+dZYfT//Z/UoF+nNUdks2CVDryWfcg6IAaxnd0uNuFvBKKZbxO1Cs
ywYoc4rd20qpWxY1D0GE87n9aOVGY/x9zr1sReuReq3suOi1o+IqOP5/YdlnVuPteXHeHBIfi1QH
CVK5yP2B4W2UldcHCRtJFX4njo2Bo8b29QpMJIDLizYowW4qW8vA0GV5cNjGdI0M9znBMB+wsG4T
B7e5OIznNcBlKzvzDMfwuHf3HBASnqxUvF3iVkZpJHtn47m1X9tUOSSmgRd5GQWFvE+nqtaRSnY3
fWINKhql2cIUF1Hh+5BEPAfwAVg5ieurz3T2jteVQPa7AYNb1Tr1Wo6lFAmOs7ltIulLu3IdNW9d
6zUdWE5MGvflBwISI92/oUzsQAyKv/EqgXhLJbzunVmhzwVVuElLfKGpb1XRYHCRPp8V8ttWqVYA
LPG682XRRo899VqfRksDoaKRqac9g6ozVGdIDRH96j6QDhJjFJCiY8BbkZ992gwDzMnEGhXdgdI5
Kch9SvCoAmz92V13xGfyKq1gVThs2SZZMQKnOlojUdgpoDIclfbsGO1Xfrv4gtqN9NEUXw2VOiCw
/tqkCuXyC/BlaUxZ+qURgnIyPEC/FYunzCI/rZfyYq8aS1XVMFR4x6KSMilkMyWXLUByrjEtC5XG
TF1bNgvgms+xrRM7IHwCHM6InjRa7hZRd0fRHZRZ2vA2H5VEWesFQoO7Mx4B5O5/SphVCLypS7Bf
ywn55BCGjBnhTEJEXUpWTgHuoO3jOJrMPmgoKePreCf3j4wuqQdizR63NbMDKYlUb84OoLuhaTut
uGwJQEdu+JsDhc8kzrxkNDVanZE35I61X1AtVqg/+HZ71hQJnapcXSOXOLZGe0+XEYoSKvPCYKTD
NiaUoB42Kv+j45Jkvb+7h8fGAAPOXlGmpDqIzYm72Omir+uszp4AkVbEOf/1uwbJvIssR+xpiiqv
ySD89dxYvWWXf1Iyqba27Iug2lLNxDgG+Icu25PVJWJhKdNb8TVCKhhobInnrjaqxdJ9HfDg+r30
X8V/hlZ9DX6FfaPvOfELdJU6EI5rKbuKjxn5wVxBl+u9SUteow/GfLTYf34/t49q889/FkrIm++v
Z+Wplkx+BbJzGHJrBrtxCWUDdsb0w0by9oQ4X4JJC/WBZ5Si7x3YYz29u/GR6+7vdikek/auik97
Bv2/mAq86kiOLHhduHeQkvRqonnAC2CvyxirMlOjsQqVi1fnTONZZY9Aix8Qjzi56jt5IV8UOd+S
YZBIJTa78U62mWipYlvbY8czRTnltS1HFSUY1sDt/14KZXY/8feRLa708NcbCUnI/SVRWXjvNbAZ
rodIH74q2XrEQhrt4qVCC/TuFP/3uo3DTJNeWxa0VVGHDC2NivM7nWVqGrelo2LS16ZbT5p0IFr0
c++SVvioQl4XmtQ/ngXusS6aXniTsrvNUphQMK+YU2HeSIc6cPpBWV+d8FgTf9Ut2lu8jaJivjPz
+vixxmCj0aS6G5DP8w2UCF4uEv2zvC3ffNEB99R6CN68q19SJLz2wF3ECtOmkOdCympmi6Fk3mfG
C7EHt7Aju2MpomfUWBlb3G/tsuJ5ghAN078unBjjshFyB2roPfkK3o6pvwG6p6650gi3WQf5vRg/
VXqmEUnPCDcnKTIdBuWjNwHlxPkZmfUI5IMDW4VWzgLkjPENRn6NHqr+LvU6M8EdIYf9Qk1EKKoY
LYJXbARcFmMMOpR8WY2VmxpVbJ2aNK3yYxqjQ8SqI+iv3AO0TVMSHsj+R4fRZCKGepK3oyVF80FK
YA+3moONXwa28HJGGXyyyNZhn1D9+d4/R7EWCcMInrm+PoHoWK3vftzw9P9GZxr3rodIZtoufCwA
L921ww9DaTyPMyiC9mIvqCuca0uixm+AntXev3hX+rAjcf2v+kxRg5G971mrJijX5ZLJo/k6i3yI
z1ISuR27m9wtVndFLEY/U5qmZq9mpZFOBpyrIDksCxxTff7Eew/PHxI63KNpnAqG7UHg+0FCLcrE
XjhEDwcl7tBtjIZs4o114du0BRZ+r3AoFCiI0skDYGnjxtdJWxYDILeSwZna9TaoaDBggadncKCg
nu3/Rc/MZW4eTqh9zt4gEo4JnnAG7wP+mEUp1/PrA7bCOdFLyJ0xLoSHj4YeyHUT5sKWHU5FkuqD
8AzgxQB/G7m5LxX6nSjICH6G8FGBZpYBmAYx4UQtLcA3qYOEcdM/e2EJZkrJbEt39hw3JFLvLDJN
TBT7rkY8ZRvTIPxs+936LN9oK1xycNdFdVUQiL/mWv7TBQoR7Q4zY9lbEbpvKJA2SpbB2RPSIW5z
2MjAlZyf3MnASGdCYRB38WP8y0e2dAEqDciVppZ85ciELgIgkxPpKnjBeVKzjI5yryfZI8Livy6F
RZ8T5N9tNBYk5qU7DEdgueH6QK/yuq9t/gOp/3x3DFW2rIblwDgU09XPYvZRZyC9SGNC6dV680wN
FLJ0mwjQbhNM6vS+MZQDl6XCKD7RctTn4xThn42vJtWS7Na4wnkDGp9+pzHEnAfSKjvNN6HSEN3F
fQTsG0otATL+LA2qDslmAS4E7m2lKG5Fa8OYL2R2OUlF0Uh3Fy8TTKsDjr9ZTCPGjCqHB2DXusqj
tfE36Wv+RK8CcSEgjAEb8mj/wOPk5N5b9+ZSkUO2gKVMKtLrAQxtc/nmPfcQMsqfZRic/3/W8S+p
333hauWgtKZvX4B+KOSIpdT3kUG1TyBvznW34Hl6Af/5EnAbwW5jogae1h0TUnxdPB9cAP5BtZ5s
VmA0MM9WVbZvduYb6gxiq5mZF+0wFzX3YmlmkJhLPB5cgbtBORuxR+oCvASyzzGBnIGUcWI3oyTA
fiNT0iHDBwbBW3BZSjAF7yoJ2fEVERo0fij+ueAZTbcuAFyejNjhAeASlhBFRdRXYTjUUXqO/I+J
n2gUmQzg8PVOwfC8e2NDFqIbl4muNFMuWvYozw3wPVb3us2hV+jdxIwVW5wUoSbR5Irg2CoQeNVY
SJ1WAyeqEH7e06WNPJMPF68Jd/LaA8Dtvj4RJQVPGj6MjXpucSk45hahsSvs/digiyJl7NC53rnW
FoRsfgePX3i1OsJSXvB1BNiIvfrvhoH3EQBXKeTAc38p3MEOHckGP6Ft6CEM/KJX/aLvlzvqY32Q
cNh6+IDwQLywlyVD1oAujAxNECky/KGsrYY9mT0BUL87G2U4dTLRKJaCO5KIAIBH5vyEsIGsEU10
y1FPRVWWfW/Vh2+W9BkkerxohHkGEnSy1O1XxGttYUXnSZjISdz/s3URgnU1i/n1rqNpCeEOsqbv
x/jcCvH3qpqCqgA4Tci59RzG/FfGiLFH0Awy6SDn1/yt7NP6Qi+GEbuKlJe6Mbt6vzQCSA6PGhs1
Rxmber9Elm11P04T4lGi5qz+wtMmKDm5E977M7OMEkaJQhbrt4Id646jCyZvttqDbo072uLjtCX2
VSfdbV/23aG9tGQ7nVB1r2+ShSs6kHeTtoh3MjGRLkwin8Hz7lY42dPcv9huHANwUZLWhCaBP40i
mR+z9cOth08hATau4/AX1T6n0h//Eml64uV88YSGHgTrGUdcYos5NEPHbWZQmH5KHYJDybPVFQ97
56CoEVsdp9MGzdW1moMy56dTKso/NJe0beymUra4kpYVqHo50Uu5iOLwQYK3TI4lxWXNlfHwkoXq
v93XA8YNh0g2G7MyFzhgSy4KydFAiOmIW5+N780O9Vhx/E05U4C+mnJL7fRLtlMctMeAcgFYKRZM
l+wYhvdvmoEJ9p+cZzjA2cLr9h7ZRo+VuCvtHVGmaoQBNzTWNEI8pzjvGScjLpafhVKg5uILPVsT
FdbPVF/vdlH6Ztqw0gKIxXDqMr65s9Vf/fjVoSjPEbZGo6juC6dggsBRk23AzJv6Cd67RCpnFFWk
tjTh7Ryyr5JeDwaJLtEF/ZEmmopGMw6DDCAT37hCPlQ1Gr7daMieLLsJuM7RyIsxPSES1kQ/NTXK
22w+CcX13oSZFAMyeDHKXwvz+lFQUFrOKTDbepMrmFJ3NJVdBQdkp1JJ6E8feLdaXc0SKcvoBR3V
Rd6P+MmdKcgBHgZ9Yw5nYe531IgcU0FiMXmIBzkhKHUKDJpMpMvVRLEWec/XarvIJ96aP1/v7KdB
SsA9Dc33Oedi1HYmjtJvCrqyJbRlZypGUc5GjluzsoG7pNd70TXcMUyvP8Ui4D3szyToBQtRgSnV
34sSNWmJlwBmSULO3u3rx6JGvuEFL1sFDJ1VFHRSJP5UpK5gwSR49YGjHTmR6bjDdPtaXMiGgspq
DJVLUGytLwK7txCcp8cvhhML5FFRfRm0RTt23hHMvHspO7YbewX+GhOrkWS3m9tPWLdMT79S3rlD
xOAunisMME43gCVj1vl3dYprC7+UFA6OyjIvDrpdTdykGAcxT1eYroouBNfmpYCCNXHJaK/XEhwX
+2DXQOXZUzoubnEqFJ01M6Ru7jbB/KozB34YjDY/pmrhPZdtA5qhpR256B4+7Vzzp0IA2xjV3yM2
2MRvxlrAiYaq9jwomVBQdZ0l9LUKO9n/cEvi+z8ebmewRoEbD3N69oAR6++S7OFaMao22rF1gKbA
PIhljwnkgA8oTLIN6HRYgsEF/UIYGSqcvcynePktiiUZBlqS677ED5p4gkPLV2cn5FkDC3TPYuok
o2bzn/HlUmkVvFXcVcbcijAKPoaHVgZmQLni4JqeRgaCxMH57P1N40tnQXWdcmCWbGLg9jLg5Tn+
cRg8mpaG5tslFTslccUgHJro5pHbq06AjgZVWMzD6AUjZCrv/cVNdhy5PT789wbwyv0OJ8zmUwVA
vzj21QQrjVmdUvhsJ3STdy18Ph1Vpw0UhUqwlTvHwvpyXenEzhMJqhDnhVOG3d38KXlr5gfNkXe3
XqJ2vTaudqXtvugtnIdMnVf2Oc0fqIMVbLctSLf4pDYMWHEbj0Uhl9njpSG+w8pb+TxnZy89Edfx
PzQNI+weAuxlaOlB+bMhOJWyLfYnXMc/MJUSxMtp3sfabyayeC3aqQvw8Y3nkm7q7dSlq7s+2H49
87yZ5MMIgm8aXRrDYKPmxLlkxmF7q19i9K+yEOR8tgRNcrQzDzI72FmLjZBGnMpiQ3FfSEWG2fkU
U6+izdC/1FexbXO1h7vJED6Rg1JJLxskqlSHlvmWtoAdFLE/IJOZCvgO52buUZntwbK7xlFhSbD8
dy1vZ1kfHEW/r0WFnaNvHIqEPWsEYBuxWWqkKBujWYUvAba0/0T6iql2sEfBcBu8kB8avGJoyl1n
QxzEKy9yzb3OHBEkvkVrOSVNeYmC+/s3mNbUyLYbVItgEb6fjUE99iWmCYHbm2chqf1ndGRNwdHu
3PlTboEv2p1IEhgQxS2wucY7CuAt8+QlNun5Ue6bdgHAZvY6VsDIDPKunfjeqjaTTP1awdxmdX4Y
rV72w6RJqUtiLOzQP5jNzMZA+/BdGhE2+X8jjVLXIuvINn7g9HcYnYU4ZSV4n+pIrz2VQ/Dgkkw2
03YMjxE49Pn+Kn2BW4eo4rPJx1TJgjN0gsIzHHeKuWRDhFajuE6xCqEJMOYPjmdzENd38xXmKLIl
eo0P+9qgA17G7G1b9EWdF+54HO/zrxFoJAfm6f5ptq6idscA89B95Mmv7Eetj+NCZUv1u2tgWKVA
9/NDhGIqGzi/HdXjrHB6oIQkBX70lma9rOJQgu8VA32UNqudz9p8Y2qY7G8bbsYonKq5oPYfSTHZ
eyg4w/XTWGgD6yT7+aLU11kTWuJFWz/YbsE1nnVVtNCO3zvnOPDyFQU4QbdMVw5NO/7VgDnsjCkQ
w2k9XOUU3WJm60DAWy6mtAP578Pf2Ew6Nn5hiG1n5/V5mLVgimTw2DKVJxcEIIj9vYLHcuD1MHKB
aTd8rMM8dSkP3vzaPIxtJG3KvANoip35FCmEhlFoI7e3R+0K/EabyM0aDuqZYPrMtAMmXtvZBGM8
xQksEGOmsiepog/RTfTnXTyA+7UHvhgYhzs8cqG0uLSUejRsH9V/ZvILIw15bVCPqlRmddeGGUbk
bSitYvXtKNWyFZ+eCYdvJZxXseCZ8iWI0h9vS2KS5DDjzoJcVwsdYDdyTsCLtN9U++d3kHdY1bKr
hF8bKUVgh1RC/xoJKAcMlsg3b+VZ+4MRWsl6z1bs0wwCnh4lmS4KNDKAahsbTxVvL1nDBL/CBRTT
aSYSJPFSafhdkDTsE21xQr+EDPCkoO8KMP9ksIWOZMd0hYL8jeoeoAVu4NJsmKMx1CvdgY7yh6uR
QHjidSNQJDm1FmrmjnqpX6tDEoHrKM7DnngD6EM3BqfHk17MrkZ8gF5lHozCTYPocDT51iKCHoL0
Ll6ocHWB2UgbDCxX4AFIVZSgdmaYHDGzPYOnSwJWViZN4dyONwr1TsG1i0tvdgzgAs7zsqp0M7KU
SFH3ka1XOD50fSYBLgc6RKvhOGSVDXfDEMWWi26lPDReObtY81TIGWtM7LGPTW2HtCt5DNTF92Kb
yCoSGM2hQ228I+94SvkJ0TRdk7zkH3kSZexLwKjUSPr9dO4dYUd30q19Y0N3VGjBECAqXUVaqmon
KsHmbENnAgcx6NOnwpe/0EGSRIK4YXTDYnq0gkAAyJt2cNE5PZHcVRhlIr6vWuc+96CpuQdwH398
ORKdT1T1FUGk7RMWNphocYHBOjXAnKx0gAKRwCeomA8Z/WparbcaiwRfBDfDekRYyIUeMUuXh1fG
bcVhM/EX8ENdyNOhh4bSWYo6OdHizpsdIRzC9bGwC3sbLH0mwdrehwulQSPVqQqCfs89btPD6xTc
1WRk/UXgea6TPsp+C1oq8yvkru6zQ0E52MBrTYYczAr0BJ1eqOt+PtQCMpEpTQKOons1YaSFlqfH
9koZazhYn4FY88Ks4IoDMMt8Rz0/1GCDsuGOpqs1qmgKo3EPtaQigmOzJHmt4JKRfS9XeSCklLOS
VZz88ZsiwSlfLznOj/kkg68P7JrFjd8KrrH3jO/cQPfMVOf6A47gN6xoajjBKdRBn2Csu4gzx9k7
uw1mYhB6pB0sT2cole0nEkYahLehP26KHdlgbviAIfcmosrVccFDynzG9KZBtn1SciFQuzeDqIUT
SMmse3sMoCDHwCCvlLO5KeGoS3VQX312D7RX2ua2YcjSxPfNCzNGS2OxP7DGwRcZ+RgZCDvOGMqT
3aASwLbq7EPySoof7uQRANEm5HQxacwVfEvprhkOB7UuunvJGvJFgddxrplaD6B4Skg0ojkCKbvI
/k3h3JN5Y7Ty/ip5Fo6ZfGox5ODobN1rJVhIK9um19LYDRh0qvJvVXRXZ11VHvp+MCUXTWRX0vl5
2vUoqdpTpNHQ1esv51ZognlhmueMIHaWuMeh1WXZHYsoUMIaJJU2sk4LJgpbCvvnNPVhyLH2qe0Z
hyRCMiyUEdiboIAgz4UTEY0q9aMo8WH914x5eXp0Ha+6RujxKIKTouGEQob3O6chGJ7alt8N4Qqd
jTUR7SufX5GCf27iOCAbgHq4oDiWHQ0MIEAaGsFLBLoC+DbuYc5cUJb6UpLu5puT/4KqzjnZFWlo
mvAANoMfZvYLWV8hM9hiKCa6TVXiMH4J0vk96NHLpCVFjpS+/gYQdfq2QHTFFkqtRIr8NGSq5NQW
GOunAU46nHB//o8RnP9AseuWSPZHKCWPvTOYjYvVejpjiqWKPO189wA5DEIW+MNO6CbUzjKkZcGt
2HwnJR9LhbDKqrtynsML4x8joxth0BNRaJ3czDH0m0iMvO3ntECFUGJXKlSV+HG9HMvcfhkVU70l
irjM36zJSqxU5fV3L/qO4u7h5tQWcpt4wJSwzuPu01AztcE6Z6z/2qNPFHmKC9kbKo2BxCRCbkE6
7/L55a69PijrvzYAKl0b3dEKf25fD/KRzne1d7XKNeVSmM1ywJXsI6Z9wB6ZtU67DKvldvl9ybMC
I+XOylusxjpYwtbu4cdDAYPHPzPMwZtwVOvOJmJ/s1lABLijX0pc02nsTfR9HegCB6HXrGdrHhMM
TfHlH4fkTxr1qrjTyFBWxboKRoUqtjSvXBxacJHtEerxA3CvFX7D6yyDoGyF93fpWGqJwQ0R2Y3P
yv5eOpMlCWdn38UVVH6k2zoLVRt8oQybqyaE6qlUUw6lAdJOTXyP5uBWY+6SK0Imf/AtlrEf71Qw
alT4K8/Xhuj9595aeGhGtITA2CJX3WcooovB1KMXLggLDatfwgAZJT657n2eKR8a0GH4nHWdWEEI
V4iyD7/mp19ujLJKmFf0PH3172wf2+dZ/zqlab33i/aGavLy+tSN2SKo9DYThsTXK+bxGCaxYqOI
zQBmmuNm1wIad+igIbCR01R8tQ0LL6ioRbWMSinqrFrx0eNyKsLOtrQFLLz3tWqPlwxHPBY1ojHx
vGvIG9DiaFyWhqcEYZj5ZTvpds396kqRTubd+ZiccYJdVvw15spBFONWGFy3U+ojJu9mW3t1l3mK
izqRy0PikL/LyD6MrntcnsG1Cp4/wjSM2uNkmVJ7OwNKrBmk7MZQrkBGbIiJRiFrhYVDHn/Qwjir
riGapqh43kJ/XHL9SEW0UpRy6ent/Hiblv724SI6AyhTrEUn19udbB20+zhRVvhL5OQ3PtPOt1Ny
xE6FcB0xGy3gXgE93PKpqRNYcBqOOXD9oqmqPG5GOrw0QNVvuU/UH6BZB4AwJJgi3N5d6/lKxhio
htknWvGvKa0LloYKj8gWbiW+0yW1/DYfuKgDFO0IbkJ9+FRhvQdwwRmuf1++pkYq8zSTubvjh/+C
jtMoaKtGS9BtRW/wewRDis06Qwv9Ky/EwB1AMI1o/A6bGONGwVcxCxAMR3MTyeJDOgtjosSHAZ8t
69mpBqjABx31hDRxPu796fJFrHXfL8YwRVonojmZRIDjXW+DfrztuwfD/IEZGzHyEa0pJ1sovcmc
iWbe3uq3Xi+MHqZYGSMWT2GFagRuQpFwuCQq5tcPVi8K5CmMYZzXHvZOIZWYyddC4y7mB+xvvFTj
NFnT08/07/v/yg2BMPmzwsFbiTC7Du+hr51G4FLr6wzdgoCwD8XpNkDdwK+TGUqGPVNAsSVS1qU5
6imDxppHrWfaQNVpYfoSlYVg6mN/6ooWPbrufhmUUVAvia3zW4XK/n23rQVuTSQnb+1+puS4pPyt
pAuA6VDevyVAyXn+BxtO/DW1nBe1Ok/wT/oScpXn6TO6CW2a4tQuEaKUrdHQT2Ua/JjGASAVPRO6
VLrSWt4rNuiT+urs1VE4Quy2PJzp3ii+QnqJEPTJgRmK3zbzPEqSXMwcQtDynsWK4+z8I9rHG6gy
4iTo7nCbCO9+AysNFxE/nuGpqTjsNKRxb7GMW/saPnAlQf+LniFaIWirK/66hWljtolTnj6z+i2O
J8VIymjmV3lY9sPKB+krqgycSuBGQJ2+42cYiw8WsW1EU0E25MJ4UtWXezaiC1kP+c9Fgykj0b8A
Wk4DPOiUow9hdBSumJFuSqNQBCVCncdocDWDux8b4lZeawe+G+LWSxaw7U9pNhNOaeA2lICgmOIf
SM9sEN6QzSzNIHtFrPbWyICTKog68MHYfLUPtj1dLRppv5AdF5sTkRM4ChlWIcnYHRhqofXsexV8
j2qoqch9EAi+ZS5keGeMlNtmJrVY+ueZTTPFIMeuMmDANYfJ7iVaWj39it6nIKOovfgyOFkMSaUG
7iWgI8iOtWEFq5syrPROJedjLlkn7xuyvFVsokoOtSjDedVj5XL0jpFWoe5+xynW+8gldICV1scC
vAex63ch8xHv1kdblhQlPHv17PSr9Mdu5NunG1ZNesP6p4zE82xzp0ZNMBDUJIKNhOuZCTUH1B8C
EkvVraIqXt7RPJQWCBY2U3UmrbBdpZVmduz+57lHrnxqZGIIqIIZbG0+OpweBIjcd+uTeCI6jUHL
JdNBozEoIs4w3sWcuoDpNRd8X++9YDGGTjFZenYbyecreCqNdRkGwADPiatuCU6BwDSda8ZIIqM0
vLuxSQT4+CXE0e2ql/laXegy7YbevZ0jSDxtK5qwnvzF2GQmQoSFsXfph+cgISdWwCuAqWlaFCQ+
hEHaZM7ImFN7SS2vP+N0EtPHtop0GjHKouSCHADP+lRA+KyYSm4Q2L2swRMBt5s5EYVFQ9YYy7IS
t7UtWkUGcR0ROASpHHxhF7feX1m+zaWGj/K+5qWJfg/cQGnIvdAVUp9oWEnZ++PLB0FloG83JpO6
IwbVbZwMtdfEMA0cZaGjOGGXt4yDXFLl6TlTQCb/1eg2BzjMMacNoGEcc+DKGynEwnzGKBUjNEkg
kU0r5ywywqXlhLevDeOtaF8eShXuD8rOGq1+Tt3W6hd95CXqygUXsIp0bzEkGeLEYBzPuSF8Nr8w
+5UZbUKxyMk1PhTCnZ+I3ThJBX+PmqvZX2C62uV5PsVyUNUm4gv4l0C2TukabTb4iZ4t0Bgex31Y
5gfgnPgBXJBh5ToePQaridgyVOKSQxyhVamOm+xl+E62qU7MrGhO9ieMYcM4IoCwmm1kQrn6FMUD
ow64LSVJ9SxTryIm40Miar5EhSHnFA+Kyl0sdvTh/+SO/Nr0HaU1Qm1qQgjTdNA2wWLsdzkZNSfg
UedrhWbRwBWjt95fuXNdmM1xSe/f4ixP/kzx8ZFh04oMuKLULZ8k3IwbVhjOFb9ptE2fqZ4mpUsg
FBBnY/c1tYqXZA4Ht/xSzXRGA/CnPVVqsu9VfQ+wSDDFJrez8i8COOBVMfxpd80CBlBEEYP5WCoU
1qj3AqMfx98BtE0EGYj0jRIk6hyNTDQiQTwx0WWlXkPth/WEJSQGVBULvN0UNB5hV9b3eOQ8YR2F
uRuFvtXJqWbNCyu3s+sp2DulBH0iFXSekpLSaMwH7scndSFHdjvWI+pbJvGPCX2R/b6kA7ZOtXHs
mLhLxezRAPmyM0OsiexIUWxpTUtWgdARXJrdqGsSgRU1J+56T6q9kelB1QhLsGJ1gUP9DYWKLf2G
vZ97d/DQIXMeZ1npUeLXblgdgTM0N6oFKNAXwRJprP5iAuMLT774RS5n+exUV5JMU/O5ISAWqZQE
f6lv+lom8UdX6YNEs8bASb7jnYgE6znxR+qrWwdSiR0YpJpdgFHxruBB9qMP3OMKXFLXgV3cK05/
P+1qsPtr+LMyY9f+X9K7CMj8jpU878ktuKByQWsYqIzSUDc78S7ii2Y4CrQ6PXDFiB53dQLfai75
+8yJEVqHDc2FvGU94r8NL7GKBR9gityYlN01/qXJqVDQu1J0mErrAMn+DqsHSsyN5P8GOikeSSjt
dgVPiyei6hyGR2WohclQGCYlADaskQwqLhsP+WSc5NVI6+4QB0X0SMEJGoNmnG+aLX5TIGiq19z8
MGZwp5bmF+QtjK9IHBq8CPpTJCaG10hL9vhNSE4mnMUPoNIPYJf2o5KZJU1wP3uhSpaTG7zrnFTo
tBDvGJ3RnUuGwCk+HzyvJM2TdIlXMH5kW9wqNZxRRnwNroIqSquiz+20XV02A5ERQd+yPQH5s26k
gMm/o9vK/IQ004tgkrrdshvdpPbCnLh/uPTRiqMen4wA0knGWVliC8hF2nEAEGq8Pt1/Cvv4OWr7
oLK+6lHeg3XP26Lrcu2DzaVfEDe6YTp1EMPOWiUMVMkkLM62o3ZVPm+kLr1bHLguuFCyHiRgNWBZ
UJ6vZN0yuUrzCKh/O7zk3XG335KoU39R4qOkLOeeU5zRQhh0YDpq6daA2oFK2OZ4dout/G7egY3g
F890cjBbCyzhscY2/J8wxJIBceyepg3VmMskC7+3IE7Clrh0Nr6kd7FktEHoKdkEF4RYGpxXOdwi
OWO5cANKnTGPAmb7XIbQNRIFduNl2rIPXJQGXH6TyXmJUFA0OfCl1FwouP0QmD3xRhpwIiVUsBId
gCZDJdsF5V6PbDX/SklXWYAq/NGgcIJAbKWZ28IKYSvF8Fi/d7ALel6Jen7tZxfn2tIyZ0aRabzD
NkN6Kt7Tk9EzwJZCMPGIY16XSlyV18kPYVIhLYVv9m6sTAbFPLzcJxUrTgIfvHMGCsSJa/YhcBsV
jd2MnAajGyE0KS+aTBNkx8rrsYygmkAS5MB9Ya947BXWburbbGKKY9qwbB0UJqkEVzDiGbwqx240
BSFVyVNih4vs/641s9Z9JZ1ikp5niAu1EBKQba0+0MqhmNeCAxnlr1/sWcLaXinLDeQo81jipWV1
rMPG79Dfhaf5902Wtooun9rMU7MluiecFMeegfY+KbqHfNUZNq4UuCNdGeGThL2v1tBSn8zOA19T
4nbTpoFp+9UbpXdZI7Dzs2Mg3lY4nMMm78e9++HmWgHT8s46WpuBIUSXfLdmkLFusm2MP1QXam0u
GD5MvdgJ2EJF2r4jUNJ8ViNO9Bsux2+T9A6tvxDzgpcF1gwCQdVwrKe6yy3iaRk8f+3ibvJvBcF7
oFqkxz+Dsk9evVzUZmjMmiQBc4TkkJncOVN1JE13rQ5XEP791LyBrPKWhOLhED8IhPAdH/RuAPcN
i/+EIQ4lrxlXfqv8t6CLfWMVP4RbGMkQE+lPFdnN8C444oSXDaELRYFWMrmi5OBXYqL3aM1Ig2zA
wD0mYg6WliiBVLLFMzwO5PU46flT31UnD6eHw5jD+nYNcQlg0IqKZgH01SIXzEAMDtc5gf/x95tG
HScPLz2y6tba1HWzUML1Z86jPGkVtspI9+ui33V7P78ItXeeqnpGIf7gss5ZaMJ0gQGnZ2sJRl1T
TIk6OS5D79+2GsUcrMsJLCbL57p4h54qgFzJix05x0chBLVz1vGxkxAwv/nQDDLdSDoXB+37q9aQ
bIyr85gVvTd5fSGKaOswvPcOx6IwXUGMWEaxXfPOF91hQOtfpPyBFjo5GvnC4cC1bmPc+42EtkxB
nbr5aeTUqds1zh5WTfs4Sbq8+2urnxBok2XO+f7FLrFRjupjCx9lx8Po5irR49elyxBlTYOak/KC
gs7QQrtNlVbHIQXrlOJVJBAIWrAFwxqZKtne03oC3/DcCP/H5xYbr5aFDA4Oq4ogf61bT6wV8a0M
kBU6Dy2smj/5jb2kvVuz6TxD7zYboB0Ur7ONjV7+z/MfTp1GaMNaEQjBx7wtyJPSxiRzN37YMGdw
CGKwSf3VSzaR9bJWi/gkBqF7hRmIM0Tjfsr+LA6FXEyj+aJgmRMeOoTgqZqBA5BJFwy4gS7OQFbJ
Wg4MGX1jvT1I/OgP4YMgn+8YI4P87HrKpSYeoi1mviLwSKcMeCLa8NsWHGwPgX/Dw87RtQq2qF76
A2F7bTXuUZ2ba0YGvUuCElCS67ppjgcU+rPr0MurlA4h8JrRBS1ncyBKh4Z7IMGiezN7p6+Yt9Wr
urotX2FEmpRt1UOQ7KCZsiEdPcT20p6/jmBKJq/Nt1TbujElWR13lya0Iv6UmIoNqEYymajdTfoL
Eo9dgmXVf1cztaTXu5aIWF3B5mDxBxLNHlcxjG1lwU18l1bqlxJCR0ITLmfOQnd6NH0s6KqXYBz2
fS7x5v14wTWb0rEE22n6jRfuTvf0o4PynVbC40zqfdM4gTmQZ6Hkn/xIytQmJBABorHDbaX4KCYm
xBCzkx8z77z4IIrtt7OgzmIhYpzyK8gxFMj5cgRxJIzDaWiA+IgnrXBJmExYGgZ9qq4cK8ZiA/cl
KfxvzqKpEdrNA1rcXnAbb83xvYq9popN1sDg2cXaPRjGShDJMTq5a2BaRDaPVC5YKEhXOndZazMr
5TR1oJ+DeRE0Xy24kSl7XMeYmUYTdGYsffiENJ3OiHcatGorRbMRbfOpRnYuYD8ENJe1LLF2mJ/D
/NstKzJ6TixoOmjG0FFzA6AtsxEvwzb0iY1jDK4NU1xY7P5cuBeJb9VXhRUEsVwrWepUrB2hFlPX
t/WGXj89+qQ/s8b/YlSMTOPSUHVVhuJu2A0/ihnW8A0+J/mkCC3GQUaKW36aknKlBh32qePCi71C
rrGRZ2u0fgT5iUNlNSdNEehlEPMTVNX3T+z/u4DKq+S00a8nigFzpsmSnbshdTymyIpBMJNkJ8Et
X4mL7dkffCrFv4YezSLUQLkJp/GYZn1pKHCjCtAIGmKfBSzgK5Q1UpAwaNvrR8UTicKQAy8QHn74
i3ZqbuVS/D6U/DLJ6CFdhf/E9nN2/h/6Dx/hJQMa8nLc9hztoojyr3620kKhF1Zmv2IFRm51W+19
n+FOW7JyM34EcUKe0Xd6kpMqsFx3X2RDhaE1FLQweEy/SJN2xlgoAzYB+UzOpyej/YVUX2QQZcih
kLe/fAhGEq3Lot9U4F3MUOhvis0ZPLV9/19sDJK/j6DZnmxW+SXj6Nl5YIKQcnyW7raPSru+wlVd
P9PH/oSxTsTo2fDTH4Kg2fluuRfwYWF+sUZTEZFL0TMgk8A4X+pjcsNwJ5EyrN8go1/vt1rnhqRB
G5Bv+to285PLIOiwhFqgdAiRMbLnR8DBNQaV9GVmeOaGet7a27hvycsracsyzWjkLt8VDzhZ6a9B
XDK2Bwuyb/0N5eY86LVX/A0syPyMJGJIVSG2axIqDhxL3utK4R09CKSmoqjsjUrvpoWUYLGgWQ36
Xxc8q86x1UtQvdj0LEa8jJqJMeYF5CN+WG8iqGTYakZQQmKEao3XaslHRoteQROSjjLFhFnxy1ZX
fVF5PhYqg/rrXn/6da75xUMiQzDeeRO9A19C3EIoiOqPgSThHCjYZP68MYd6ons6T5pCt/P+VRoJ
id6UKX4/QjBvfP8JPC/BHgK8d2I8lZxK/sUxq5IF7rr/H3MLMrvu4IfSjaVjMtkFghQXij3Pa+DE
p4rsVAqwYYg+K8iNqfSOEjTJy0yO8XDaJ89XysG+r7wVf/sZEmQsLnayGqFtGzWu5Z3U0Mk7U9N9
1qQ6jTyd6ovhCAyZ/zcbEsth7cel0eiLPnj4qLKIaztNsQpok4zZcjH9zmffqCIPFLKsDmNs46w0
ZJp3Rd/G/MtLG1XRmA58rAzb1Cn3dXG8WxyWexgA3Na+A0iQqubw6V08JKHrkbzQ0TyrjhaYTsIO
e4WdcQDhpZshodqd/PLOh7hdp1dGWcx/4hIX2ALU2903vRsZK/6ARUgRU+J3h4vHXK+WuG1ZJRd0
qAXoOCvBc3BTjSGfwx0gU02TP6wqK4PbXkUXDjo+xNfHDwIKOAxBDSR0wBUFRZF7HkV0VlTeqChy
8wsOt08MSjSX0bDOiT3uNVhWMDx09EmvmvCaDRVF1VVdOEDRc3xf0/tKv2NQ+5J4gKfFEDH+8CV6
LTAcDefDSn26dXnpzBIQEI2HQpQHwgtGtT+yC2YbO0t3lTNSJd1eIHAINJK+XFbFL/+jia0HaQRm
SU2pWQadYPX8ZR2rf0JPpFe1B0BEDZWjomsRka8SeNyoZqt2uyBBw86i+oT7EoLOjBbzYc6xHVjp
sXjeNmqqZnbTDOo3Tffj2Yrsv28Jp2Zxoq+ektnzKQUERtMZAkIjTLNfSim/2KVRPS1tZ49Ivt+g
cbuhW1W9kz+RxQeRbKHBMShMBemn1L4b0BoeRkZye4wEX8BfJfjL6ot9m2UOVh6HyO2rX9YLYgv7
bU2bccWEU7QxLxru7oEQT9iXARFdP2krpOK3kaFBxTZKrJQkAiOztznMHkuZJVlUWTJDHvmZx4K7
HaRc+piuuKXeoobBM/DfkbmbWNX0UpvtmaXaIQmwNcOlIDRAFpLolx5Z7/EPQcnQmg7Tsn/fblf6
POPEenqVZzpibyFlNbvZqmCGwbUxjPVKa7RKBtwbDzs5bqwv3D89H/ByAYZIa7pqgFzP1R2PlLYs
G9ciC3bQtdT4w9ehw8FKLN3Oaob/hcPyM3hiNGFsUA66GuQ14uFg7F1n+SZx/x5gLJgHMxDv8V7B
5uVZ+G1oz/XdM5/bk+K2j8DF1voT0FmrCMqdZbyyMU21ZEZWJae2X/gctOFAeohd/tqWTTKpoTlk
I1N9F4FXRZCUSgsyluAGlHtOCjOdLlgxgjSG003GG4aWrBvIv9GTeEKrV1GpNuhlEschXU7eryUU
QiqGd2aNCeqiUJxVenW2lftYjVEBKLbPbCExj0vtZ/N3kjXuNzvAeShwbbfP7YNw79Pr+jbux+aO
f31XVVDtyUtro/XBxy4lKv6A+LjD7h56iLA8nkzC0PkhL56dY2OUuKKjmt/yFc5ZVczs7xJrtgeB
st3PlEeIKthGU4jmwLlv5KAB4WYJPHVAmMYWc8rQbpGmQg7/bM3UnQHLBTfG41fIRJ9jR1rUUeA0
TpZ7swCWEi15khc/iyGj+nqKrV4fQULbxM7ZByaLPRsgeHasn1g4XZocY/xAq4Dbt81DOFsBVzk0
QyUpXoCBxjY/bkz0MMPlnOAL5uiMHFNhVbc0rE5zLHTR2O3zacMX+fk2LuHj/6MuMt16Av5rkAQw
4rHxCj7iv/4iVpd4HEyXAoVKbWOBDRqsAtqRwhy8DROj+V8JJY9o1gdjqV16/vcrHycpuwY+Zb55
UtiHH5XpRGyPSzIpHC3RGaD13znqpnLQ7imhHlmNQGvCFUgNVk7dQznMxmbu6Mm36rwOW5grn5vL
0ypO8M+vvvit3wNkXCezBzcTU0PRi0c3dWezIs3TUnd+GBFdqDuyZ6bweP/uZkrQfkWbSDQ5zy+c
eQvumiaVeFIjEjiJvDcd2Ub5vEBwThiAEWuAqEKGyEo6m3ttQ5CG+PPPQvS1rL7s9coeQs1JKMpC
7n6ewOMcTl4MryPxu/2Rjl1m/fIe/OX8y0/YCbJCnVgtTTnUdlQ0++ZWnXCxH9X8hz4gd3Cuuz16
isDFcJwKiY+E7GNp4zLVI0PQ+563vQlDHV8obI+vpxn6tpXcQ6FnhNV0FMpmocjyLIEsxx38rB9z
q5yIM3XXZ3LyjynQ0mayHbyiJ78P1nzFQqfZ7rjdXWts0lNx3aBcqrWyr8aUuKuh++wW6rHekAeG
OZSyG2jw/KdHbVFPE5fMPAPkiLqyBrjTs+lvsgYRDnMVUFyw3uZyjweiMAWLuVVguIAAW0rvf17y
/fY0nBPxkiHFVCGpoEbF+vxPqCbNmuAeKsSvbwRa7LjXkRMiDJriu+S/Ok4XJs/rIMpDJAEA6Tep
hh0Yd0k6kdi8CgBLGqWWrBFHNaHl+NCTqSAdRUuq85v/H3pi051Nmjbh9X6kb3lUJUywC/rhP5jd
TG/m+pP2uje1V8XNCrBR1dg5GdLHi8rjKBF+ZjY5YqULlQg+SMJK5Wa6qfO2ECMXUDPR4XBDJmAS
eYRI7ati+Fm6bPR40EXAQjRNdrlm5Habad+7MnZANwv7Aw2Ggacln9W9JQL5SKKl+ILLYhGX3uQi
xypgQCZFiqnokQytea5X1x+qnF17PvEi1oby62zNJvLdQ226tfLk1vBJgvN3p9UIISgr3phjxbkp
b+bYlcliCo267gF2XxN1keGaHVLBJJ2BwZ8nMDW2sZ5NaJuHNRq/QHVo6fdEF3LD9NBImrt8J2+f
nwGQ2NxGq8GDHyTbKos7mRl04acX+otbQi7sWNLjuPwJjdmgvWgoe3TknEJARIaX45L4eWRiWZnK
zco7lXJxk2BYk7MDGXFtmyvQrEiWNdHeDxkWzq4AD9zF9P7dRakIOE7FvPCROmNf4cYseIxmOuJA
bTMLj4BTHV4DrE/v+3V8+krMGpeZL9St+4NDzSI4NvDjb7qH8racSR7VKVOHoxyMpmfxwUlH2N+e
Rb2nYr6+NwP3VrbCu9VN8ivQ1Evxmm44pQscx/hyL4TbL4asv73NunYjjvKW7hPvgggchFbR66EE
wZAOr9zfmtQGrzmoAdvOZu3P7onRvqbnr2LZ3A63gkkfAjNIp+FvtNJmWSlc0Zpm7qBImVfIc2wv
XN0G5kZFa/xc/K94gmlB27lNsMkwhhe6bs6mxMtxednNGVjPsNI9qG8o/hqko2nQed50FNCy5FXD
+JncRcm+nWs1hryYxgcWdqDWeSFgM8Bs2N//q/0fRsExJBZrxjY8Ie57MDiDDHC7Tde7p9HHRiP/
pd4/oLZLbFBMM5QeQu1K8i1hzZjpqDT9VHlgRay3p+bzKmaD2Q12ATbnaKIgt+FGqXrG/JKxKgdF
fkMHKWFRr5XJLa6iMo6LRF+6DaSEpIUtHslAukMEzxmCtBdmooG4sBBLR3D966RkNzmFJMWFwPWx
5G7ipnG5TbEni4Bnag/epE8VeTAvu/aLEf3UIDts0Wfg/e+d6ox38d4NKdm3AKiKmiq4L0gwQp58
TMIkphNZ31ruVC0ISjIzNhTVqLUyHd01NUSBSFmKCJFyqa89+LZ3ane7Pou/hu9qFkj2mJCfaXQC
TbzC6afjBrJjPwAG3b3S3ilN8tf1oRPDcTNmjg5qaHkFcIOqyDUNG6ofUUISlGkOvYcg+WKRxIdr
+mt5FyVM3ObKXzRhc2wx6Y1hBzAV7gnq8IY+ICmsoTVRD/hDurWD6r9YYqIfIEN5L+yQh4NyQzTO
Pv2JRqORe9Cnx5JvlIa3afy0Izl5c8Sz7B3srZ5HsDl+tLOC8l/9pxq4ZF4cbru8ylrp8vAbsnpa
CGOH2h8xpl0Xr0/+7VvBEy82T/O+SMfJH1b4BOrIB40aGlAnW8hgJivV0EqiIqPRtK3qxl/sXOy2
zElRQjfvZmUrnKcPgPo5o+1eSd45Y98Gk4RICWrSOQP9vfe0lJIc5enTrfH8hsVwRT2GLtkGyxFx
3S3CDGghNrwmxE45dbh6UObaRj3JOJiC+/N2cy3vkOIlpl6nWy/10dyyMZKSHOvddCij5nrjOmt3
ZlR2fPnYXxCbSU/zM7y/oXnCxcxpTf6T4GNcluQAb/FbqvCbjr97Q38kfvnlZA6MOaQyYmQ6woza
3vbQcmZjBlItk+lSZ0hBR0Mdt/uS/JLqGV2pkSgjfg4howFkfSLp4y43uwtTskpInrpABviZgX4V
DrRwJ/6kmhH4uCUDJA6HKNiFPI4vvS/hNq3giQpx+hYHwdNxpJHGpSAH1+5zUS+AuHZJiiYCFx92
gQ1BXp8Z6n2eGpbaELWb2MErjPFJ4iPr8zj6C9KM7xNd3Jl8gDHkpfrde95fuh1KQxNAGFdHmVuI
XjQ4Fd56Ncxw/kGYkvpNKFvZajFfpKSshRSUz2w5EtkWD3B0mZSnQj7MSmWQfPRgwPxs0ukvKv1d
LpMCsfZuwPBi56dSxl1xFLyIedICiVFkIggPj+Za5IusrK51dbnMGRnua/lIA9LW/pHa56iFQyFE
KuMWALMgPc7DVJKVMnGxynqOj5Xny38keYfU5ldLAmPN6p5J41D8niORDZppU6oo+Qvz7g0XZH7B
GxYm89W9exFRh/URTM7+CuFLawA/Da/Id3kKKJM6HP87Dxn2eGvTM6bVe7kM82srMebYMeZIJmM+
viEMlsJx591yiFjnlCd3aZAj8X32x65rKtSJInKIw1KTgL2bMUDluHqEnwTA81JpK1BD6K50Djax
aQhiSappw5AMElOi9FFMjLhot9SJP/pUmTktDXZj5Baq7U5Ek68uApuOYmxCXdh5NtDVox+5qvx8
7H8jqJgkJZU4e9/VtB6tnWZF5YEmx1WjcUpOcLfXx3qxbzmmvzt4bKTldD1IVh2ooucT1h6zlWC1
/Z23qIP4Tmqi8VguVsk/cDhh7cbLA9GC6CYS4+8AFVnQajwZ9rAijsa21DF5B86neLsf1nvwFnZ8
6JFahlTrAE5IRde/P+I9lkAe5z0qNM9piSVC7uXJ5n71EJeYTL9nYWh36DbwSGPPP6qGWuPfnKKD
/b+nWHSwqZmDfwrhVg6cR4HW6Cs3iHYH9GOP9q+Kh+hFKWggKq8LjwlGJnriRjGGBt4izvfk/aUU
pTYTby0naVj+ZKmcqx9TPEP4sA1KjA92UtC8fppiapzDI8m/QoZnyCGDriupSBHs5CDBVpjL/RxQ
t+jfuU0idQZgvlZP652zdytRbVYfzNxUbjraCmgTZJ4OxJUgRRlDBj8BMFeO82KLla1da7tDLw5P
Q2qOABHNbVNCRlyffahcXfobo5wOzABMB0DDMWKPLZQwaz3gjt1r0J3klD5P5V9iO6/jpGzNYFzZ
2vImCCwQ9Z/UuWT0UD9jF1F20/CDxUiSFqueA8agH8n+qJu/ZowggXjMZI6Qvdr8cEl4yK0VLQHf
RTveDEN+mBYSM18D9Kont/H+mcJ4yYOTARjweD+0ubTTVkV9oPqbjykhRXMoC7eR4QYiY0FBiVhC
9h0lBhyQMB5JaOFi+xGfxoshrns78iSedSN5Nr1SURanh38RYd8RA6eT0c0+gceDMlgwcUFzU2Yp
CvZ429QPHKh8+1QmX5czNkL2GdoRCGFvIzzC2HmpMYOlSMoVHVMlH11OJu4K79naSv4gsx/siL6Z
5VpxXDtDMHOgGqESfrWZuk0+wYk/k/3Lf8HTz7F+JpWUtSu1eqeknCfe52XuoF4uzj1vocvkixTH
m7nd8eJmSaSqhi5h5OdDcW1zSxOPgzRTKqfJNKTj/f2fLt62UQ0Sg//UA8xumWh7k5K9piHM5RM7
XyZruQB3820zJLWeoDm8KBqIw3dCSQhLowN8O0k0kgk/MlPybLU43xVv2pRC2ucajIpa08oQTJPU
3PITACcegiP6WGmE4cy+hqr9Fbg1inJ+gq8TtKu20lyQYUwo1zisU0kGOpDc8VW5Aw0Tw/tl/tIc
IEpK2PZKiscOQXkFvXGg4Ntm1JD624RHl3qoQBG6pWo/B0Wi1tAPshaxoTaBE4Z0kEUs8UwZ8S4i
963Js5vH/6VqB6M6urNLIn5tvMSKN5T+2k2BcnB1bK5QVb/dsJJp6rBk76Ww9Eo2UE69rvvFCTx9
Uvd1VSYP1Fs5UrTCGnZQ6IgZQQVer7J4SDciNdHIVk1MahVoQB0YdP8LGhNHvbxq2cflaAhaoY6e
3pJhRNs/I4nen0POcIiNlAVpI+E7kt9XHJK4C6k2ChiwqTpKJF91v+LDUgXByfG5pq7WrZHpXpmW
j/lT7Ak3gCUcN8imU93hX/dgCHgrbyPU87LjYqLwmYNd5zJEh4F9imKRX0bG1Qt1HDi2qAZyX4Uq
mpLRSKSod7b7t9IboMJ6CBgsZvbht0I35Q2vaIrgiANbbbxotTEcDyp4hDPwqZ1qcWCoulx5CGNR
wxPOk3Y0qKDsZ22cbcbYQC6SE1q+S07JuAXdhntSL5v9KpKxQr0VY1Ay5Rm0eIok29LzBAybDqgg
6pRCBI0MHLCqcKmHz+eTN2aSfl0kfdcyRPKEIrl2wxa+lBNaIIypP8A+RiXG7HA+WzNu78FD/I1w
CkvcIdSs8+okcYakFDsmLP61zOj+iTB7VGNt46Ev7KeqHhG0UjuPO29MdJqNp+xMCrzY8tTJoIqL
oBlZV3BMVOKe/EEtQfYjnlfPnUGvxaAJr3UeDPJh03XFcR5W2fBf3UjAG+HbWTc+U229w2wxTFKs
BuvdJvr6K+bn+IW3CN2wEufESwz7RZh+nxb/dcG+aPdagJY1NepfOVJfVZl8K68LqY2L8DRUg8y9
Rh9L7uM+NTzqnXCRKRb4Fxn3i0guNc0g7ZsoE9nWBQghUzAJ8450hhLhgOplcfaYmoNSbgjz+k6U
ZlU2ED9oMnEhG+ij6QQ3xY0YEB+nG0MluYMHHMU+xrbg8+V7Nk+U8wwjP7RX3iBNAFGE1IR/zMpf
lX7/FciFey+K5NFH/+MAYVrp+yUxUAITbxVpJm1kQylLF/6LSVWG5/ynK5JSa6MlJA4UT3szkgaL
rHYwGY1hLUjqXqR+QnZ17F3Gux1j/adEY/rK3k2CK8BkPk6qDPJQUIJef+JGUnhITb6nadsweYBz
DJZKsG8HVDZ1uhCi8i6peecJEz5T2WJUD32N3aucUk9MiTp+U/Y4HPVGTXq8f76m86U+F5O86i2/
vjt2wwmwnHR2kfO37ZUh/7LnMhWIPBszq+QRmLSlk5pEBJyFDClf3WbBFPk/EnbYmavPwHSeW4IS
Hvnf1wuFf0ssHtKXDlamo2eGV/hy4IxuaqLO2ZPjBDsFng7gBvQoRwKugH+yVKRF5mBNCiKqUACH
G0G2CQxv3M6qenqbpFi9jwA2wtSF+OhndgD36qxNAqMsMwMQBNfmpcr9vgeMe6cgufO4qwoXBZt9
jC3gyIUBldMt0cEP6Y+VptUBIM87SE4yGflJbq5hUeOMbPM7/MXqE58e0jxidWSbtQys4fPJanxP
7pXF6nWOulV1AdRl/D7T2OiYHR1Hycy35R5DVU6yqT69Xyl3CrUpVL9UnZbNrMhLPx+/8q6R9wAq
8VNw6pV+gfw/p5GMoKxXG0PeE+9ZpWs660fY2yBPQiSiVzDcVRDELY70G8MlDmj8Pn/Mv+RG6NtT
RtP/mee6oXjaV9Ze/OgieDtIdVvbcNegqVzX+etINawr+vQTUGXK197jrhRKmGatZ549zBNLDWxk
tIqit4t+aMbrM9NqHNkMg9zwRsiIbf8HwMVWwP1E5eJN2ScJrS3GOm8BSgih9KCTfVZUtCWsYFEX
f7CB9hPOAFrDjn/yojhKNonbN72suzi5p43vLFSTzTuGAjfm6LlHtRry1fn3fS60P+iALIRdMdrM
OzMwDgVErKsyqd/yn9w7yqGYbEHHGRjEWHg5LlgXv3K1wgrt/DjTo6ZSVq8ZJWKFg5vWarM4dLZX
5HClG+YQ3QlTzMJoFTxqUmIMbtizgn09GZdHgYGkjuOkoIAMaJxi3TkqkhLJrC8lmaISEMpB/upK
Lg66B3Sp5qIUqTwFjfYPaZRt6BxTUIYhYOtnQuDNKea1ITfWnqq/hSKCCFRvtQf9vi5uaEiSX0Ei
y0ZgAAtdTYp1cBKrCO90lmUQ98FKqskkoBizDJoketBZOe5qsBxGbfUJ0rDdy3PNdyr7z/LvHv5t
pj/dPDjGxC6DvsXSpesyxYs0WXJ5Mauu1bieuC6rtM3UyAOb7u9V77NJQDHe133VQ814fo38iZNS
8GRzBqSZWoeyKI9BUB9yZQ9mAn84F2zBaLhYdaOHHtE8VliCKuUEZGgQ3HLGf5QUkDGedx9XEh8b
VKO9o1W+gZYnTLgT25wDiCddcoqRYua9o8LSjGxQFmRGuz9Xc3F8Pj7Abkzm5B/5uAvh+NDqsPAZ
oEKpZetcCaqgeQAVmr2Gr6jg3VKYyQZgbao2hQpqaOT2N1pK8ZhT07DIFnhNbF+OReD+dFDT1yTW
mb2glEEzIM5LNsUIMb6l/b7tvWYJb/xIUbxp13AIb3vyCvu9USa+4JzD9FXag+d5eh2ZO0689aIE
ofEbTxbgzHDK+ve6U4zuRkMK2S04DMeqW35WHgtRp6aVfqijglQNsiBN9MmXlljLvcacyF9M73VC
0LtwhYEWboUAT2KCXNd8YCYwsYb+W+CRtTJLqCb4b1zCWGN2+F+P7u9aO5FqJMW7ciIiulJnHEpU
JFEPls6GJCHN1TXjNiJS6loUBDWInWPhai1jQ2t4bfQSHcqH0Oleoa82cqReUQ7AvlQqWsmbL4+x
TsoGyxLGe/rtaOsYTC9t6t+bfq5bOy8JpPbgFqSQVCekt9OQV6UM1YCnRFZ96hhsAIbmy2uMr8bl
GJeebjYoE/slacI6nwMufd8IsLstuGu+0JKFS7GUv7pdg0GHASlQr6FeZOZIDVT2rw00pXXn/Faj
PpB4xc0ZYfSyu6LskLm/qmHerwbrBfkdkuExukFj7ZEpWYJ8er6U5yByFhqPyCrMNdyUGH8DnwS1
P42w8LbAhruMXNi6Lv13qX7avcuTv2k1X7pFHzqLoKavqdb7vQ1aQyDoxwDHdj9cHl3SD16pprKI
lUzy97jn91Luv5N7xLba/FcEruZp+xg82qUAXQbKnb87hB4xM7ChQXwgLRK6FVqPJF0Kyb33uEpa
0aA/ggntwgrp3o1gIdUFyuqbL8wQ3lkkqBVWQBgQJHIflHIelWkRa1oFfaJ+HXTLrOohkb5b0LFk
VwT16h/BZg2O6RIF+/4MDGXz4IPyV6pa+7S5tNhZGmF4jZtkFYhVkF49RDE4sklSq7oum8mEwa+L
EBSno62/7hxJdy+kiVmMFjw4cIW1B8JtZcSDG9uLSt3W/SfnkkV90EHPmPqawO0VhYbuZdOc3qbS
s5hOYRL4FyZWUwGmnDVlBRTteUOY/FeNs6bpmwxZS4B0o4EAR/YSkDnmQ7s8Bd4Af5MAnIjJcNHs
EOlASc54O7sITGVUAehAlwh6jLkZuYDh7fUNvPBp8cXG6shRu6hDBeu6GHVbRoimnGGd73B2VEop
DZcRs0Zn8zqGSwGyBEo87AzB4eTOFqa25n2PAjfbG/GQk11s+WgyAJocX185LfReQSbwceHKoHmV
Uqe0QshXb6+6KAWgPu2WElHT1uBbDwvA8csur0tBjM3JcLFdEe+c2q4MN8OIP2CErKfGpNK6Dzqf
wYilVBhr2f0BXdMVI6fQcilopdPLT58AjtlSVMpfGpIiTxRO8l3L4awh3DZ2rYHce8SSmzSnVH85
8swpzVMsluzjBRk+DNZyu4w6AyEpWGyQqotca3F5riAqf8oFIISNt7LtgWPIKwcUPfswZ1ZLehPU
z0nsN15tk50rmdr+1hpYF5ls/owDnkx9Y/VvYO/QI1N8m8FFKFNy9YQ4cKy1J5vpLR/8tisH6SnZ
PoGkMj0S7+6i+0gXl9FHzqid4yRkH+KjkK5iKtI6VeiDUB64VTB+I4lK9VBsHJaCVH1uXFwMp4lF
7+kRwRJBdeYTFxjgz4lWB/1dG+Uki++qJVlP/B8qeVjyr3PAp5BX2Wg3uvkaGbSxTbgD+4DUpgTU
+5v4qD3RLcba8anIPhy+n0ZIiq4Y91JGwXR+mxQcyRIpMfPhiAJGpedw1SKY3GxanOz9rtmMb6dZ
GIvR40F8aFNtcBq8gB9PSVXThTpq67DgziTMvJoq0pv5GyZc2i1lSkTAsj67CuI6mUSmvG9Bb8g6
rg11lArz4/mA48vEsKpK1MhaAT37YMtklN9u0OvdtFQGK6Clu8qw9BD+t9PMb9ecrruDdgsVJlxj
5YzNhoOCZbUYQCAHOgIOjUJDf9lPm68P9k5MO2Q2ifCoXQoIYn8uWReqYyOUssz+zH6i5e4KWFS1
lurTmCN3r8jgLbZmEKFhYl07vg0GLWbmPwal4ETQnpQw9OWb6VbQ+S3+6fTkEv4ODOcOjAvaul0V
VEcMH87pUJFtFK7c6ZjKUdSJrPz5H4UO0voRBjipcUPHLQLjc+T3qJzlfQg+1gzgCosYAepyi42t
r29K7TIPUDNcJhrZ6KSxvAMYOI53c5JxEmW8SpCXRFSaNoWHV3hMEWA4usef04Z6+ISv774cNsil
97PSDBdUzzxBuguSwSkxLcdRmRDqBHiqooqgZiwDvHCdy8cO6aRkzm+6FIBQZiAxrKXOJ2o8wpkq
/MD/3H3AfuZlyifw7Nmnxc5SCGfF6OXxcnms15eAaWmkEYxHjF4dFsTZx7k+kNuM+l1y/lsgxl0+
Z9bUUo5maW3HiLEYxzILvbFqoePX3fbW0ANtWdMtJJ2BatE6fdyiuvxL2bHReusyiNx4hu6vkCs8
Kknh4bC8sNHYrshMU4GOCWWbqYEjpyHBxSAI5y95Cm5TZzIMxdchygLEG2Oc3A2uG7yWQUQglREx
51N35QTtg3XVp2GTkTaDnqqE2vb7WVHQwkTnM8TaUtaS5MZQSKABgaiYCpyKYs2zvEOX8kyAUbQl
VD014IQTP0m8zistmljyQse+vWTHOs+WknWu4tjn5134Ak3imGsJKYavTG0QL7lpimHhApqM5fSr
cIjpebebRM9qlYI4N3XiP8tnYC0yEebBTuDLQI6EFeKaJPHhCXvJWDNbreGLaVPX6YHq4IxA/XRq
PvGs97pX44sP9ECw0or0DoiicutDtFDjXbdfrAdEoqRaYRrdFO+IQqLtkzigI3ECyicn9sznaG6X
J9BI9h1PU7rrgf5fkdMiSwaQM7+3SLICRRyIwGjNWrhuZBcYJORWeGx0C2L7aaXgAKLfg4YeqCcw
lzN+wuYUOuBbpk/CtA9o5EiaQyjfRUhKS2UjDCA3Ox+tlTos+2YX0FNPmzNfojTQhcmFnsdCoOwn
qbyW0mRpIZ+qs2FAlCIRDWQ5oxxhdPXD16pj/ePPHqWIN6xgkFZDPNr1p4HB6cUcraTJ+IaC9mU+
RGw7IPhjfIrr5TaPvSroK37ZetFjdS/meYFgRFuW/FwQ79Zfjya8Z3T00pFs5Ji87NpJw5VodByW
DbK4gsDWntnEjD5V2zxVMXuNleiT043XzYjGCk6mUEN9gxBpaTUrWYGjQQwMiCjsaeUfUhJPOWMC
jjMvgOdLm63SVAUMp5M6gIrs0U0hm/KJxwO+8KTL6t5CvVANw/gL+d1+rr/UH4MFiUJII68D/UuN
hbWx5s+GhpPaWyYZxrJXc1WhlRNH4zSZZKrlZgP5w7bZaELKdSGZYtNUo9Cy8Gpul5hmcdJcCVod
jmvTncjKtE0DkIYIomtBfaIP1PQjcAp3Tt4l5r1aeSP0q1h6nZjSpcgScCVVPkWoQNIRfPSuzDI8
flE2rCt1ChbBQPZnQqny7C4qEl9f2H2P/xExdD29NmChPNcO8NActlFev6sovIOm/u5Ox4ocJnXs
nN/TNF2bE9MiSp/rzicAy+QZvaEJdMFhaFbKaFISfYhoQF1bhNp+yHLCV3Ue77xpVBd1r2kXFn9j
vvrXN6wtJwNP8b7GvkOR2v85I/g+NQRuxKU/Bzta6VBzr5eyAX0U5v0U42k9hudj3e1aC/2+xj9g
nu8AJt6pXBSghjShdqIDzIHDx9fKkV2rYKuuSS6JMJklp/h7Ax2LWerQpbQA/1av6epSiGhVDqEK
hpjQqOedqYj6QGQ2xak5jzoUVKxLBH5+fc5e/7f6WUwGS/O+u7uThiDlN0vUHK9XyZxqIf1yHoUW
oFHUqP3TsxpTDuOPXhqEhRsGeEL+Gr3ndGDAyMayFCPhEDK1oRIhkVCEoiai6lp7Is3L1Wei3uqe
zPsqf4kY9RUn4ofN5KQ8NnOeq4Sp2Vx/bzi1NacuMFC+kCjvjrEYgBeTp+bY+/+hwYrzhJp6Wjob
7Nbz9PENxGWdW5UTGwJxJ3JeDko+RP9uPyTPtH64/ZPRrXvHESMcwK6DBX6Zeep/xUPWm3j8Qka1
qSpwlxzkcLOUEUI+Du5I8rzbR8YDYz7XVEynwoMRnk5sY28FVCRzJhQ2gMfxvOAUhq44/IBiroxO
YHGyyMlXBr+iY66ZREy5WWpbKbgpCuv2OkpONtsDDHMYnb6wPk358Q0mI1jriwHucSJvcrfotERA
GT3uPAy9H7QBAHY9jXJK/FyC2zYAYsWZw+Ksh2CQAhshwz7TZalv1Cl5ydGGSRy6s97KO6Q9XAvX
QwofP928ldsz98jAk5p1xN84pS1OIZAAs56DZR/g7xzN3ozkuODUFG0f3BkrTHD6YJdWOdN/WLbv
pC43FT8qMHSDMtjyFTwXVBb7XTIwZVmh7SdzIwMnLR3sW9wz5STDHktJtCj2C4A6ibFP8opo/D7i
bksAGiCCzdpbaVREvxPKBKSkEh0CQZK2sspOZIbotqB5hQMXgOsE+KUZaJazw/ufRqCX/k76doMt
YTz79QhjxjqVFOeMoVyr1aaZsUHx8Popn+V9D2We2LUfBGqUrMRY7kDPM1P9+PwURJG9H4jP4JOM
94sM9h+PPmFAeB8H58hZbcW04vuz4pzUSYG4e7sjdnR96ckOJqjEURXEgF3gzUrNL67lNik5N/wh
3IR1ocy4gNENftRAAwKCbVCaVfCNc6tGtzLE13AgR/+QnkpNgoczsZOO5Iy3TwR089Q0pcq3Woli
zlwExiwHD6mE/7a4VPIDUexm5UDC5g/Q3zwFefX9RWkSs6vILzHkK3HVzGb8GnVEMle9BGKKo9xP
a6jcr6WB80PDumQL/+nGZLsRxOp+lVsKk3ymBGCz224CJjwU6/QkWn1VzuQk8/XutqIoii5jWwwo
NXzZ0v0rAFyvO3jeVcs5VaMh8OvIIfwrDtLBfVd5uVxUPB1pwooYGUTP7bYUo/m8P6oNPf0EleAy
+sp3k2mNVqcwkf+5NTahEolweJCbQeSmMBcE3FDEd0IKnLzlkBAliz5nuCeVVB7GucDVOwjzHAhx
OPs1YCntZ9Es5eFc8YT8Wird9FbDXH3WC5NHi53PVZPCxYhBMzc/5nva90sFT2ynNC676VcnOAdF
4GFunFZW1J7GmWMqBYAZyLsx1H9OTqt9xyotfDhlN8k3HRvNqmdPvgVcsMsR0DPjz1qFrWwQUhFg
FTJMJuxVzBNJcCloizLljzkaF12qZ8/w/gywVivja70qFT3dOSAUSpOm2GzjiiAQ82yWuDbO6n0E
Z8RrTj4unIiVhbmtOzENDthOxpxfAFatBD1tvIo5NkBtSAHR/du2LCg4oiZXXITMYKggXTxNOJtA
ZJ24zZ9dJa15LboKb0dVx3BApuRa+MhOrJ6peV6NDe2CPSFsnjXmc4oGlgndpIc8w067gGAHa/FZ
Ods9nDyzPdz7Jez1aLbpHFuG/tkDOLwnHIb6rLp5Xfx5Z5nxcYADorkhgiogHW9FeXEidvXrkoQj
EYn6UcFbGC45QI9cLAUuPWGeYRwLHjzkIw8tpkH37+pFy9cwP9r1ya7wvb8RbBwqDjQL1D8fFsqK
l+WckF7UZ1Ub34y9VHq3d+9fg2C4TaDMU8zmg8EAg2O4sShgGVOw97jIMPS24oJ6Y/2k/jWbWuOd
AGErULwJYvMA6o06I0Jp/i8kV/hmuir/2OMkKFMewAxaeyRcQRYTKZs66AqOr6unzXdmoKFsQ4GJ
fUlJzmEIY91cfPMxnQ5GAcMZlH/YmjgV2JeYq0cfu9AYsWw64CW6M53tHopq5Oj04Gf4mlA4+P+f
kzP6vlrD1u1PEv5v0//nNG2ISSWzxyatKm+QVwPUigKMCXpscV2YflDbYJf5RHUgv3UT3G9SjeMK
VyEzRWg80eCYN64RbXeTKMY6ce0OGwDMHIA2xlROhxZsM3eZNFqJiMmE8udlN0kYeaYt6/06jJ7Z
sdZw/uobZ60uWzBvCzmfrDg3Q+VDLJHPKYiV9n9VVqL4rK1v92hnL+TlNgc1LN3KJmzNPc8TG4xU
VxHC5mw5KUlZSQcHVPHJIHLN/Wtx+wyXQ4JUJxPGQDIZfJZSRDWeINzBdm9GCC7eehJDk65CgOUb
Vk+8L4379W4aqTLepm+nYuBiswTFxFhZD8qwAmkXSxUhwr4PH6luOoMx2kru01lj+YWQ5AgNoyw4
XnxF8p1gY6xL3X5TSpGvDRa18f/W2NFKd/S1auxOkBhYuKeMPf6wTmms+z6P70UfTZRlyUn5fWOc
nXbwpGZ6ljfHrXsJTCI1KtBTtnw57G8Ca6wLjEYoj78c0+dzZUuXpY79gKriRluQkMvWOcUr8Viu
98R+SnNpTcIk8A1HoPiZdEJWjspRi6T6fi0gqyWVi9E3pxQstr3bGm2QXIb2p2U4hYQtRrVGgMLT
hpFfMbsGzmbugLV/xk890T2k7JzD939qJ54eeGo4ltCdcY8HMghl8Stdsj4xHup/58/id5FHrGGO
0RQjrtn9AHQwtjiB0ZI/2CGr2EAh2Ln+Az5HK8cmuN18e79f+oYHdu3hWfGcjGD9geEVFlhvgf7C
TJZWJxQSnLL1zvZVXUr8N05U3g2s6DFzOK/E9itIxel7GojNwZfkFG7xeTceK+wmu5x1gY9C4D7d
mZHx+WhRQjSrSZ5LXznIAF+cEHQfhqDZFuNBD6TUR3/Vw8WwKXIF+LnfZdX9TmlwL5nTJnU2wOL4
kv/hIkcH+PYPZSp+N4oLuRdfvfQ0vn8OTXYwtRrpbSn9eVGpaqOlx8wJQrSUOKJL9O6M/PzGMkMA
0G8xxEr0Ua2uuJoCmmw3UGQqbg24XulWj5qdlZBFZARhSlJP2gdYLi30jgQ7T2S+1ojOTmLd4n9Q
9YlngdSFU16VNM226pkEEQCc9pamzoKUZYIGH6sd+Ho4gAdKmj1QQ1eXNk9MU+RJZP6HUuaEG0uh
ADwMkgyzSQjbnz6weZbRpdt+kr7ImSXZfiA+EiO/MJQAPhmLd4th4qtzNDQ4iyEWbr1w+JTkPb6x
GT7ptoYsoa7SiGYwiVcUF5i+asq8gEwK1AYfgNMNyB/wYCkD83PbEuSYt9e44wjQ1akR6yCqt9Ns
euqknPaW1kRi2QwFE5pvnFdj5/88ROEGjSghtEtsz6SBEuvaKDmipQx+/VzC+KPGQoPRHzjQw/VC
GfQ/G5k+r3PTW5FQtPS1+KsVMUK03gSwATaFOzaPCjydftbN3iVGIikNRRoOOZMlB98B+YWwNQpO
DrJtFCTwNTUoWvzLtcpn2TKIhUuLLorLKuFxKoLFErGlRt0Tv7+PqjV4i+zNr1ID/EftrGgxE644
rsppGL/H57E3zJ5oYwMJIicWdbNgIsHAAwXshhYTXILh2X1CjaIbtGjPLLfOdg54my3OHy1l4tNM
ecyJ1oD+AGo2S2bi/LYdCU82s1JxDDiMG8FN850gGa7xfNXsgWEsskSfwCXBooIlo2c8S5R8WA1I
1iL2efa3ajw5lwmvU2WtZsau3RSZwDe3N1TyjwbxpBV783p1Ib8pk1cYCpZLumALONRGRvU9L3nQ
sYq7iA6GsRx+84dHVhXzeN0qoJolQG8JwnJGj0Y2Wm2zvNJn8Cd2Qt0AhlXgCwq0/nBK8xHnHyTd
6BFaX5XJxMGPMClY4zE7FNnEBXBk1gEXeDwRM6U5BbXnOZcHHqtxTZNSyFvL67/5VBJHDkilHuAv
TYwfwUHO7Tjt9oaU5airt5yh4dOl9+3A3SdYTy8+tdD/ftbeLfjl+X/R7Xi5HQ6AhdT3ASIukll+
xY0Ub229uzvL1e/dmXZkMTyXrETzEZ+bBaodi8LaR/uaVNnt3SXpELUPnRoa/nK8ntF9ngNUFbMZ
5HOB+Q1HAlCiu6V6S5Ru3HjlXJSPo9ybWxt54/sf9z7bNizoeWsdVkHL6IEVFuTISiFkS5H5ZkHd
VFHN5vztwesU8JtM1goId7hIyCzHxpcEHWTZlERYRdEW/UV5+XP5BIcquCevieX5AXP33qtBcRhi
CGiGqinqd6GTUr+Lfx0hiP04VttLzXvxrk9N5BwJNeVZxPH3BuKxgPsuSkqNlmgDtP/XTF5yONaV
6JlgJZuAblV9Xv0JKrSVMkGbZTIUoUoqBGelYA2+XS29rQsYSF470OMxclqX+mC/vS40Y8IkVO52
N+TZuxbUgs7cr+JR/4U2b9wehZDtndtTvZSQzjXTB5Hc30pne4Gd91Jtjfnkv5sm8bt9uML0PkM5
8iqmBv/ikzUaOFX5spMWRswqef6IojgEdeRKmIA6Z/bLEoeO92HSMXuDKVALJr9gQ86dJS6gD0ZS
AcmFricwgS58udEKptP6Wg2WOFRo7xdOy7L34Pj7s6+AeKi3VvK1aEkOEVvHo7PkPt6sZJrfzzcZ
CjIETK2GohuN7D48sWtkBexfGI74dQfozvhMDEGjnYmk7Z7y4FEl4smYfBGVsugkW0m5qVOW3Q3R
XbUbL9lOlemabbywBxCnS1ZcQBb6y0LHjwL7unkklTRVprcg0jZKBXhhkqCc+okdJcprlYgPIBVz
TWj9ZtKj3SaCith7udJS1WZ7D4+gBYPfs7O8OsTyP6MhqTELAnx6W/v31if6CFmN3TpET6g/MwnU
zJZNUKsQDIFQ7esm+VI0MICcsVqXs3ECZU/wnuany3Auv0XRF6IpkD2m3kU/02FLFJmxSSuVKc4g
OgN+g7ABo3DdjrY+XVMC8dSZI3MJ/PSfoPlTVmwD56s8S/54sFdXL8M4fpTwRplzikDJA75aUw4G
1PUBnZR8jLt8SHjLlwz65g5kP0nMKcv5iDWFnSm2xYg6X+ENId2AS7y+/aqTYhVE/P/kxo9TxqHQ
qhPOxHy1H2A1iJlaH8fepUJFxlAZZ0kBvwxYSEWvbOX4jJQcEovb8ft9Cws05uw7sO0brPETMn4B
ueOsJdCHqN8qhPJsdHoqh3RNcx1oDG7nxbxQPIvReclbcF4HW35uHwVbME5twFdOShJAElysxS/y
9rA6ZjEJ0WvBQ0L5FhvYcfVUf6anLcq1bgsP4JrsVr6tRHgGFvDSkDZXFsVGIEEAZjnI5YbfTIRk
BYZwW9+/QoUDiKMlU2iJW1ERBGFq2mE0bFiQ2onodgxyEdve3RTh1kbzjTgxsy14xJX/5Whogj9S
3HGC1cc5QqdBBqNJuDIc06KTbqFvQHIbWssW67HCwbXDubT2mHNUVh5kki3nneJCnBE5r/kLEBbU
1vSDyr1WLyUdlbOa/9Ho7bznjMbnwMNIXguvskaFOuvyTGRROThKMprTpg9kyArZHU3Nz1z5yyvy
fOLtQ6R7DmU0DxZKYoexFZpYVubNb/wfoJ4nIJngE2motcL9r7oIUkS2R8rLw/3Up6PMbWFIELGH
4j8mydp66/8kP98EPBu0J28qFUhN90sKRQQvp4HX6oUke4tKjHAAfmrfpjD3KVMkrPmvNmlUeKIk
XY3pY0R+bH5it7nYFBffuWAsMerBgskUECcaaILmbfhMNk6QUCojm44oCL4Rs1uhOfFPjVwExegP
+9O4g3jY7PXlBXx9BaJY/+FeCVRZ7H1a7saeGQxPrtrCzPXkEzWUcNe6IIER6XcJsy65Ou/81pKr
1i0Bq3tciDYFRTVu7h2BIgrllyK129ljt5j4+3jm1GQMBQHKIKQBf++dRFJ5Ikm5XCZZXj+9s53h
pOxZuLxspyq5b8pebEe+JdzlJyvOqSNYAZJpcZDRXzfwysk39fvsiT5Z4c8V1DEyOK/TlnHOB2JE
3K0yuY3u3TBAPZCInNa/B/Oyxli2iTxk3bTMO0gyzmJZSqX9qZI7tZ/rhiQwwBxiVSI4kFI3dfml
Zs4DXTPN/dIIxBNJBG4tyx3JwzP0pFyqtbjuD2D/EpUhrV2cJv7xTpPtvkQnWWY3bjQKEBIvDi5E
uxAXvGq7IdWz7b4kRYx88YPy/855ByR84K74TrZzP9g/FTxr1WToHnhei6Pj/j6juH7+6WdAjQR9
eNd4a7VM0WBQzaGeaqAIejPd5G2cDWkFeDUPWqX3ejBo2d9zPrYvJbjwT1ojoaOm5wUEngjYaakq
9Kk8LpXGZYJMkOwL8Lw/pP72kg8MdYeQ7N0XJwFq6JTJ94Ur7VuaoPrIemAq6JoTpqb5Miuu0+PH
/6US07W7a/wH/Yy3umrcYNnRwwHWQMI/YFbK8W2/N0q90jgFoG6OO2BxsvMMXujxrWdZRXNaB/Ak
GO7m2e3D4yuNNR75SAPm+d5WqoynBJq+tHjY7taPkVOknlMzbm0VWjexQIP4z5M+jq0kIIyC41f0
xEqpuFtBDCHyqMZPmV39iwCriY95ETCOiDg7POrDr1IOj5BhvGh2jWqjhRrocw8YzN9UlPy1Sjou
1IBB7zyYD/9scObGvgbYaBsCSv6VAffPRAnRTtohcb+M02ma9mSTTgaO2HGDwncDyk4PMUUOqgnO
4nHQMoCumgK/OOTQjOs6du2AgO3gd8gPPM70KAyPaJkNx5xZpyJkcCGpdcULbCQfusp+GGpapwvd
B6ngptXBqI539Ykuhqxu2NoL5KhwSQDFohSJvROZfcfV4pKUOTisSpanAEfnbod9rAN6c/pQiu0H
leBxn4fQywJNP2KePnJdm2ZhKwv0ETPcwbMDmPVKCexUXG71aNEy9eEvFEHc+ID9yEDg7q/02EWf
0wTaGdOGYno+/IUMEK2/cKjkZlPaIENnZ2u0XTVNgymJHeQNSacyT1oAcXtJHjKz4C3PEfLXMHlZ
4jNCuS2mlNIwwuiYKFPrAJCnTyijZM46LxNAGVPMeUeTRtMymuNG4nHH1LYX7zZmj2xsyhbamtRf
OAxiRw3/uP8ndVAAGqsup5kEZFSoNKvk3mjLbEeXEfJoGD7rP9Az7JzTA8v/H5hlfxDUxN/DArit
+MKhdZarwDq0NcyS2RYcDPEAqhQXvvAYngwrs3ZPidQzRWLJvQ6HVkcR5/BntK4x339O/o18sJLQ
dRGT5xbz0BKEQF/cWDCIlY3zmA6lNUV48sm2+NzZl1KVY+LTrCKCPUakkrB+kpRKppu9/LuUJ2DA
cCjd6ibAk0rJKnqF/M+/NVWorl66TUuG7AbJRwhpxqrIhF4mymzSZwtq9nCIx6bBAMzeVPXPs1li
4iAE9wGFWVn17ZUSJFLKzbmsgFB4KiUdglNzeXUTJy+RafOvpXWIIihFCK4fVIhjYs4IMpnUr5xq
imysu2jeVNWH040bzMJCCcgikvfZYpuhgI2Jubh5bkyXt9vwV8+I/NabM+8tPOrywWlzdaEvCjUx
M/k5cqSqoq/9RsDjxHJfBLJUheXtSHsRFyDmANN+DFRlOFJL6/OIatYdUiF26i4zVWur4uQgdw+d
gcv7gmDkNIUFI5TGeqYukQjmBT0DK0Z6ryA6AERbbYUlbOHmuCbm5CDSK4QcNYJoNiPbXKe0zxLb
7Lkh9DW+QXhqBrMnkiAVs1XWuSitpvTBYpZygE9cjcrpMlnv//QquqqfZhAF1rhA0kSFpY+yRMN5
Jn8EdjTK4wPIqPLqx2UfiHliiuI7vtgeGO5Zr8RVU7f1Omc5eUCNQfW2bhPyBqBJHehU5IMaLt+b
fMREd+Jngn+UR+3Y5xBc7WLkLiy0uAFxhZmzxhQw6NxWYUiKZhfpKo1x6GZggCRKBCR/Y/OMk+d9
YEPTqUhivaTjJMgEJoMvZdnvd+yXdJgvxEOEJWnE5YjJhpqxhG5/VSjWt09cB/EPWff4a5HJxH5f
RvNFCkDef29mOfiILmkLu28eIQzWlE/9ddv/7aRqD1nzLeWPPUKr55He7dfR5twHBu5OBnMaV9CB
EZRiNFBS9Qdh2sMFbqWdyn5Jz24DNaMnMjjE4zZ7X4a9snTHhT/03qD/Evc22ERdgGPPjc1RUUVa
k2J/XDbKJ62Ypjw2uOAixCW1icZCpDUvONXDwieHpDFEt74YPnPtS0yQbnFd2fkGcx3w2ISkmp13
ViiowNB2Zl7YA8j7DaPyTmXdBwtXNGHg9sUMue+Usvxo1ohA4lZWBPkpkbtv6eHa9zZaN+OZ0e8T
JVJiimeYSG2ooHbgQqa+UBONomOiMjDUZFHcMU2BTaLVgUidFsDezX89CEeLwsO2qmVB/wXKQK6/
m0bgW9rxWWhVIOQKKxpcrY9SEhMdgC3PjtEjNjsaF54wP9CXJlCGxkUA9VhlxfUCUZE3qAy/r7wT
sgLXFBDDsBvzu7N9Ffg8T+FzbtetVzbj2etW5eXR1HZOs0Y+xgijkT0Jc2XmDpedNxzpszsTiOCr
+iDOIbBQKqkLJibazNm+YHYqmfCMDVGsTSqaSdbZT0fJyMfx8TsKlbH0x9U8muBpE+eyN2uaZl8w
QyIYAOD6AzV15/Hyi8uVSXVGqXc7p1Lhchqz+qIw2E/sd9oMr6jpz2x7C4YAT7g7SWh1YvJGyA1u
KH1CtEbI9XskomctpScRYr8oiu4BhSwDg2E6Zsk2ShU9C/sA5M1JvqOeWL10RfHawwgQ2G6DKDVc
SpPKQcr+wSGsEMEuWNXDMe7yBUjiGgFyfCqhUqNRw5/9U3JoFgXBr2WeUvd8a/VaLlCLpM7aOda3
iUftVjTV8/OOG/zR8Gnzn6/EN0nMa6lR0fDk84kEMQbme/IPu6/j9eF4k2P/hngyCQ/a8qK7M4VE
ysicp3CaHD6MROiNtOWQkjQ2RlsMDKvmR6gcQKi/wlZ6XZpkKH8/3hFrfj9FHjbh5mK9anvwQ72X
cYeFW0aNW8wgbYi9PPYz3YFimsP0EX9lRyjaq+Qzs6y4MstHUm/tsdoNcXSxieM9QV9/3eFGWqqq
XfJeaAS5dbgn4LDj7wzz9PFKyb9oaNjKWFoRNCxodvAquc2hIRV5J+BgZwCljfC0lFRSUTZCwkoA
lETusSRU72/FhGzCeMkMpBJC8duHkobL2o3G/eGqnp31ijvQk0Vnc55glpBZVCXQ0Ohh3PLhvZuo
8bQ1E0JECdWIcenxEuSLiMeRjlDd6vcPjfBhnupI6tQY5WEOSYkhMRrmZjAndME/5PkZweo3ScE/
yTRMw1FeXHAAmY6qM3hFdwhqzvQ/75SCEK88LeY8XxSXxj4tQX3mCiXGux5/N5p2/HJ1OuGrr2jJ
hTpQf13/Ilw/3qvoej2jAG3ZOfsBc78KjT/zipUQldGg/aRn3V/Q4iyp+S8ouEzP2H+DLlsRKSkU
vy7oQmEekex/a6X4Fm6P0TJW4H50Zn7/t9T95/QcfLuy4Pjw79fJUBoouEJ9Fj1ObA90L+TVXwtV
8miRkpguED2hvRr8ddcI12odwPeZH72TJNO/b8hdtkb/V23iT7JZoqxWhkpThywdFW5OzUbiLkRv
iwPovU6CHtc0OIXct4oD0ox+2G30vEA0BzaahVCMRinluC82bPA0gM2KN1X/LUmzOq1MgDU/a3wX
8WjOPUSfHr1VJjKvN7XC94NIJSd5XaYmJUXDXBU07Yzzc0LJcdbHqwyLSXcslSznvFgpD8NMP2Jw
JwN/dWEbHWHRBPwibNaOrcXuty7HbT+rzuG9yHkFt3825QaKrMl8gcb/J2BdCWuCZqmnp8rbnSu4
9ZOgdDNu96P4BvHVbcVsEFwXt9TTYkReSuDHXllC5gxkVF9Irkdiv1hJ2GDyRghQ0qlINH6sCNDt
AXZmfuMFXpumm7Wu4lSAckF72wXR1v96eLsWf24s+1/+Y7B69t1xYO07xn4Lkv3yt5/uepPwwfTB
mYR6Ve6SUZqFiDSbxCRpZ+NxcyGYu+MpDzqk+4w3wmtjvPZz3gnxZVHbl+UfEWCw0bR8cCfaS3jV
Ta4yl13PmL7m1dvCunUlntQQZDhMRwqrsOrTCL0046uRlSoF1qTRJnbhaIlwJF2bWCvb7t8ne1XI
R4nanzu2T1z0SokTRV8PU9f3wcgxYs60/5TTuEIMeDaVW0dlih411yep+yOUKNzsfoY+iaqYDMcQ
fR/onwtU1Wx4s3p6anuro4IiqKt2n4dMgisD020KcfFG56PF+//Xa2a/rcMasLKsMwZHAzlNKKMq
ATw+ERpz18G9Uh/ZIdrgGg9COzbaqAjop/u3xnv5KnuQCWwxXUBdutIzlNIrVru0hxZKK0TU1WoY
yZ/RzXvrHJUJ1fDRzQKZBjdXdGKXgPo1buL9Eqm1j249xbGLQnOgqdz1egYvbLWGD4hdOlySB5Uh
5O1cZIEdGsUoL7fQ2jXENUureDZMP5W8zVg5+ir79Iq7v3y25m2hUc2SE3PVCavxLJcphx6+tnSg
hQX8KoRKdI0CTbVrlibdsFqpfyGRW1RktD+kHGQ/CFrpSLjEjhnwaEbaiWHc9TYWXyzkPsToFRiq
dGWnYM6rvsxvmKbk79oehjpr/Ipl1u0RRjlZ8oyoIGJgq8Q7C0+THTIxfJ/UCP12wlwHlRxaX/Bl
71pCMLnGtAmig9n8x4sZytESDgfLkShyswGiUmptMDOyPmihyd5PLqKjv94xdz6zkecCV1sSBgYY
JFN0LiK+CTIisbe1yJM9HDM6ghXdz8LhhNR5+5bNGeT1FuUqaHhdmOr5ZdOr1tMwI4te3lDH0rkq
jvtk7UmNaNNXhD4ReIpmxH47xDvUsIoZe+CcPR/VSeA3UiOrzZou57nMFdZvYs4dnjYbK5FQxfK5
HiNhSP9yLw5wmfdkeYQlti87UH38ae/nHXq1rFqW913+UFcTxJSiYzSI4RPzY03/80FtYkmIRV4P
ed6iCwC5G6zRgOhU4lKEh9Sibv+8UQBbVXDa5gHa0QDBO0Y/bZ6vn3dwqaNaRxEXeoCH6PwHdL2D
PQqOGZUGfKjs5PuMXyydH9iOfKkho+jyxsUXzlZdvbEQcqudra5nP6UwXORVZxPr0OvMT2MAQxST
Z7pEkdPQMu9W34jkE5kmTldOWlUrXW61q5ztRKDj7H8DWEss7J7W3x6/BvK1iLuYtXKSJUcNyMDp
erEx/LV2jZ2elKk2ZrbDdM44XTmrS98mwrYfLChSnpU5QqoHMdM1YLUUGOMlCsgQj+SYTkbM8pFD
61rX6S5TRXacWu8O7XsZGyLa1TkElv6a9v26X7fxA0klsK9mPknADzm8VqLb7XSN10AEwaFVgGPO
ptFHF4LU/Zwouh9p/1uS2ACPd3S+MdLW8FtK9SgrfedhJf7xeYsae4KnIRQseyA3Aaiav/5YTtj7
g/MsEIBlbaJBwYKrIqDEC9CkVcbqhXgs6LKQQBG/C0/p6XfeQo/OAsgeTLIQ20bYbcSQBOj5B6sy
pIoakLVSYozF7dqoWGeVm5x0oxwEqOwG6F94VnS/XN6KpDsbF0JTCxcCbckXWwLeFZf0rOmC2mj6
iMz+yxIkV4SE92jua+oRNI5jc/qTRyqeVyJBdDrifor3ZQKSOfvapXIPJiKW0ieavDp+FUCQHM2L
Wcbpn4dhjvmRR6ahTlT06qbGR9o7oLgSuhqOswY09tsQqjqnWCvToauctB7QQJp5/r14YxtvZPqw
AD15aGGP6Z0iT/zT0RRi8fOGu58WqEYJBud7T1UjeyRPlLsjjX2iZnrw5XfcCfcAMXFhlnXn/XJq
XiNeQKkR3lqf865MitsSeYFkf2+bN9aCdVUZYG6DXdbg8++UXpW5cjVzcZLuQIyALeRwwe+tkGgz
Q99b4sgl/P+U1kub7bVvuun9Il8g55z6cOCkRkP9q0aBFIZ49yGKgoNJbfJQWKh61P0U09Yt1lA6
zvXFdWUEDjl76T72c+1P31KBj9QkBVAsNmbbGrXuGJ5wIjE+v7asDRs+jo0Rqqbj/ICOuwdwh92T
imYv7HWvy+ZylRRLSOdAZqIGszr1/NAcx39ZImUaPWmsX6bp8lSzRHToMvMwI2LyPvn0EsEILGd/
95s+3PioqdcI7Zk0nuhKh9UacpF0/99rbdVhAq4xCZDK5lFcvtmT6G76V+JfsyHBEpBLTv3YInnB
8ZIF6GASvWkGZjpsftkP53Hsu3NnUvGA2B8gcOYbPArRrTOrkBlSdWgy1Qb/bNZzLwnUd4F8jfHe
7BAiJrQRwp5ie8igGWrxobhL199Z6pSmdmGQXnOQrTOVQnS4laOGnTgKDCZQ2t+JDE1/6C/hQ0Hi
Yg6sEsgKp4So0ATpdQtjOJKaIYpBU7w5f0ysCkUKJq00WoTq4twSNUEuYn9U3Odua8rtfBfDtkU8
2v4jH4TXIjgQ+qA+0H7d1DEof+nWmR2IHvco7ONt4mCjRFTjW28T35t15u5gP5zZLI6jhMsAc9tX
BwtPAjUBmPvD8TXUvmGU9suaWXTAgH96Bra+AzUhHu9t3CVXf9zVWdEFi7DEuJHfgQmjR7ZQIhcN
Nu6nwtBdax/zOu5XQqfDZn+IcePok+R//aLbbdlGMjlLJXw1a0WIiV1qQ71R7T4NvuXsyC0nDJ20
UVDVT90kfbnCFE1h2MWTjedGDS53uWdTcYt4qjKCtzbAvMLyhAjW43BK2lqAZRXhk5JqpWUt+Hvq
O9JJ0trnFYGs15POazKqM/okii17tEVq737vCSQ7pOHNNQEHir4RTOjy03N3dl4u5m7GeVqj7cKs
tJfWSJcVf8ofCxbj95mGcec6RKZlr4anhJoFlXS4VjsrOdLisLPKKe/fUAkHj5MzRjTSzHzqFNfG
eRAWN2leey4IJ+gvnGeVpw3SrPtw9L1Ydw/OY8MkJKpRZ/8xZBEKXbyLyQXMjT13HOAX4K2nMoqk
ZfkJJsK6XX3Jqeo8cmE9g0aSPfxRsevfNFWsVgqOI6mJ9+90RxSzUpt5eVH/V6iGHFfYA2bu4LO8
vwm+lAHIJY8csRGKYAeYNAz1NSn7aoa09nTADEoNOqqF60FWPqVkwqUbwEIXkQzCFFpaK992asP5
+Nr4jmUINm6cuWELjotbfywgx3YMYKBQFe4q7I4vBh1JTsJButp593mVE3pI4cMAIRe9dd5pt0GC
+G8eS8DGs9/RsfdoEX2RGdfa6aBuKJNY4JMtC1K68WbDPGDUw/gzHe0nPnVwCetD290IimMK2RxV
OFwExByKdLG+ZDqeoS4SxkJBM7oLfnc5hTbstaQeHRs3rNtrTknyYZ3UiZrBsuq4OeMlGKbX1RqY
YtmOOoqNkBICp4h7Uw0d5BllGC0yzUKvmE7xKIQNChCokUtEIwKnXGsP0XdYOwLxhSwx9tsLlHPZ
MnbspHGjIJ6o/6MwbaIWRpRTXRbMcz8fUDllFtGx0Mi94s4GtzrZx3azDoUuX9xjws3QVwjH6zpe
tHa5CsJj28C2hME36zyYYPjwQUtCwi5SIsa1ueItRz0b/7sG7KTZG/86bx0v/8XWWjPn9m9Y/0jw
1DcLO/0+6MrRCQeLz4p6uBBI75RvZspSTZMPLAUu/NTGiPUIOoCr3mnidDrJqRZhByXGSo0xXY93
v1KclelNzDjlyWXscrUAcNF16Hp4wsnmJxYRdkNpMAucK+5e031Ya4PtNf5SG14iiHyGK0j9NQr4
BEaPfk0voFjzBKV9xOBSicB4yTIQYlHcBXk0JVogjm9OlHnPwnpZhv/fYtQYYcyIGYAvCC5Fu3py
+B/3r8Gt8zb0hK7/QISTsfSUIyne34Wx4mGqKXWvKs/DgFizRh0GV32vwMc5XahG7GWNsY27OdLt
12fvj9QPzr5I3Caecbe+uhlCabR5ld+8YcLQuZHsHVnQVw4GIz3TgULEaSrBY08JmAvPv9kOB8Gw
7TFU9kcOEyYxGBMxzrHVKHEn2j8A7k8xiYzWq/UTP3VzBkTry3CQWlv3FNGTdAaU7nBD2vYzK0lC
G0sgUzRuH+2H/HFZqAo/Sy8jY7weIaOZIIlU6ZwjRhtHBo6qyVurs5Uex1PmJSnhIaZNftRbAaDv
nGO4XweStLDCEYioUnHn/vrLyTWHwgV/9BFX6wiiDLyI6jRl7dqYK1gOuK/eGjqF/HB62cag88Kw
fhpTvbe8cOpbvQLHXVYunt1xJuWQYvEwABMxct2XIMRASrKwDGCCL0DY8aG2zkqgB2KFfo3pRG9k
nA7BxF/qpXWqaPX5I+wI7wH1HL1ablT5b9mwm3npDZTil8HkxQtX2CFywXWmpL+6su0Ci8q1hTY+
jMYw84fsiwRPLs9QWY24G5ql0cU2wt29gVjmCncRV8S1HG/2piTXeQK8ftz67MFeNCuZA5nloaOK
RdtU6m5PEDWjHFRUZyacPFc3C7n6l8yUjsAYAXWhwDuhjoROv4V77cwe5lDK7T/S58bREF4mvG+9
OdNRWC2ZAl4GwBiwWiebsaQm+SWnh/CgiMtqVto9mPt+Hy6qxGcipmHBUfJsYsbrUPFCXoo0TV0H
O2g17/g4ovXVr9OSsLKoD8328bOscnLiY64N5N6wtFg834h00I2wHS8JUOsbJKlvA0r1vdVwaDOc
Dieq4J9CFLkPN/KjREpFO1/69FGAOynmXu5F8Elp7iPBEqNXpHVFX5aSnojMLU6dJ60bI0Oi4ATW
gWDn8ARAlo+Y8U2KD2DU+ug1CwComjKOHwsKNYvyRpNXopOeM78SwDUMMl+6vVq4E1wuc6CPNhTS
NWfMlpCkH90JP9hRKOryucM3upzKrYxjOesJTRVdzSW6GMjBPFq3Eu0wd5XBOqc/ArA3r/MR4qlz
8sbGj1UrPS1/3ap/Qa2/9YW/La4hOCVnj3LbihJDc5Rl35fzqj1SUE1p/ws5+40CyKI/qqd5XTg1
NnTY8Gn6lzptQSW3w66vTbZivZm3e/HpjTRpgkRRZfnYBmSOrLY5wfhMm5sf2NEb5DjyDLgmGdb1
lQF1JXoNxSnEnKdxx5f0i+VJ3M56TDjO2YgfYfDzt533P/1oa7+1BMvb1iX8NRML+XKXh/uhVZT+
XOhvTOJYCUbHKS6ObSujymF+kGDPQPNUD4srdZiMb7e3BbQnycKvmWb1I94NitFi9V2GDCyG/h5A
fiTbR1BWlNhIRcIXmPGIij9ZpfEZvI23MMBj0RKuFLQpgC+LtZz5a/rysWYNWN1M6vTFIkd/y7l8
Y9gCq35LIQDaZL9+rMxMsk8MlJ6JOhjYNOkMSJDSxnV1VHpOIMOt64yAiN3TGE2wi+lP0X+FkqQi
R2gScTdHtmkOR9guGAzxEcZnd+sQjj+Qr1UCu8KF3aPIQJqyutQnrLBO+Iby4Q+1x+WFiCwk55mx
sXLmg8cnfUcD8HHjGWGYLxtNOGKAVdowz6OKecppU09MedJcx6jznGiUu/Su57dWYCdDOjdPFWs9
iLBrVq21UQRD7kwtshvaIdtd0+i3+Hiq10dURYjqvI/7h7UT/QrKz7717zpABhQfuqPO1g1ge7E5
ItpH1/HBSMAk3IIwatfzR6XQRgXA3ucA7ZMEx6yrILuH2NxDx4l11i65rnjLt9VvSkEauKoq9jBp
H0L9L7KO10kp1r8VF7Vej786gbr7IzcB4H2+Un4YBdLTEN2VKmRcp9Q40TuJ6WG857/OvPGY4Ki4
YIDpTUTokvg1ylvNTu/HvABzVX0eK2L3e0vOXsPVXlVv5OFLCAyVWXAPqE3wTYuITwJHNSzL9u5+
HUDkJdrWgjZsq1fvHHQBLLVp2rnq1s8Yjh4JhAQveyk80G0bk28htluUeq4URzoLtKKwQGypmb6V
qxE0K8vgLO3r/pTQhUz/IoZ+aSmqczBdx6BVlPA3MSBV/HsLXuPvgcov9NdGf32GlwOumeH/osMl
sBODF9AQXmgN8sqB3xmU+39I4trCeUn64w661DwdoDkzFGTYyz1PobK8QKUdvw9IRZlKHMuZC6RE
BsL5IzQ7UdOSwEICfWZJ1mFeCZ1TEDo80U34h6szgKhOq3R1DKYxj65hsxYR4w7zRtJN969nUKWq
C+mxSBb58uaUdKGi9rzQlppBMnkEwpQjTsyilZQwxtcP3O7q/8UE5ybnorGlFXj/li0Tqk3P7oGm
uq1MZzAS8jJVvzaHloEljMumi/WoVV3+HW+z9mFIl45f1bJaURaFwP0aXQVJqkipkC4v8Wwe20JG
yRWkFkG2+2iAHYMeLCY+IC6re7SdYbP1/JWKke2ByYX+yPgomJ/8fIBeH2p0u1s6hcRrNX+az0aO
tZSvkgKD6K96kNFk8zVB9Q6/9qUoAbRZn7/wTEm5kr//PVcmKIC9teBHuIsgrLMgGq/gXGz3luQQ
6GnSXcXD5Dv2Ovlz7y4jHRF3CyNtj2Z7oCOOft94ubmweOm8rVbnPGN+/HvKNKtsr34aeSP1arPI
xgerBWwadO4q+4o0FcMnN7Dh3nMPG5YuX5n/tJ1nmxjBrGkB2d72AWByILShuIRs3JTyEg7xh5Wd
ZB1Ax+EGMiSozZripZDBnm3aC0GdVFTVycjA0UtkkSSqGW8unyZxsz7FBehnos9kzOgp6kKR1hVi
c5x36jZUYOo3rr+C773PwV77EYKteIiGDGuxm5VHtVOrVD7M7BQUxuOGbGysTTDk7TGThf/17cwp
E+SzJUS7JsbJRDFQExQo3FlrDT0DDgLUL8sWxLJ0/koWvi0ddazNJ1HBTq0mB0UH2iVMMlk6Lwno
Gy2861D94OfUjohreTJcrwlGG3/nhQtreyv67/4VzDISApEU7lOdFD+EP5eoQcr4W9jhmfUpcpDr
MmlGcJJTitSLU4lOmrk89q9qPBTWWuyE8SbRxeAX1ooWE4TXf/ITUddI7b+/yZgW4xvWhCxYGSSP
niLEMQztXsfEcc7PAuJ6YKk654WpM8w25mV8pq+6AqERaKln5B/h2/SDZJbZytAUEJ6dTF+DxZqY
yv9SG3E8/RX2irQSAM6zwLm94i805faahyeOKoGb/9y4gP1b8bnoNgvUVcQPz7J8wTxmAJwPciIG
nEOidb4uVPevL2Y1twOuTYnO5h71eztIv53bFQuSFdFT3tXkw83+AAiUWO9UvbLbbAeErjcpwxbw
hBMKPUfdNrCswJOZk5C7btZxDJEvn2I3I2QbtacheOplToAtJxTTsy++zFPl4+5zkED0f8EWEOQF
KugZUrj9GMHzxtszeKXYSA5mgZ3laMFqPiRHd91CEnZZFHJ6+GJGnud1IdkZfRH6qDnXhE6zfxAx
VKOiNSght45AblaybRdN+CVp3+OzprtnhH/J6Zda9OO3pbTkJVpymY9ADVCxCBnObpYlZ0LixiH/
o112+ypQ2gK6hfQBRECW+LCDrxnuqrOjm5PNvbW65JU9XzHpM0PUPLelu/T9QokY5mlUPYHbsxCy
oW/LBZgHwuz2couWmwv0/Z4NxKxdK+r9xyJbFXns1Zh2NXIfl3xWq1YWPYw2DSmrBFolIOZq5Et7
ZSmgOcWJIj433ligBO6JqfsR0Q5yju46FngqSSr3OPrhWP9RdvHIZJ+2ggplyDVTzqSeBOGvUngp
QNdKLCeMt7nORbs08ajp1+1ClsY4GXu/fti5ulB22OCPU7h4z1qG2ZoExbNpdIX+J37TrHO61xrk
O+Y/O3GdhAjrCiDPqSyJpSGe5m2hjzBngHfYgLx65wezOhOgrEQ4X7O9XERf+bLU380pIEB5kmMR
42m5OR5ZeQxy5KPqhKX7r0z1o5W5b9swt3Qg1pGWgmrPvOBLyQ74vmlc98tf7lz0pA5WBH7H7qoh
s08DiD0a6JGc3lsqzgHlRnCdd9jyGaoMu7O13kTDp06ZEsF8WftiqCfaXldBLziNnQh8H9by00Ji
aajt0j3QR35bqCT1ggzGbinaXI+ECLxTKcfsXYUVcTeM2nOdmnJBaDe1HuLWsEf6dhxDgsbKzgwM
4cBna6ewAhszEszywgxMP+Ca0nZFnGjpUy5BYayWYpf4bzzin1lMgvxVfsvgCL8EXMDlmJDKNoue
xf2oZeH3KtQpSjCDWuuQqi7WWH6zxF1z3e4L8FY8KwcqKPQUBikbFDrZFAjoJ/M12Vg8ZyJDfj2V
jLHLlZL/m6UV08OvBAUKv8wt6l1RZwM9RA7vDA66EPAbEwF42Lvee7FEPYvfXd+ZTLfkcm5ADHLL
aGQzLXxyVI2mzuJF/T4mPtipBGc4KA5WLoOwPwH04NajUY/1Aknze7GZaPWphWN4xV7nGEVooEJM
E4WetsElDNcKXzzuza871rZASiNrvYlOHhvtGBW8Nc5aSZCC8rrytIZjft1XIDxPNkrHatQD+sPL
H7O7p8VcspnyEv5TDPhmbYARUoeKb48kimHEfym6CVm78iJS6dZoRHIL6k+IeDYfFxzXYNXAZuWx
ImnMLwA1a+sZWT308DYInPj1kIW2d3/wSo4K6FvikZbd6hSP/RmtwjBvwi1wdqhWFSw5mUXqtD12
FVcghzARQEK9IgEz1Akt/qeSRpwuTOP/jS3h3gXx41wDap3ggwIVC/TzFPxoW5cwh3omqQcMUqZn
zv3M9pEvMdBysXYq3K+tG+o6VibInzDkE0K8wkn6A5mmriR36DlOjNmiDMGK8dn+iIhdPOo04ZT7
IiEzvDibqzPr31FJ7Nv8dn7lu+sXNvvj//zoRQz2ZKHzyR2MSxC24+/ZdRtVpwaHWFHcajQX4Sxe
okjQTn7aOGWoDvgyIDDBXo+BE6rmtc7DusxeEct4yLLvWUpwTJLpheTeUcPL+h0FjhEoYIRhx/Zw
OvbJJ24LzdPwNLhc4PXNbCGmAwlFCaOFvRNv/iBzJgpM6dyh20IdnZs6fzH8XtTUe89vNYcx/rqG
QGZJSGQ0i1E8Bhc2agLR4mkJCKnxtu3vTWQsiBYQmDntU+c+SiY4YqPR1j1YSnvLgVZxE0OAwIcz
gJjQI+KbblYYjC5+796Hlan+CBgUYoDfH2PJM7Yyjto4pGh+QUmegw1VIB7bEtIWT7qNNYmwJ+dr
AMfybV5vr7h8RPBEJXioA7Lpqodj/r95PJZthAKfZouHvfZgT5VuSQAuHkpFORe363KiuDGrsXS/
SejepSba8dYw89pjXQcIbCheKxsN7XZpD5Rg1CVucW3WRkucr+9xsA/SeI7q5WubPZoGTLua8T4l
0Lo+XyqV6haSxLP+Q7g/jKPVvIXKJ9zYMcSLNyjOY+9n2dPGivs3BI+1T013Cm+WWbh+VF3Ro4Cc
eJ1RcV332uJBzVW/lAkHa9R0ezVLUrl/GwSCGBf4VyGPr4dnRSZfm7tG5A2BRFFsiwYhB0ditFtx
Rro71mtE6QybKaDQqxRCSgkVkJemR4p2gulWjH4oaIBeU67/xu18Utmp+G1crhU3Foqoxx6AzI8z
T7K9Dgkr6HT1QYNuKljOPtJZrg90JHrJeCqteX0zK2ebkFPcKO2oRC5iDKE79oJhWaGfnVm2jyU0
TwpS1hjOmlAJHbrWtxy3+D5MyeX5JjK0Wdw+gVUd4CQFqTELx11KtmheRBN1Jnhd0eueVKB3PDQL
PfJ4nXYvDfk6YjP8JPE/ECGMaFQlY6kAYWwyp5BhZVtJYvVtqXg+t2n9s9iu4Ta5IVT/4srKTx9Z
9tuzVs/o4OU2c/D7sX2d4PKsf8N8i6pqxe19EohDnG5+o8PCFI0W06Z4FpQneeh4dhutWp42Oasj
JTY+czh/cGe5ROZ/vxhEX+zFfNKbJsqTzD5m5uYO+kf2BONOx0ed5tePM2NMuiy9xMp6PsGgGzMx
657A8/jbAsuhtm1zyj4ypIxxgdoNV74GWwiMiNkqHkYK9Il45aeP+0J0IGYAHyFtHoY1RGTNWs4p
YdA8y95RjIMi3jjmviKea5MBEhwv5ypWOKK9MsMLfr2GjZjs0LpF1gTHKs3Uim6ZaszpFHahDfJG
TtnQlnuCjQAwkq/Y8ym7Uie5leNkpj7Tasp9cnVjTym5i/ilfKxlhzDo5o3NRJvSfvM4i/HSaCW1
nkC/GrGTrbP7BIEdb6xym93jOn1KtK+XYINcLKqZCm2qMv19kRhWhfvq0eGqii5taUUKJMTKJ3px
VxAlugqJkmz4yuDtzo0AnP9ley1Fi1BTyiRLEpHNbgihVNl6IhcDg1iv96k7IGD3NhfmZmG1CHF0
6+dmpdwqifqHMzXKb7GGL157zTBHYq7DPsxUxOpOpp8uni9f2WB3lIK3gpKJw7U5bATOVUGJW90M
Wct0nZgPXmFQIZOR0iejYY1tM8buRgp0FdOFOhtglezP8QXzx+AtCZOTJFZNuXa/94yVyKvIMnSa
2Iu8RKNOEPKT+6cUpe6hGvH8QXFkbB1Cf3y/OlUUK9E14FSZ7fSXsA6GPfER2r44qoyNzNzhg1Dr
69+8y1ATmlyg4zLHwos7jJioRR8uI+h8pnifzzyu6uai9FvQiZgD9mgKF6i+stGF/h7G/K1brJVU
Fa9ibI3sJ5Ze05gDIytLYVaCZZ2vXUrnA4xMZml2QMc9NCZJKRSlFCEUdxZllfNqvshFtAFeWz8p
u43TEh3fSG6YgagG8e2N/zxrqnqljvm8bvvFXdZu2+3SvdaIQRRe9ubgEOcr9kFIqmxL9HOXteHW
jXA9z79MXxWQkJELYp7xOx2rJg/HKM8IQoB6upA6vlV6OMf8skYhn3VV7po+tWxrbDIJyURRFEYR
kisgSCKSjBHXZsuubicO7e127ti7jZZC3r8wINmnKwnD9Qs/kpV+jKyB1s9VPIXX2clKlWJ3D7o9
ZqKcexx8BAVSMqFNOXh16YRmKyetC985SWt1AK1g/Iq2nS3ce0BrebyOFP+WBu4CjchHQUKVXrD/
hhjRbTQFZSrLUBKyxyzzJi1utILc+51gZawKG29FVP3F1vruiyqqkiFhs/o9oQjSlKB3Jl7sadpm
/zflIhxGj7X+RmOsvbKHgFi1uGSC7DSXc37lKW3XaS0u19V2/FFGX1lQLnmxw33QdocYfcLAuv9v
7FThXhK/2pyCiBdeYoAiRRnES/PZ7Idb7p19kI34A4Au8kqlvJIrERW73RvIE5qsA9pJ1PHFsQDZ
UP3KZeLKpWPJF9DoNYHsdSDyxQF0IP/XusPpY9l8msd1uPNH3VuRvRFoacHpr5HeRtTendrM0B42
zGi4IQsvCwTbWW5n/z1Ls7wpEdz4aKI55+oF/OoPqEOZXaPA5XBgjx7rD2GiXs9PPEiYDSDohcEk
G9u+4uzYdL3gryt5mRlOZYv+kJpWZmPl9S0GImyU/m/l2orQ2rxmcMscJHTkna4RWRROXQ+ej9/3
fnl8ZketIJ1K4Yqs1fhHynZFgoLggm8LSJwhLDHZGcc7EFjRW1qsgJ5n+gDnzctq6CDKXwc/kFtT
a5PRhFUaVp8qJ3GbCcddAHwEDyQSLGrAI4lFToGDxUN3cvTld6cN5uWtmoFciwqUm7ncIG17fpwV
1LDaeYp1bwOpn6BZx4h/SRe4ZzrBmalludNllhYHvQiRNxVuO9n/19mpMOeS/vH+MI0Y36XpKSAr
F5WZYx/KVlN92QAIjoj/LPbrEMK4WEOLx3Wlx1teAOF3PTWocoxr2voAZDzv+s4urllfJKppVBES
Oc+jSyvaHKgeJqeqP6OyYlmyybrIIUnHLZTnghiq0dJgXNkiUzMqXzg6sp1Od7ZKNltBhsdRdfjD
XMYgnicjy0WdGEQSmH6NZTEHOx4gvlHymRgcrXN+d5lPMzzUY3rFmoaDrwWdqTjU+hA6HdV1oYvZ
ubH7miDyxzpfhYOIktDNbq+T06igx0bDCn79PAAmW4HXfIQb1csWROmjFXA7ALEu13vtejaicEYy
K0zVefjJlIsB8fqwXCqRmX7+sD2ntI/PAtyeSuc7nbc+YbnZmVTt6EsMWWvNahJ3mym3canIPlT8
JQinWf8xvUrKphcsUuUNFcB1VYwrPXcdvu+72Ajsa0OFKrhM2MnDisliovuqchIBtyAJ1UK0a+jp
4L1+UFkx0RO3LNO9T0Doa9Ggz5AvYJr90NfxRIIVcIuKZvOeBOJL/kfQfLZa8E5qbZNJ7lDFQc7A
SlAqfkDrK1wioJLwO6gLCFxjs2iH/5/khi86YUzvWailuy7MhWQvC4BGQ1CJiNhrhetLZcI9eixv
nq5ACRRRjdbPgINgecZbK8LDfL/4+8fxU7HInTvcnJwwEj1N/CS+rBV6cXsZoAmJomAEqBbzPDWK
P7fTmY4RZTazP18MCJAHBllTZberstrDSbB2A5eTZ06+sy/ZKYciF6EUsStiRq0QGIk8vhQVP7zD
ih+tzDnsB2mJmoW9Gyvy5I6pOJLMRVhAPqF97dSR4Yxf1jtflw7QckkwBGts8PNVvpkEvQu3uzS6
XLDHfqWhg/uR8Ad4iQK6oXpnK0neG7S4yGCnbvwf+Yww8qQww7ufz7TRWf69ydjhB5hVZ3oGKLpV
uSFx0H47BZhG7mHq3BHx5rLksKowgTjfZ6HRaZMz3hrmj0R7dMwzDDTpBCcjaai0hkRsfm0aTtEw
9mPneyyMQLb0A/wNescnxcOLcdxvEvfPAUlQi/YPnUEFTRM9s1K3yTZXscY2JE7pZL2rr7+K5rXS
hSt9c4T8G0/C7ve5dL0bfAir9C4MCOaAFETid30omXit+4rF7tKPnfkVzyHMigPSQ3qh3mlRsMfb
Ed0W2ZFMkqtQetbZjE/eoODykxF7n54pWhzc9cWAN6CaZsjFxYRJ5KdgqvreyhPc6wl7egvZtIgx
i2eMrRfUWYhH+FbIZ+fZgW6cq5hQrAyxZnH4mzoMa1eRuVXXSM1rz3ZR5Bt32VhHwwN1ciNbM8l0
UkvKexAIUnKcBFYlZ+qJef6DlnWMehGiXshxETVpFag0a+G8eMg4pTsyUvWZiYK6hQ3imqhy0DvP
Mn9sZp5V0MeF9lBzrqNhwUlePpkrIv/d9+YMyHXQh8kBePhBRI1QHLgCLmwZSRyE9TS+oZDRNzKB
P26BHPKnvISEtFsMHTbCVQOCd9OvmCWFnLyh6hxM0lmfjHYtPA6upGbkdOQMJDip3d7DrRu6nBaJ
78msu7BvjYMacl/3iI0pZ4isbOWX2QsradTuKLkXZcqPMyNhl87xOCLPCqI5gKH+so3lbdZLu4vH
QFvKv96cLODDynYrlOIdLRb29SBaa9qb1lmUf8aer7BYUGR52uqOasPdp0+u10Kj8fO7lZ8otXcG
d6533bR2WDh76JgO9pWCHhG/7kTd5wsaq1BSfGZLKcNfX0XcExmCVXisHgIJJ6clLILkAJXOONTS
ztjz1kJkWrN7ERSXAcxL7mPxiI96KNPf82RGhPtYlCBEmLVFxt+bwsOTZCqNkkh6vdWzOZv+/frV
eATtQcEsSy4seAKse7hNz9T241ets1x4OXTOFSYxj5/3t4Ubh6ATe8fmrx4ETeSwkW6d/5k3qzeW
nzMbwZYrvSFK/1swJXk4ls4DXAUZ3Mc0Y4WEC12w6BhiM0oq3Ux5mssjUD00+T8K9O0w7RsnxLTf
iH+MuYjsquGUJinYQI/rcGobdxkPlqbSTk9mAi87JM8gdHcAwRjSBAT+qTA7bu6f9XdSqP/heqT9
8uhMFqhdW2nQ3+GBRJECfno+mqKmzWICgHB9iNyYj9ZRA2Jph3QCU9iFtENTpVZGC20DAhJVW2VA
ohYSdyn/JscCN0cvgm25CTCcMS/uaTTrzyCWBRKN2o77jxUf661mHd8IpXmurySRGaJJ1reE4BJd
356hi/XHluYRnnTZd8SCYck0FPjtQ2MVTbvXkoZ9Ftk2tc4l3Qc5swDBqIc3AsU8TeB73o5QM4GK
14SM7wLzJmxFBqCc9UgNnkHFw1OEfgvP1zNGplzq6SL81kKnS9M+e5MramjPaaRoDQxubUUroQCH
UTcxNX92TRskT51Bw1Nn5NtcRYD2VxkDLkLaQYFUHYyTZUgeVsPytCXMXdT0A9IcRGj2wvg7/Pyd
Jq6WsVKODObyfLY6NhaqaE7iFiD8SraDYhQpqht7sG61L1O314oIzIOwBrbe9Cyqg+0qJvraKsuv
CKBJ101l2ywh97uXPzv9lGuJ6ZN5MHXoS8SC4WfKk3EwOnmfF8j4+V0iRGcEjwlJb8WyAAfQ60rr
YpT/7ZtUKahEe/50/qezWzdrqxDtMg6hfJJ6Ly0X/KBipnPIUAREO5njk58GAQkocDbJ/YFfSTB5
7OsVHRerCxWV/XPAlpCJGmyaeQsFyJ3KNdm3yfF87uu7aJNFuqOEMbO1ZnOk6Owtt6JZjIPM6KyF
80EHAoN2Gz8Yz0lKJqrif/DIfdTy1mJJSwARXYqT4AVJLvsV6a+/S9paKn7sywGFGVWfwPhTGoAZ
9p8Xc0vWiSmts0b1VKnqFmmhXTc0idYndxwxBd9RtRpVHE+2XZ3a40eaUFOqE6xKG9evZ40BL14n
TdofAfG/JohhdnpoyDz5T4VpPUMFzHeQ2DofSjm+TTsAp3d/wKu1JE0tvb+DcXOhYbFX70pgclY9
cVVldtl6L0YOK7bqnBd+hSLUscIhxYc1nCIbPlN3uxfR316ixRwZ+TwVJVIZzUaBYMPdtYP7Nhtr
N9i8V+U+6/n3wBgYZRUqR2s3kKCroTg4a0tIflu36Z0b9MJezoicT1cVGGQVsRLS1uexw0oiDMEX
dG5P4nO+n+RNRySuI04IcjPr8/uoPdLrNSVmUZffk0MHhQ/EuMgQ4lMsYOPtx8kqKvGfSKVFnlnI
n13oX7derbeZf9dBiPgp9WmlqZ6gLAEpJHbrFyGyEMV62lrMlTGmEMMw3fDJxbEIXgIL5vGx9QNV
l+1mdR8RY9jW0T2knuAwiqsA56mVOIlPuhVY5gTaMIPKsmEwh5HwHgSkuEl4Zoqvf6oP+L1Veg7n
zHWGrPKfhG+jqZESK2JzQo/p4/NGyD/sSRy/3XWvhBzOxwoyOT5K7no1EPJ2u0Bh8QJfpT70mocJ
AK51HzkviPyfpEUNQsd7KfEsd89oqoBdzBs7vCrpU5Hu8hWldea16sQdnGO+ObSWUnwfWm+CvX9H
3DzbWS8qE3OZV4Zt71AJ80FUOnkHntPvnADc5LmMEyV2wHw2Xw7zJxmsaVN+YQjaCaW+9zbbO/pK
g8AAuU/vXKBOYKwN3pQkafhUzLX5waHjbcnlpqoTWT2spkq81TKj2VAfKozcD8caiuum4/kQX7rJ
MZofyOTeaJQnP2hFyLukM/uTdUTV5IMoMoEBLupxljco0oZpjlN4BJsvWBOZtifyDKC9Os3Bgxcv
k0IAVV/9e3jvGXIQS54QqFONO6kg/DmxWg01CNS1Ugd2HVjJnMBhOB99uC73YR9LBrYl3natD9oR
BxQ6QGYdAuWidUWV8t5pZwTYW6+pZOo43SqV2rLEOgWKCEqyqD2T78h9wsSqjNn8KSRI5MPpGzaP
YRp9Nb3LlnRyIOEd0UVRX/oyXwyluKW91hzwGFO54JbMBOR2Ce7vCIhjk2wqx5sJpQ40pzvwQHc7
hngbsIvGz68GuSt+QDswakAYJHvYXF0JmHYqKcKTug5GOTuUxlq4X1odQhLyhfzjGskzWnY23DPM
eCBWM8V218LcFS5Wlm/CwakdqEpzQV1R7WJTJkV96KF/8JOhO8tLDsA9hQ3lIljK616SFI1SUVaD
CwRh+4FpD/kjU1cOCXfNXdr6KfTCMBg2SnHjtgSVQQHzOpnCEtHiM2j8zwrLmyG3wPOdEEOqnEr7
NrlCYxmJLx6jIQT7PLp6s46AS2PP8LQGoZ/pvnYxroBboflygqP37xqDydj2T3G7uc7UhSXU6PyP
SBWPBrQ+jyE8SWr+oT6Cl7aeqHebHZtFQth1sME5XhF0IUiRNTZ3QqgOXD/LFymCOiv99wXlS5Ey
cJVAQkGxeANftezY4HSjmyekajyGbKt0RRoqjDyHlHg8K6animzH93TYHFfygVcoNr5isWgDVQdV
jxLfkidbyRpTO+FM8vo9+yfvlU6GYl9+yKvfUph7kzpR8zq26c9e6fr9Cbas8rkqYqLuVit1OfBx
4yMPe3QOfPxjGLCgeLLXq6jrF9JV5xrY/bDAZZMq/WXEYifEo0rXEuYi4ItbflQU5LnzeV58zoIa
scOAMRJTduDD0EnEd+2WILjZN8D51rZDWLb/RjE0ixX54R+vVGBVWQS+sT9jyEo1oPuudE0hTnAs
a8iyA1FK7ShOdgSo/TnTxA08epY5eh4BR/cx+n42rLXyyD8EA83yL3JamiIa7W8NjhjE7gwTYEQ9
KuuXFQGwnZ4xm6Tv1197l8uHeayomC5iOJRSVt+VovIwVOb8cBAZSLGVSy1XvzMSUxB8ynbqOObp
b/HV87ApFQi76VHYPo7j5P8OGGFSkWDY75K1T/EgJx4qCIGcgZJG9e/cUOdX0XbxexI1NnLQ2KyF
J3JJhIUoGBqAFDW70JUgzDFHGgj59qheDWQyLkugLn71JUJZMFL1Ovt04AwvBRTb1/Vg6xpgkZx3
j/CjReQ/QcBsExIz+L/TrQxUUMJk5VFl4WfYzBo1ohX+mjkywH5owg7FKllMNvIqybF+dHzS7U1S
3LsDHB8+fLlGr+2ReUCcmyO0jzvvDgezzFVjfekSDlNmSHNxj+xrq95DjNndQ1/58/h7V27z8Lec
32flYA9zVzyAMbyveC/HAM0w39h2sNXKOPkEqa5bMCdtCxeoM+nfEWykqA3xnCHgDseutyLRCzJU
LA3AqF4GeOfC70StmREPW7e7K/iv/QmUzk020GulWXSzBP2po6nP1fUElf3SdoX9RzUHAcfqlvT3
qkV+qKtCLXxFkuXIjjY7pRZ6CVsIB8iIuZoOS9T8ijLaH2vFoKbzRldFUaChJQ5aTihTorHYXcaN
MjMR9OkndUx3TeHfvZlpS/xxT5QjTCHdX3aMRuPM5Q0l9QCX/CYWVeGteHaSupnasarj9J+L5C8e
2Riy7GjQ6NryVqwvfUlM4rk9FT3uIVDl9SNbCQEQe0mWNYAQEpB4tDypCSlYTvrq59YMoMO1Rj+6
c8pOQDpMOdc5p322UF+20PH7PTyA9rpJGeZ3S2Eem87KANcpCjRUe1TeZj2TnawaMc+ZRxMTvWzY
fdJFKIj235wd+H8LnmiTb3FKtiaR5Y0ChDG3/H/d9RAkeKXSX8dOYb/5MRHaJXm6QEw6B3NEPME4
eWQVpIS9YIYOII46B/YgzWsaoTNjs6HUldCCnBWS3XAAhB6l7KVB3kZ/ENzNfash75kC6lyH+owT
3mvNqXbTfubdBZXsti5caRoGUxg7YihkW/v9luUeLR/tE//9SFI7Ch0tVPxrVupUj8beWjrjMlFZ
3LVkUg9DmUxUXOVGW/3vmU2fV7UwO5NtarRpRX9CeDjnOuvJ2aKa4ADS1Yb9YcJEYis7QT9dCPvd
uKHVVemfNO9f87LKNKNsX9NcxWWFYc4lvnb/tzm9LS5CmIhT8GS+tXtOxW8QZaSG0BsCOdlOAfk7
ELJ41kbS1frQl0GHgwnATxCrSZWxsuHNZP17EyFzlkEsW5F5VjoIjTJbY/uhbNWWdh27ZAjSPnw1
ZCzjMrUoewPohiY2gv9I9eES4ND7m9voJ+Y6mh4587ZvsUdW++G3P+mR59cnk7Kfjdn0hSnCrLj8
Mtq3mbZ1rT2/zwzSr/hOYa4F1E9BiefRy0lfKgCjYsFfRegWWVy4R5xdgzbQXh2+Hx0ZGp1nGeMp
qnqVctCtHsAJHwqpusP84VNkPt6P3zULJDh9+hjLbQY7L+RgXuKiD8PzfZM4hJrhW8HaYFzycIoX
5f5pMryYZeBaZ11JHnh1rH2SaX3J6FbxG0oO5HyGYyK6J3ghv/UyPuEf+wtUk12dPooHuN6ognvX
ew7PQlGxb+KpVPLhv35MmrsK4gj0OloPOxD4JVedkf5lW3BCsyYYklSu7Fn1qzYeDEMmXxuGrPLn
4wXgVH4NqpFz5IU7gulgWKmvlLrOnvFZlihcxLgxhdXrvITvfvgygYAQkC28PsyQztqJLuhuQeUL
zXiLGeHdmWClVOTgUTGYnJT5l4em7YXKBa4BeYAO6/sz19vxfaSZ2aF2KirSkK+5bagw2Gkipa67
Hrh6e0XxGXUSZyWPA6wrS/Q2u1aLj3i55vCrScX5MpaF3Hcq49IMloofxB8rMEtYOrPhfllC2lVh
DuI6KiXP2sW3f4YK8/qUCeS1FXvEZnGH+8hYLSB+q4SZlLGZkkJ3tY+tqcjcq7UxsbSIgws9kytK
ejhpQcYKJwPw1pqBAhS2BIPpWu6X/CCS+a5mnr2LrO9EogFD8Gpt/7teGOBlM9p1TrenR5iLXMbj
TVUPK8trhtxJWrRuF5LmsLwvGhIUaYYTPI1T1TehqtubCTxh9NFJWqP+VT4FFi3pgZy3+jz1Zwn1
cwiex71j9bf47Mw1TNRJml8n4q/jVuhwoCVCg+jH4u+ug00OVEbfb3WFIQnrClWJ9dyj8bYg709j
dNnIqvirmpeAOTE+F2HedgGHJC2yo6J4fF2l1ztH4JuvBR6NYRMV6LzS2YQCCSw1B5CkbC8xI11x
5jBe/yGN3l0sbDoRD2gfq4QGhzHTZkXKsdKRY+lG41SHe6/G2gfLzYUrsv9coutW8kuQTb/GBC6U
gXmHWWBeTLLeZQ23rUpK32OAi/6emtL4pzrxoA5Wr4MR6QxmGEG3jBkeXFUpcAIp9rKkbYJv4csR
zgB2zrauS/Rw1sGNng/IkY13OCM61szuraMmOobQ3tl74PTStggRJaEbmhTT2mh4oYF0eJB8EeW2
/jP+HurV2gb7CXqD1zs6fZpUe05Mh3UyF3sipI3jbQzxzTdwTzch2mdu5UThMA/wcBywIo0Gl2j0
3IqsWHKXRYDuGkVG2ocYua19S1y/q8T72o7SATwgMiHMqFPx626d24UXrB6xB7uhFfvb15i94U4e
hB35jXfXjVZ5Fqh+fOo42YAJnzQxSFJm4uiHIc/FHr+ClH0fPwp6ay35utnrA3k+3j9Sujb4e1dq
V35ibbP3X9cojJxzVErfkbir9/pIXMu6duyduZuhkYCwn52N1YUULn1rjr4OmXNAQKzPyobPpiCI
f4xMKU5ZFsl0aBT19sNvph6Ptrzxkw2gWTQR+lyjKd9SE0TL5qaF3q5z56w8jVlDx5bNO6BPS4Pu
64udFg9knnOXmefXoJap1XRDFyRc+30/8avTB/5z04bvN3d7AfbBmrwczX7ckO1QLAOf1FP63gIB
6U1Tj4EDw589ITfugMXmgQr8s49EtAaRJVsllNyLtE9e3aITR4faXGJzqNrbRz3QQUvnfZoS3/r1
kTYcOKXMliNQIV7QWwyZmQQqTowWJ55P0RzQmDOVAzd3QxjUYXKX52MjvvsyaothYmd24M3RB9YT
0d8XAWXgx/MkvbqzbM5Sf+WWQdyn94y1+pnw2TzFexIU10AOosK/5bZdb824+7/mwEvKTHFe8oEq
Hy8icAsmm8N9qCahT5roSwvwrvmPcWH4JOb9EcnBNPxEetKfAFkyoK/2senegrgYQZFBwg+rGidN
4yMJJvaiAZGbVvXwEmeySW800lq1flEwyKyWvs+njTigtf73mb7ztbd80nHzq+8Uyyg9I6GhNppy
vB2AVFz4yEoUmtZef+laLprUxbZpqNZR4tbkRXpxY0TzqvvMj5ntnxjZx4Z4u+lX2V6u8DX5DXR8
9VzKWu4pGPZk5A8JPxTxXgN1LlmNl6lxDWl8kdXlyXtDMP8YsTKWVZZtAXtVu9Sqlwh7xisXz5pi
hqcCjcGKsVT/QvZtDhCKcpzkmHrOuGCHIDtJn59Y43MHJnS2NDtsHL6zd5/TgmJBHcRPJuqf70CY
3nZGMOkgWGQU5wE4YWnqyX7XNQiOOqp77BivTh41R7hXoGlvf2RCBKBm5UehGG/Xeb4Prt3wx2tL
w7NbkPirKaOSEt+ZJlsFE8HVoBaEKnbG8D/yPhKB9eDTdmTUrecwfiHFkhbwgriNRDjokQLPB5UK
KH+NRlAooRXmAp/czgGQcriLeIMAQ8/Eb2KlApjRR9qUO1qPtJL0RYgR5lhI/5nSKOCefobkZbzO
2XvsIodwOfRtI0z+3UofT8ZwfvE0sfoY1WA1UX4DILeSviDOSpHc4iBySVNVarTDqBDhGnOFP5rZ
7QbUyTNCVBsRcRkV20D7t2ktgdUDHa8ElWhHFr6v5RhBqu4zQtV1mJ7E0hp/NXqjCO2uHmZ956TH
WWl0Q7EscTEWALryt2fzi3iS+qsf6hVLZyN8KcuN1kY6pzGooSWl4HnaW5A/GP/FRWEIm2CkGAsG
R/Pby51hr419DHZNGEqfFIvNh8Zt1qURxg0Q8RHDENSNdgzC3q2dgBFOpheJQZxG2D1C4m02bg2k
l5kE2vdVhrm/tB9NN9e3+oVLmBWEElo00RHjoMmzYcBsvDeGRMh7xzw9MIyd0eJEKRtVLQapwbW2
lCHJJPGmDCDrzCeYCKLS+xQL4cBuoqf+wG8t3FmnrfYbhnAICaPTcAmCLEjiuVWoFN2CoUI91hPm
EHENI+bHYEgNMlxgw1ddDDwT5NbpesK53+MYaZbotZ9OISmFvyXI8CM1IzuPP9LOn/eWOE69U+43
2anC7/Z6PjuLGn8R7jFSUsxePCv+GwS2EO9oyYpGyFrJrO5qvOuRgDtORL4zvtMgBQnO343ekG1p
ElkFxKvHEYPdDbbXKB56nWAVlTIR0todtEUUNCFRjdctVTsYbNL/lxw2NT6NoAacvxthq5xO+VoZ
slGiOsGOpNA+/9/fxVQygFyvOC4sVFqAFN/uJfnV/acvfv+/XFwuKghbf9FTHzwpxMPvbQ9V+/Fz
BnXBf42QmOIRpH8WeSiPKP7GJr7MkMNjdgpfrhxU7UaW75NYO+7+IuaaqYpiRUkKoRuTzl0/rCWp
lbhNb+QA9pBRUIJ6l4BBvaUzqnDqexhoBSaQxIpOzwz+JrqsvwEo/2zggpuzHMdwBsU5oLOMQCyg
Qt6byb8z+fp8BiQBoSGhcEzUXAPotoSuvPavkgkYyyzuP81gJUOJ3Ttx1E+lz+zYhiOS1MXRnJFF
0JcOQ1XaXrYgL7iJb7iES0WJxebCYpWXz9VtmKxhC6Gdjt2aRFCIIHszwaVie6hVM9aCjj+tELtz
9XDXrYvKBdOoOHhvlLMIhjWZf+GNg72ySlVTShrk0f4yX6u9Jl6ar2ORUipl4mPaB1lfJf2U7uPF
7JK62Gg2+vrYLI5pH3cZighe7ZWKfHDoLqxBSh26/k9UxQ5iVsh6lRu/FIXx89wvsx/NOvQq+yil
qIsc7BwFeYkURHPzelqX91zKkivxnkuHXU21Fv2Q7GhxHBvV0xc1ARR/YSkTJC75auYHfI67TZOB
BTn8LqmL5U9WPqmErGpZ6DhCIO3b5KbYqH3Ljzk8bpkffaBQUkKZqQ0sB5d143uU+ci7aWtVTqIx
E5f9eB+uUdtKQYv/fsEa9H4nPfkLFx9isEhN5eHtO+qOTmJVt5TZhn3VLCaUHhh/WCa+iqUGnmEq
aH1vdulrwQF0cz3ftA8BJub5zjpjg4Lsj/mpxO8NmSUpZughEaLMasZq106w4wdFnsKUBh+iUCPG
+M3jERpxv1djWW3CZAm1S/ZpTiRJtm0AGy+hYyuqK9mc+R16kYM4pPRsu4RUSZVnATWvHznNMLHE
gEW4nSl+iuYKqWfHOqKIH0miKjZtteNQOX93bxEbNZ4NNKMrdDi2AEWlNd/M3iZMns0bH6EivwOS
bqM0pU29xpSHHvsaZUfj4H4TY8kcJ12v1eAUpZZ0Vh4Er1n2AYn/OwyXoXUMSagOtI1+bgC1wq2j
ePcqOpqvoUrO2Tf3nQ0qYAMQgVraetlMsclgIW1gfNPS75Ub1tid7l27BEQq6gjlkeFFNV+TWkU1
iErkvXJaCsN1RybTYCnwadISQhCoNo+s+dT6TrJumUIHAcAhzFeRIKfFzXvh2OxeVbAOwjBYogkm
e9e4hRgMRtbMomdmFOffLVb1gvRIpAhBDjTooSxxynj55t+PX9uQu6QDv7Yd3m6RMAXJn8/gQHd7
LBjj7kb98oten6xN7AVigj5rHR9BHDhpJXuFGVnd9YY4/B9T8Sn+tZ94t2T4v4zNdW6wYsfuX6VX
AE8r5qBM1rL+85aTFEb7eXdG8fAaRoLU8SXdJ2iJjzcuU3kSswuKNtZwTPY7V/fm2Tyeb3VlIdiH
e3/0PyM36LM7a6jMMeXHv+gCPiSyJxN7Jxd4OrFHA10o1Ho6JI/208Q1bf4I1LqyHg8OaBKzne6O
UwUPyzLbpozRNQtN73qBSprjae86WA20gcyxKkCuGoZ1KqB0hgUnv5k/ius6b61PSjQ9TE3vi08Y
z7CwpmBUHfcK5t0+VvUp5uW18LqjbwB9jO/iVlBXTnCQvVKYKbu1aF03FuY9YLWImeKU1URa65Lt
cvnuHwqt9g6PWrwG7zNwchrwkjuruqKGJRGdOHTMiPAKMuWOnst0WFoy0yowMye5EepYV07wACcO
10Oyuvi8serx4STs4M1OmzGfDSZWmyhGAnDISekJME2wpLJP7hMlz3k40NCU8whiQGPuuNQahW+A
+B89su06Dfxgkh4W0/Zd+Mc9iF9sDPWB1OWYbEabfKChJPcOmrq0m6EumZi9+544FQ+Gvuu5Sp0m
B6pR2oTygVOIqOhLdxZk1/HNRjkPUUJVX8Fz8YIBeLaizinuRlIn4XDNUWaLF9aedX2X7k9IGD5G
4dpJpU2ZsHZVaK/WziyhuaujbPfgpZciqkaHU5XQkqd01LIA7znypIADFpKdkDh5ak6QciVh6ZS8
0/KdwU0a6e5uEBFGUeEwnyO/C2BJbGRfAXntdprxlK30fNJsyBQt+1t6tFS2iZXew0aR7rwqB5Na
v9uXLpoq9u6myaslHIOHOmTF08JNccZfFcQQ2Kj7YML/Pz0qwzy8M8mJfy4lfV8tGEcw4/uCI4mU
kCTypk2kgl8ShmTPOMsOdg2VUoOZkPXzIuynGbG6/TAxP0Vx5j7xBc1X/LrcdpeanpgIGFiMsf6+
vHU7gIHCbQRYYi0ysGcBbUuqoIK+SWbm0O4IbGihvxJuHmtHNENCnsorN0F+xue1QCGGDGLoACXu
SnJWp1KCLgD0wWDBjqyx2RATHshecQ9XhfMd8vb5pU/YZuKOXVM8hI3oPfTSU3494Dq2f/qlSr+q
cvj7QIwcP+pUd9crylW8t1/ZhgiujJQIoyH8MBRv0kKnAICQvGAX2zJDvwoM/eP5+DwPKwbgjaHb
Hhms2NYVOOJ2Bi6yDTf9hcwNM0zRPj41cLXSNEy/NWNgLr9cD5eZxjLzuf7GYPcwoR+WfoKqyOFh
mngnuCnvIUx/KgoZ1PXG8RnuNkMZavRKARF6h++4Dd+o9aNzmwUxDbZI5c5Vi9fGmwO/z7xA1Trj
/nvNU9lKqXhu8dcaH622yZ/lFY38IXNMbbvxV8Yci8NYsCXhlfJ4JVngH2YZ4KJJ7V+kGLX27AMM
VFXf5m1okWzhepSXMtospuz/OQJVZN1bSieHqfYg84twXAam13YAwscVkxPauuOQpPSwinlFNXmK
NSLNaqKoRNvwVzgqlOBaMhPeMfEXrKN4ewz7sg6kDdLHqgHtkS+R/3gsVgR+4eTm+2+2q+kjvFkm
n9mJgTRqTdVUv2ow37/QWZC2nwG1PJAntg3H6JmEKoY7UysKYd3RD9HBElGmCvzdNCTIyYWnsdTq
uvIPJr5Ar4ispmcvQhtdM/sSIn2y/Dbi6BGJGu+gvkNziqtQmpoKdvZA0cDJfygL7651PgmKlSQm
ZTaOQE424G9CyiaQG+N3hn8Ivr/TDqg0iI4U5tESk8raAe9qoK6RLikc+Fl9iNkgSQhdAhzRdXum
XM+44cwYVYwXz/OyQz6Iz0pT53NPFJFgHVQnugaR6w2qZ3H54LRYvSdBTxBItErxebRvLKzNv+UZ
PamvINy/6NaEMp2Hu2/0xEGlginh64LyuIX2Wq/zFM3e8OPVNDu6HaaIHpTTi9ulphQaJVNj1cc3
J7wovgsuL715ToxvMRmkN6K8sdrAMYufN41yV6dCvNzn7/T+4lNFM70Dq1aV7rDen3LRzCQHULLF
9DunfrJnwtaj+VTTDtLV+ezic9CJEv++CRLm4h0Zi4F/h8kYWlfbfyky3MZBP8mJZJjae3YFNKZn
PL0xa/9rFGAOXZhGZo9zZXI2gunsGxjLklXhQeuD1rTKZPBTQeKLGd6yoGGRkHTt7gynp+DtzO6I
gkmwr8ruKTrwO7thr4OHcE8sbJSHqDmTOCU2f1CkOxAG6l58Vfki+BRFzO/hpm8SuwO5NWFuj7o5
1bup7fsHJ3kHp73OgowmbzKp5JrkfSVMyopq3+iIjjAOAg5VpVucHmRpZ7rg770vQ73RYplQ26DN
+JvIWeK2ECgnN++FefzUz/irHt1uFZ2q5bivctMdgmoF/RYSnqYzldztLmZVBE0GZozaJz5eE922
JEEUBvJfWhQGr4fyqaBQX0T96MWoJ0SN47zrECO9EfGs18EgINhb+19mDBtEFxVTcm8k04XO3UBi
8gMbSLKVV/KJVqy+0exdLV2K7yGzFT5gAW/DzlF1jP6oPNjC/yQ387fda3+ZqVmduKODRVQfxTe0
cvUMXIk2z3KPcFsCzD28pGZqbzTba61hTdrFRnwCxE8TdimEp+VZ6YGcmrGuqdQLpGObn9zEJH23
WfLtGg+YcUIPTq5ZaSkHt2svO5MMGC7F0pwTI2aOcm4O2nND1Gvy0pF/etzXmCODDAO1ikTCegt/
VmwQB5AEAlKwujO3dcLRAfExS8yyNyT2WplViYySp+qE6fZK5NVwo89s7M1ab5bA1KOWrffcwB5x
DxqU/GXed/j81nEYi9p+Tn1GrQ3xDYf3dWNd1sk/wvsbjSLH1ZH1hGYn+Qpa0CwfHabw1axrTJ+4
phCTBKe+gpXYv9zmDEZJntX/vo9Uc3/x1xenEDOt6THvZZe7vBlOHR23lYqls+Y9glCmwuk8UGuq
81XEgAWMqN2+PuisYO6NeK/7cx9y/xFgGzkIVrAC+Fuwctyf5hCmItugTMneE3S+tMAQelnrlkUN
ZdIn9vZvAaTxsDE0BuKfDwsvsosNoiATw03lzEBovvTTtB4799yd46VrAaYd81Rt8gJFLbehmjJw
XeA/XAm/hN6uvzPyk2A1lWCszFhBkMMCjRJSqPt/l6eWwqVbDedbTxq5MgqSW/v8NfiNioHdHZOj
tntrZRNv3zvclKbSWZVgpxUX+YeDN9fJrNWGpzG7mz8/d/SWTf1But4oIKzGSxH1bgMuQPrapaK3
HczX3x5GY0QnpRhUZZIsgEUZbf9vlNBmlFh+mFi68lSjQH86fFuT+UNADyDKkOESAr4RjIfTrBCb
93pka3ZCpcaRdsSRFwFhiYOaJPXt0M2bmxWIp43B2qBBBLmhpBJZv5pe2iFmKgqF94uMlhdYc6iC
X66vj5j/IZOf/7jRPE670S6VBBgrLADxb/HVZgOnvNiSEr25y41LyG2HGuvlfaEuR29UgR295RwO
O9MwutEw6ciHz6/Di+8zoKfetphz3jbgXpxENaCrJNQ3eeWfa10cevVQuJJRMOsKQJpMUs1OgfA1
/9dQOS15j7y88ahz3OZVuLagNUM/inCgLWisxiNlENhczjQZqvkNngPP20zRxxZGVeJtYQXAuQ8X
VceoBToqMsZaTOcdeUPCi5PWMxIVNotOpGZQW6iNK5Qc/ZjPRZ0qvCekIr11Ki/XHTJaWV6hUYus
7pSgJbFTDfGmt9yA6tlQr1D0wjfdFAQ2LWt48A/8FTHoOiy8uEEAJxAbbrzZc5BMwkSE3DVweB19
BMwvtKbQdwvRRNjGpynFn/9v7vRy9O4WlQFnFVTwGFjFvAFXYeEmoivN9UAMb7KgCNuLmx1CVuQA
+A0s/kml+HQAUUI1qh6zyzoj7joxkzIFGyODw5jHBOYKWHz+ny/pHTB9WE6mEWo0kMYbzzFv+Dt9
1RgUf/Ww8s7umfN242NHxLQ0WWUIOtjF1nRAD3l2SMPvImyjDa0Eqf7Y0kh8374p6CAYSCspBBPd
sY59dJD8eVo0lw9nC1L07Bk6g7PP8w13xOgNulSmVlCj1hTydU0FL8z2yWxADzfD7Q2as+Qx7GoO
rn4AXNLsdhm8NNPCc/kIiKGG5NjIxAAvb+0TO3yvRkncwa//2Ew3ENE7y4F8bUYiqMO8J8wJkXE+
qgY7NuaadoTIfeLxNtG02d46qJuaL49IITVCbljkU5VlFCqdiwOp5hyIJE0vMVmYyBmB9LvMCVV4
XxxNAm+bnMPJ8qlqtZfLvweKwJpjWDCsgchXkg9i1S08m0WA2iWiN1lOcY0S7nQi+Izeb1OA+Y5K
8Tvp6xQy3Ml01Y8QJr+eiHrp2EypBXTjd5P8kwm0cSY37TXgThOR8ftg46IPtXvC11YgriKv+2Pt
iXfE0kcZs4aWT+NvIaeV/YjDvjqidNOACaVbHGj9cXT3wk4ptf2estfVW971YXJPIgGbQWruSRZq
BO8rXIv9jcYcMrXqm3pGIjo8Sy9eQ+l0P6OSsCZona2QX/3i87Q31dSMBsTkBXF3b/33TZIYZm03
Uf/0+0Dk4xtdYOnAV9RmOLSJuuria3s47tVTL8wdNcA2Az2UTtm6DHsMh9wWnbBKW8licOHfX4cY
/qGSus9a2Bl0eMClwOG3Qv/spbYUB0TYOE9U6hlM1vgLs4HKuCsDBfvh8a2aF9+8vNFg5wbES9Of
Y9Q+75rear0N8p7f+UFKcZk2AUH2xEfC2Z0Emmg1/VX9SpPrWgrddBG9PJvnF0KtgFfwX2SOuHlm
1SX9IsouB+ddoMROQGUwMLdlHYlN/bCmfsWmIWbJqleQXJMQHjLR3faywdlpjHkE/kE9GT2zPpR1
Rhs+aHHtvxNCrm0sqsDlL+GTTSWZZzHUVZzzSsf3FSjGkyLJtcmtXrWbw4AcSrvVSWHRtW2ZNbIL
gUU2t9NbD5qxIHudxQg/EiOppyV/ZFbC55N1s+rxuIAFY1TCeEPMZN99Obf3DWmo1T5cO5lhl7on
EP6n1BKdiYBAxVBp3z3q6/jLOki1RFt2okIzlhRZLHAF4FWa43oToOfUq33ZIRkVLEomuacbh0Je
RPoQCETWwy+axVrij+GLulPzuoWOJ8jR+hADvddcCpFIVLaKn/2RcrGm+uB0xp3ujfyITAu+cgPt
Hfix2QkdSsuOvv+ygN7jS/qtgnsKdAlySBRgLh5Wzv2eHnhBZqDcjVutOwqErl2VHFFJ7O2rAEv0
6wMVqLqyEx6ve37u3qhM+xfKeQ0C6MPWlLFlxyLP/PArPA3tn+Ew5Mi31Q82/59yR74cHQNDLmsz
NuaTXooVH48245i777CwBwQcY1bZ6SwB3z282TC68VD2RIvSpGs6MGFcmYOgZRa2DYSvAwPScCfQ
J8OROGRIhh68KDG926mkUB2SRDs0HYZnwP8yanqRWXts7Fx5EMmhhhrQXxAm+wIWlJN2qko+1mgr
AGuUlqTDwfE/GLDo0nxXGMQ2Xv7Q6uKxbOCcoObmTDKSjBlRXLzY9kJISfYugI2fs5J7ub0pJpnd
eXnCVz8wE1U6jXDeLqJ35cRWdLyh6OZ9j2g2TZgiLY/wj5PXglB1ydV6MlXTs4Wz0JKMv5sryTjo
G05t0rdWixveHfcigyziIOknuQpAyjLKIIV1/AM9389sGLLN/ZhHn26mainWeabM4YdGVhIGy/CB
abrXJeQfFkB3kxsGT7LUKjDoY6PPqIf2c7kStuwkwBO/9BLd80ut5djNPdhAiXtUXBrNC1YD6U9B
lqNqdYLmN41xgHm7t2uVU04KpPuTj1f7TQzEoc1QlfPULWVmxnQjsx0XJ1zpm0xUlR09ezYtdR21
GFfttU6G2IgoOLiBmDbIN3RwDhBbYOzTQK4fp7vcAJDfKwJ2ZIB1mcxwky1ZcgFA+NCrYtO7pO7W
v9o8tv+K+udKr8/HLXZxeyeEMuUaYVAkz6dpvPhCp1zjSzuDoleVh4QzadIxoIZH8prEjI3TWvIE
HgyzYTmAZgAJhKePuANl7k06Rfv8iaT5nqvKeCBpJO7WkHDGSveFuoPo1sbZY/5pz+TiCFxxuXpS
sDYHZoGIRrHM1n7Y4d8JQ8epQ5keCKmmimKMPoas7EbAIxExwqhKYll7fhbpXbLWxgGHqweS7lkz
BGW8oX8c+a8zyd6HMmQZE0cBqXwlE6GnYGdL7bcoam7dPvnJYoSmG8JflOUQR110QFYyPcGEMGU9
jdg/3yzhFIE1lCM/QtzlgeIApbd+VzzbvgQx0+4aQx1YUkcz0ohw0JDnk7KOMRc0qJmUCyu99+OS
p91irHhp7hFJq+k2tk/LsFODNtdLNH3u09YfHtx3V7orafpqMK9abfsVJ3s2uPqINON2jUARPDEa
It1JagFtA1b86ix+vrVCCBYtQ4big13cUcsaRh9cRbF5nQahxBe2TUaNPPn7vFP6Bbasdllt3dYl
7BlWgFSE5kI73xixeItKlx0vDL6XNszBeDCrFzSpq/RdrJCyawneT7L4KjlrDbGMGbc+gXrL2ipq
cX9KuXVEzLDEVDzPIhAMDbeX9qiY+Yyd3rz3EAjOT2IyDRcg+AYY8wqhBVeqpmMKWIhCFv6//Yz4
FmXnhhYJu2Q2BUzXDzMqLzkiL0ZW0aAp0TfD3rtyESfhqk3uMgr/+e6P7vbUdk39jdy0QWm7uIFm
YNcCz0zr0wLsQvDGh3Nb2MMgCXUUK6uDW6rhXNHYzDx8m54oOca4p9HH9zqbBvnzMNaOzVLVs2UQ
ivNmoVKtViGVENBZ2ZIWJIE0pACvcBx1qnxRGMJQfsRLMFPbYGylKYtycdJElTuCk720QEWrVAYz
yy0bBbQZtAWjSQq40K1h6m7AC+4pqxvVeQo4y4nBHqOSwRT7hMakYtREyWIXNUKGl7aZBqSxOwS9
Ba60GgGYIOVUh/zOYcUtL4f2j/k8hMsIklZLI6TCrXhXSQS6E5Cnf9IE3PD1awWtS9dO88mDUuca
Jug6TCtXCwcPINNpjB5dYKkRUZ57nrmZLUx4SBpc3zs6ocphP2be3kQvla9wjGHtsvoG1nspqjOI
0JlucuYh29AM39mMDwMx4PRohTPtD2h87wSt4NJajWxIyYzyZ3vmsH2UmMaoetGstpLM7KUOEu5r
0vsgq8kstHFDHx8CRIJCPu8087bGEPY/BAd81ri9O8GUqKIjeodEG0gX9YXgu/JHAFYCOZd/fmPs
snsWTnooyAEnbiRY5DYnpQ9c553JInY8fXawMh9GmZa2jos/UhCxm6G/+Vfo/8dr6nExPRRuW23d
cwiiaGPJLEU7ay6sPuVaCfEyRF6GxexcVqFolpJvsa4vvOtdw75KGcTfirQgdl5kztzDkM4Sov0k
C4j3sxx3m5rnCp70WJM+lraVN+XC8zPu+uvVLirVPzWBesvoMFOY0cmJNxR9zpci8O902B6iV64U
tvUX1kzDLNPCURJCKYnbtebGxbVz/jgM3M+23GeBHrkxIKcgSR3JM+QLZFr/4YuvNg5s/fDObTwB
8EGMymJjHa+mO3szmNZfXW5tz06SE362H55iFjn1lGV/tMCG+8OL1biAD7JwjMiWPHYcZdPfnkRD
+qrBPU0HYDpmv6Pt35Lh7TxPSeeOIRqLBxhe/+W6BlWbkpSaw6X7ZaMGRnLGhYmxremmkwOwIwH2
uRhoi+zbe7J9653FXr7ZBC//tGV7RMt6whgN454K8UB0iB9TLZNnN7+43cAkchZNgAs8QUPbd1vJ
S6F/wL9ALtFJCcgewAJVt92ofMdTUTnfPLlzfL3GED51xi153UR9tc5ZpVJLEcB0NGZJjpr1ZbQy
lX7AmaGg9HHdPpMfzCingkgmL7CdWzWJ0DEOaNpcCUV9Re4J8/n93v7IhyxbdAXEyM4YkG5p3LVg
j6RffBJkg6uTdj4s3sM7m91dEQ1rmXYV95Qxwk0trWhGs+uhfK9aSA8W9Fz/F3EEmhCLKhQcNUqt
Q9x+OOjH01UxLwoIiZ4v0GhxUWCnR+2ORVg2gHhTxc3XsP31I+tVayUMP0T2IFzjHB0qR7naIYld
7OW8xst602V7c798847fR9qImU4OIO7J132RGLY0g5+CGmAJmQY1xqmx+/tkQpvRWffoeqk4/IMQ
zlSmUm4eTUPTzdDo3EW+Pa+hyoFzrUKkr6eQOI37AeQDmOVAcqhoYOR94ae/jxZ41oKkaO47PRjf
K42WH0XeW0J2QJWC/9hyj1UFgy1fi675xcoL+PvWrcc+m6TAa8V9+YorW1ZcNLUbBOPbcbacaM02
2DQGgFD5CbjaYUUApY3im2HAtXJa+rMSxqnLyVpdGY6+UGwp6XVyR91K8JmYdWtpR07IRHDJBD3D
Q3HElkqYHLallBbxy6H3iRwqSBh51Uuw53R82666xG0pG1Xg8x6dliJt1QShet+g+YbVz4OSX6CV
Qz62jCveZhPXnNx31Z0EI0TgRprqUezDzhTNuOZQcKx9LbCBcalM3Mgh6hkYfkvnlN4xLIF8sFEd
+wqh8zEyPaEctjWeibxbHZiB76vP4CxI4/4Nc+we3MyywE1iufitfxzy7CaKZVzXqeykVTxZCZAB
kbs3kKcsxzlRDCoqq2kVkF56mP4kRw6XzEnNz0L3DH/YYOOFRP+yRESIP/TCvYLHrczjUbYxwKQ6
OCJ+1z4YJ175/+vD/ydcQTxg/6qotKVma5qiePy3Do0c/O6ceDCnz798iSY4954weJI03sS0CREt
FwOGA6+aCRoO/mD7MTWd4Fex6/yrzirSLgbWy1+1c5zU0eu5QR6Dum4LdW+dT0HxVXteO6IDvl1R
CaTw34gV5KsFyl7SQ4HZobI4w1XbHqJtX2Fm/0iNcDoWkBDAohcslFwDchcWKTAkfn9VlUyQyhFA
stGZ+PercKFRJqerXIIaiuvkP2KD0JlsSijlk7MOIYfAr81/uJcTo5TBKjLZ6y6EU6OZ/b7pWoKu
xu99OaixEtS3T4VaccwmU0lt0HAxI0HVJnAnPKD1aYgeY2hS8Pb3Yf/IGBQAMSxYhSiBcLShDvgA
8BwXmYeYP5eCd6+EXQ/GjUKnc8bF/eFhcFhVZw9Fkfp9/8UpKU2RasGpE0/11DL1YS3JD/P48NgZ
aj/vNJ5v7Ba4x8SoEU8TFCd+vBcOf/kjLN9nZXUfwBXfv1ENsGPgOuGiDz79Bb8lVr0QcTxJqz2s
KeNmzRJIkXIXSlWwR2uAXLuPV9aZzRg75wzAhYaldUFpM5YEdS+pn52TpcCvrZn9v51tmxB8OdjE
3RdOwzlLHcqXB13v3yfsGqukfzkMf4bqqGylP0W1qDk/kAJFPg/Emy7iHa9QztLF+Rukx6Jby7Fp
9BntEpREUhYKeFXINNnjxklCyrx//G2+tFe5FZMwXi2htSKESWdd5sRazfAaWWf5cCUt3593DUvC
7Gdm/S99ewZqoZdQyKYjoNgsDvBGvfIw3ziCbp1xmiq82dcCd66Uhn0VMpBaRyOQYh3UpzfJLRs4
VOVvgAZ9fAPIHKvaBbFR+X79GHsXJqC2gXe6XaclMMn2mRKUfdAvqA2RhGnu41K/VhH6N+gT1kSE
qxsViGzWLkQmOAEp5vwHd3WVhJUoh4Ita5E1EFXSfzSBuTaYGY012qLoL42lC/frgaiKtUpzuFOt
q2XJb6BT+BBpI07KoD3kLEctxGzzoW0EfHLvMVktFpfeNXX+OeANm0SmLlDfERkqvBH/B5DUWac1
QXmqMFO1Mevx+nMXUml74dzIVaGH3c6Ov+Jslv7dHg1+2PvKZ7Pu5Fg1f5jxKCL3iOWdyOvlouzt
3FSmdKHLgZlnd1PmkZ5eKCS+fYCzFL6WS2C9FSIsIMnzlqTquvSwjczsLV3xZaWHcRSiqoZ65fR7
GYwZd83OoGiaRD6W9O7yJjzBHhFNjmc0shiGceA/j4QyqeZ7RM02vGt5vq40qM7U32HNMxtu9lay
vJhbMtrNzm8hgBwWoFMfvECtpXvpBVy8sJfoEGys4rTHpmNhDzuiVY3qn8g0R9jU8I+5XFapZoHr
crJcL62YJ/4dFqYbET8+JXPMbmbmwTE7WqhFAXZmwwlvua4Rk2mc3+zu/T24vUDkF7d1eJstdHuz
LEB+SNeUW7dv/07+/kp/ysB9Em1GQPFeqQKNAtZSoDRChIiIUixWIOoWaZN2g6mcMCFG3r54mRJh
1heuViM+Bt+dGl88hXsaqmMTg9PXWhOuGMuyKudpDvuvNphlCYWxjY9dZOhuPezEzkHjMcUNbDex
C74f64OQRgFsGoh4rCNNuj3cbxkJho9rptIiOrHjKrtRsdqZD3HTaR8XnzSyTnYx1ayjsLjzscZa
dtwE2xmDc+nDalbaY+ezrlVWOQR59NK3c9xI+LOSfR4GK6HML4Bt+zKBSG/lYh7P/eZctGnwhG8v
tq5WyDrbViO9Wl+Fr8hIVPFU12+XDbXEdQOenQ+tJxnPcwYHA/jEl9nREqvibGeo3m6QG1tBXnz/
h5uhCBvMZQidtdqlKpWpKXXv7NnGQyWAtXECgO/zHsBJNrG2YZx4ufG39ygBpeU1LUKfr/PY6sTp
uq7ezAkfTx/6lqcUA//AuEiHshHsxkHJjTqnTt7OnqfGDSbCQdBDDhjv2YH8bQMIJ1NH8UUxWXko
6jzB02CjlAmtaxwGDlDzTqaD8javuQqi3+ENXHT0tgA2hqjdD47+ERKC4yCN/Wy4nx1rFN9HoV/h
rUPU4nrz7+kRJDu8sSyLd10XK/Vv7sCEh1z9TKWNPnLi7xZi+Y57wxnMQ2DrTU1Zx6Cou44L27Ji
lEy+M02Sh+JYJOoL1GWQEdqyBDQCpi5tHLkPLXUb2SnNf6qYbTOWmrw1fdaz/xQS4ye2/zQec+5P
NyOqftljxGJDXaxplRaGznrEV1GRljqRFjqYG2gJ+SP6ID21rp4UJVJ7O/eQ0zspuLD/srQVMat+
pRHp6kC/QhwUe96yiDKq+ySOnlgbcsoOivp+QRT9jiq3hW7zLXy0sAcjur0ewNqueIbiKMbqO/6M
urdF7sHFyhkd/OzcPU5p33qNSfBjwBcrnwH+Db041h7gFDZJhpyrgqlatn1qS9BQtol97/EhHCTM
wPn/I9nTI/uLGj+PTmRYkgN9KbpCBG7QGwEfcwD2P1EJMwIpY4sLri8Lhm0cXLJR9ij4AYidAx4w
BXiX4pqczqPAGL0jcCZRaIOpt7Q6TGM/4GgN8glbXAmM9wqOzKiW/Q7TGNJ4jmoN6fRV37232M5l
aE1Yu+ugogIG3zvQnZ3eJBFK/sO1EbOzS0h4Dpy70ESPnUBbFxhTVPk7Zb2RC9zWJUQhpb0LUgXj
Btjsf3h46aQaUU9D0o5CfjFnfo5ywlTXyveeNlD8UbE6MVuDh094klmBZPNNAUzoyQhYBQa/Q8rH
W1Qdgn0mlbeWNaB/80Ecz9Rxmr9pHrEJmnRGadXVfK1ElwtqeJLQMCKVFwnITHD2vgc/haptJxRP
XsZ9M3nk1ETLJpQqubVBHQ2997k9Uo+RxrlGzvCNLdeNyM1kS8IMAiM9ln8HLUIAASK8NaY2muMn
MGBSgkM0P2Dcsp+LSZYQqUeMf0/1HJgbZzlJO5Vbv9O+H5if7ghn21oFY1M3h/GeU7v0cS0+Nm3O
C7WeCg38/FAece4taZmOEPH/p0sLZMXpG0GMC0v5UkcRUBnQ/apuPe0fxymCkgiBJ9QWXQKulsPR
VitWcpUuGw1MvJSGI+LflYnlDk2lpLnWtSAACOXPiexO1K04dBW2YE390K0hQQkshiLOcZrrL4AM
1vB0Qraopc6AUDKCl8yCUUojAfoFPHbnGmIGlP1lCq9s3E7YGoVUN7P0NMAZhTPjBxinHs04kYLD
JjbdoTWSbLXRipOsaBFyW+7LJ4n0VKz9T6xSbfxmErUet7ioXGIIPtB9hx3eSfzgTttIoYVQnmfp
wd9IjGT3AAqED04A4a31j3JeG4aYA4m61HqCf+OlUcDV4NL1WccUNsay1NIRe/HIc/F75dhfqXEp
XAAJxnCtJIm3yXwvWrUIkIeTbecW75sjqJwkxmhZ7Ovp4x3DHyAW/JaxATGqhkT27sy+cBCHycYU
xC0rTHk7yX//ZvMFBNtYRPgqudjuMQldQL9I7qNYk4XLPO/w9Jun9zRd+yvHQWCNDIFHisFNDbfa
DLCphhflZBGghXXuZbGj0j5Re5qPX1e+3Anfpbk9VXLRiKFVShIgiAPoeV6yk5b2/3cGUBvmXFdv
1YUtVh5sv4deHgjHjDgOif6P0SAaFhL3C7Liq1+F1auJetSqH2KzKzQGHyv3vohrKcrxsoUaj3/k
QNeV2/sHid5G7t6ymaw1KSYVmeCnaXGatChkTCbN2CoCqgvYRv6Cpd50mCOcFqL880yG4Tgj/kQI
lhXJBbqUrnO6pIBorclqaXPJqCP1NQxjkL2cGeHKEyXmCg1cngopTgZ0hzvMlYcyIMNFch5b3zgk
pPxBEN49sDt2pqKWkksQQRxOL+DcUIfLJiPESCjlUIUyyiUwJQVg4sCnM6RXH1ZE0YwoHBtHcQrK
7fkg5kjV6yFG4EfkQ50Q2Vz3SVxdLipcl9Mw815eMQttRiyCW70dvyU1pZNh6ZXASQXhWDalEUVe
OKlMf67naselNaff/NnNbac4tm6puVIVT5wuCmF7Uy1wtB6Pu6MH+DCJjqWeJJHENdK/BeMbpbGD
PPXINlkNJ4cw9vmTUrPLZdyQSesNa4DGPr6OYX0KXRlDsthYQ4tjUtx4P78fsZ3FIscCjJP5jcKv
r4g6Q0UJeWpA4e1AM29LvsSbXbMunjhx7FdOOM08v+kYZOrZJ5sLXwWxAM+1Qx4XKFCXElUZQDG6
EOcIZwLeEhWWYZIsvKWKA2SUx0p0S9jQ/RYd+QYQAMkPWLWc763gOe1Z+t2b0roEwr0QacYJK1AD
1iR0v+aO2AURHogwcgEqnRQeVWUZiCwyX4HvYTkNRjvlO5c2lGAudLpc3UesZvOCR2rPnUBL0ugR
igpSnBQ1oXBhMpcH45s6xzRYDaQSWJ99H2bERbeYjUwN6JizE6qKsIW4oxkKcqjN0hzir8QQz/Kt
exZ81nyCnFmwYa09BIwEb3i5FbQlsysvQyOKVxS3UsSDsdf97wKj2hpmg9C1DR2jmZwm82qDo93c
bA+iKJNcmh3fgW4kDE8CQQG4m3SfKCBfra8/iSft0EF78g5MpXAT0Cop1vH71/mfVVbAovYGf0gP
BtqNzor8ZcXQAN98B3YSuHB6f3J/P5Gw2WlfT8GqFhVUdLRHFY7AvWcAEPlZ+f/DNUo6fLcMDd7z
ehdITq48ir9CJtxY40W174UB1rp8NY/je7rfzMMolwhfKPOkX32c0fTdnYqjaj00M1kyQXsK7X88
5aqViSmkOcZ+ZMjUZSg/aGeZ+yP3MWJgZY2abP6sM1lx/pD9U7SZmV9Rg6ERtxkRRep5QtcQ2Z6a
wf3XXY5FJqsFM4SFNKfmV1TaUqHcle1lj2tj7E+4mFJAFNxPm3aHzaCwZcr0eLltwqVGke6JIihE
sQTPac0+trbRORwYqrTAeVlTkFXdXGHpmMorJiPaZ1W6cJZZsZi1EctixRhEPU+Q/K/fqyPGgdWh
EDnQIRbo8w73LdkN4sGv8ISbOf3QY4A7vun2/vk1YtD8BewLnuEqVh2DZNrXqBQbvkNZLAQYOGjs
h+WHtuVh/SqNOIqBsAxJDkeBSjNcmhWgPqpk+CZ7WGtun1JedLl+LrGZPoLRegxlH5UTrzUlgP3v
qB+3Q746kujL1CUciQdEypoqKBlDm/0TIvc0U9kpVKr28kg9zKVim8XdLkVaYg2fP6OWCPmEU9mJ
1q+d5L5wr0qZYR7sHl3JR4mBG7HaPrzVpVPo0dlqqTQBsz/oOLR7KCZOghU6HM77EUxsbN+Isiwj
sVU+1Cks014PX1Nldg9obENPAKhhckuSufmOzJhqG8CEd3L0Qz+h86uGiMPcXCeCjF6CyjznVgYS
KZNBs/uo5qdUjcGRzucSChbfB8j34UkRmrfCv/nCQH/XvvnPlhFdernaZo6OjTeY42qc/f+Ag6hg
5Ld5BslJSanFzqiBMWAJhZ3IDfwpFgLldxCs3jq9Tjhm/Rtb9AfMGu9BP4OZT+Y8UKJUV76nh6nr
9TF8gcpXgGalmGI93BvntcPZqnZ1nOrVdO6xAjuKv7wSlKIGcsAqFu1gNA6blkwT4gpNjRDiNIXE
w9obRSDIb/8RvvBYWjizEe9pUsY7w+NUs/qPo8Uq71L+7nqFIRo0tnEln8CkRowFSOIILUkrclcP
uVxmeda1g4Zihkk50qGMH8Hxlupm1YORknm+uh9Q4nPa16la1G+uvbtiwpatdV8gJiw7ehCPJzq3
41OM9OJWBwqUl/2EY0nZHqpwGNzxOke2NJqBuyUrsUyOw/i32mj9g0eB+T5D/Pfnqj+yQpXYLeRZ
iue1tcUCiic8JBwNtbh3FC9/pFxv0ohhvVT+fLQFD6a5ODx7hwkTXxtCyHQ1LasD1IdMzNJ2mEGt
IT4IuYyJloXBZQGbfXWhqiNVSa3JO0d1aCHtbiNSoqkj+2nYegD6v4HYzXe5w+X2LmTgwU1jpduw
IRkRQZm2ly3TV1i78iq5uV91hMXtG5tjgtdgNM39QztIbeYR/rEpxRNQVlgr+00l4lC4VlRqTvet
8esxSfVRwf5qYmWiHPnl9oH4iNwvtnlChNEgPpDMEpPsYI6xeDf2YwknKxcTFtnz5BzcendyHbiq
//p9omxFsnwKtJxgVodZS3tq3Q6f9GYVRlo2dOhU/zxrgfDbeM8zbddmXGmkTBUNx/o248aywLi7
C0Bf7HfBHkwpxUK8KSw+h9Am7LLb0Tr5/qHO6p8KmMkpIBYrALIgc/bWVJ0xgZbMqMn2EgkehTAc
Gh1dWT4baIYqDgGtqk6m6HMiZvEiIz48Iwn8ciNZcr6tB+l6NttE8XTbc1faHgSAjp9FYHTZgVcE
/jzJbRnqy9k5ohIu0t7qtDfP1r7fv1oasRbBh5zLm7C9JsuBNETC4wQkaTFnXHRAf5P8WORpgJfj
3d+CnedAUGv+TCy1BCm8O2H3Bg7gSIV90OhCXw8Dz80yOODNB9X848VOsF4nw48YrQNQCWCKAsB/
p5c7KZtzRmaztVnAgMTPp63tyTVMFxPgcF6vtEBOfO+Y8/vswBJITDjwK9SFI/ruZkhm8rLUBs1G
kHHlL+6SBFrr5VDrp0XwPTZoOcgVn3qTC6Gv+yfy66Zy0xNh+0usMyNMFvEIq0zXc8DQu1IWh0lq
JR9J/ngMUlx9rxNgXYWXhOHYbcJskLk4dZj70wwfWKk4+/5HhYaIjOFzpKvsUj61a3OTv6yJXJzu
oRNGC0VZm+yJFCYDNa+BqusXSGWOzwzwEN8EjPt+HaDf1br8AiA7Ycaj67hNMM2skhccVw1LoLK4
QTXE7j5b8GUrXRQt+Q6DmFwepbQ5BdUIA3nItpH/ZTEQZ/5nNdPHFChwCiULuocSSnWfr9FcBeE/
s4hUHy2jNsy4on4L2UYBdKdZuFx3G23aX7VhSKu9wiV0fH0xN/jKHeicGBe5zs1DGli+teSjD5B7
l48cGpl66fdaJimz+uRCPj3jABBr3wGgQ/cGJEW7udqwkKwk25yVQQH8mUCDXQLMSdhSU0xaTu5M
ENCbyJ8vePALWBN4+q+YM+yytc0w9mea/hG0AUk6jALF8Ng2l8bEOUWVbhkN14/2zV25+iiX2GrQ
CPA/PffWc0J9P+H+jeV9msbYAjT9vSQ4lTCQCSgyGdCj22Z73crv8hEpxAVBhT7RRCwXvuC9TwEU
GUuDTZhf66GKhb5r88VxppIWcImbIB4e+IzDHu8dOwEAfHtzXp8C+hGPGEIf4qzbuABigsvV1WIT
aiAXtBNyrTGhTo1QZmEBPR87K+UIeBk2xp6ja9zMIBkdd8Xg+kulEgVDH0Jhzp94npLGjtzifnVF
zxzwhUSWyrp2j9sNXkNxJZ6a37Lyai6KV/I7hHIjfII5+5K8i/b3V8A0k8WcLGjWEQrqjLpfirvz
48TCbvFKM0JiFFqvH88gtDwr+1pzkp2LMn+kxy/6+uHvmchioPom3UEuZqI6/oGwGI56zz18nyeh
7gkF6F7W4hod3gzlXigoaJm1RoPT6PUN8xylheEvX3/e0gnKtUgZqrwuXe561wrG/YZimca4+goE
FzMq60vXcPONfbNNBVJe1ThhHcT8250wr+WxORGR9p+/2a/gqql8jzkjHcuRk21LPgaV5jESMc77
Y47fFhn5VWMq7+KmyqIGsrobArekArMDTQP5L8FH6Dcuf0ZaWUv05aJNbyHBtqqKOjOv+7ZY7LAj
CkA+qb4PPyNt/QfEtUYv9dEq0vPLGAh5uFtGHG6vBPh//FViFjlKiZ4w3tfwpbhjtnwmCr8J17qO
dcXacc4Cp3jtDmuxEF0ApY3VDvL6SkcyXvbxwVC7o368vmTXh81BvvoNwJjgBnw+Pb2Dt8u/twhK
J7gX+Bil+ppGe1W7HxwbFcPdxLiza7jyG8BLofu5KCSVzdVGLxRKrQ2yTMdAgtK3McIyInVo4p5b
XpbY3ClxreScdU0/knfESzfN9Hs+oPg75jqrRoEFDQvRu6ILmYd1BMwP2OsbiHJc/kwA7yGY3qJe
eXghdmlMz/f3FmBv3ihsPonbUXQ14Am1afws8zua2sTIXyaM5/+tV7ug/YOPFq9VIk6wuLLVFN7Y
ymTQchg2yg/EYLyQU9z47bHUSxxNJfaZq9PbEFmibS+AYsuZ620+X+yyrHXie1dFigwK9kklwRqO
wXZz8Gr+hNvzNsehuOd+yPfnHcD0nOY9KIdbTlT8gRizZ+YkCTDgovj8IMnJfsJ7YoRIhD6P74Dv
vmVd4Rm4Uo4REOOFa0zx4Cl1H9zJf0Medk26+rH1zq2+eRVFnLKRtYz3JldTexgm37aZXtF5XJy1
qNwXf0GbCRaCscn022xg/EstToKWUSdGh/NTWNffKbtIguyUFtnzO7M6WipJCp37j9qcqTFovHEG
JxNoXluiWI9fkFeziH9pfi0aishA1KM/8k77fcRZgwGYVHZ7hpRmLrKbyA56Wx07gUOHERISCzLc
/1OpiqJxzGCHM6CCWvyhSmtsrkJ3AUyIM8L9dGBmjeH/y4Zp9qSmgciqbt6p4Y+2YIc+2rIq96SY
ho5GtQQMScOwjekozUQbG4wYBLCD7zirJopw9tvV/bVOFwsidjev0laLafn7gf9Zgh0r6OgfjwOb
vA0YIb94xJ0w1KUug0lqYpRaKctHiJnXsQGq2tsEQrLsEtIgXI5Mmcg34iWN9V7Z5WI9b2Ed5LcK
gYIoelscNO1JOMd5hT87dFG/j15S4pRiZRVyqwGqaYM/E+AwiV8tAAkpaoTJUom8l0gGJbXj996H
THkVbV6+mRzJ1tW5QhrkV8Qtf8tXYBEgmjMcBNesqf8VsrzStkaDCWDxxSN21pN94q9iTtWazYAT
YaAynEVV1R6YMS16HPOOu2veaL4MwdSQY4DcvQKz/FBGGrgJW2A5MRf826iwLphULnr1VWogAB5v
KzHebr31LNFo0Y/j8g7rk4NKdAAVU/dSVS9/yXoui9Ybug0ibJybrObNvFnSJKhDUV+7lECS9Qyv
eOdf44RiG6AB8Pmls7ar57Apwv9f6JQxsHGOA0+aFYAav5zp9C3d01mactclHq3p5EowBflwpEWU
qOwYoUw5QAkH9bOrfPUVNQLpbydc+VLhOWen+zlruvGNtc4ofL/iYtMjpv07gNAPZVoCUEJs6mlM
FwomHWo3qBzkpwBg2sK34B26SkwHV2C6efEp6Wj9yv8go4Fa9kUbd3wJRdFeSHxhffSbx8zOi0WO
9UjlC//VYhcomOmvNtTzHjqjxbLyrmS08j3DbpkAtRZYegTwx9r7b3lzonAQ47jLp0CTP2ReNFTF
J9Aln1jfCe3fxER9BvQ//e0JOdSgC+Y8lPXLBylobQuTS4ZOZD9AlO9XMazCongnVgj5PkmUCezV
UKhIEmZ0Huy4QZfn6M6+J8t0SF2D48xFzl8J5xu++O5KFcuLQ8XIyWEHVz6FN06RHtul7lC9YNxC
Ysw2jhjAPwRDpmbc5hkYKqEriGWIYm4CiPXMuXCVXZT54buTNxkeFUg4bqboV2+uVwZKVcAHr/sy
flVAGU7GanAzgoTdrjKtGvD/0miQpbpGIgveFcnL5v893u2jsmMiVerO7mwAS55/Q1svZ1oMiXkv
vpsICrJBAmfeOFfzFJbUzOTgjfchrEGga5NvtWz/5sGVTKMQ89f5V7AKnU51cW/hy0NhwZ2ygje0
peq82S+mXbIMS4HlBkeyiu5mcjB6CuJU+CXjmkgLxhsnCcwgivlLEpuX8QGlubU7+fun1gMQzHt9
UaVirgzyLTezJoRDudf6x71khDlTIQOVoYlUAcWROtNWIe6+2KNXNI9iTdRu+aMhU57scexbLcHG
xOdt7AjMEBvHCvPeZgdzT5LlXSFQE2J2sXBkFEWF8unMRtI7ITIVNz0LMrdlqoFwBwy/quNapvwU
hmaq3AFUoqNG8qmsIPJAMtGY+RKBR1z0luLgGkxFPttFTLimXmfegs8d00D52nbokBAf2NxzyShs
Pob9MIzfXsDJ0FSXIGP9VJHn/Emk5vh67WVgoDzEdmcUb6W5paO9WUSXSxdpDpCyLWRPaZJ5bydn
9YWjpgjF7TZ2gT+ZdWragobNZK6N/8KFM6SnDMbfbAxMYAkn5dflW5waOrHRyHGJ6heaGUTKUiCZ
+oIOuF4ZjyK7FIIU44VKhCFFhDqcP1JOofyx9XCwoXeYaNUTf1teL5istLt6Z/jM4fzvg7bj8Sq/
t7LJfNS4nv5U87JDJET/4wgvHgUMeRZDSgIQM9EZ1IBKh9K3hB6x5Zv7Xfa7GzZa7GgHVT4CPDkU
AkKkb6HbTC2G+A97RJUkNvd0JPxP9D1CKokSayJu3LbdxD+04kAoBYxifxe5UTEdrK1HjQsOi889
dXRo9I4OLnC3Vawu8/gCuNS0nkFpyru6dHeoBKH0Bkge1uJOCysB7hkxo3gj7gzytbH72394LPNN
3rMOj6cT1Fa2g8Y/nsQpQ7h/T3aiSMSOCGN9g9MIQxeBrivsziyCrXeP2YQOtmao+LlmJAgA8uBz
tovUQ4umhR+yF53gWVmYzsFYLDg1n4L4INMEI1r7wJY2hb6lprZdiSV4LiTX3e47exHnB+nS/1WY
TuDAtZe1JTDeuqwrdEGo10iLBxYKY+6dHLhv1/IGXp90wseUwUKREK1LyEtTbOW88VdJwVMd3rp4
ZAb3lTPK38Jb78hls/Ml7OYNSgKm6W9QGApdvk53REM7Mm/0+gDoIkV1OA7P12kWG0K31wYnrN19
ls6QKB1oilp5vkCFhOniMwnjGRZTq16jKULShV9vHq3onDMls2z0xq7H/CyM9l/7ZP2Lt0HCKUO8
da3sGm+iO6ZYADoNwOXoHHcKsdIQzshJBh+tb9r6M3NL3GDRTVMUhtk0g7biHIz6X+Dlb54csxFl
A2VSE0rgFgsaG0cA1YkUAFm4M4F7tbBxNXpGG9OF4zGnLwB8rYTUU2TCFmawDP1KSJ7K9JOXW7JV
tby+VqsO1lhQAhOLm/pksMefW6CLPVs2Hh6c3ce37azdTOrK0n0tf+WZjwnnMnH3WK/dzzL+KE8u
VKX+RWkfPKc0K7Ex7HS2l+NRXaDuYuqVGC790NsRVBRXvNHtO2vABTdSdRsVCtXMwTuemm4+PQK9
ZppWQErLVe66HkuJYJcV3Ot8jr5Izf9JCI2YuGT0FDn43tUadCxk102OzzrN2Ti4hb7hzrE8KxWQ
c+9ZfpB/JZkd2Z615dgeSxTI/QY6yo/g8Dg79aW4vgASy5jiAa9q9PUnAxuqxBAXNq0bvB3fjVvW
yEOAXTCGqhTk35xAh2+C8gdT77S1q5rkFrGUfPzFFFd+GSjLylt2zHPBzORPOzJglfjHIE9l2vpb
fVhAcpnnWIp32fF7RaPLYWlBMri6KN3eDW9XaKxRhMVANGg4DM4sPjXQCW1cYkmBlHXZ+O2yyA/c
42SAZRt+ss7mO69yJHEsx3yknY5W+2loR+//GRoxaBecGhKzaVtKxno+T5d+DaKGhXSRZ9DOn+Nq
SktU7BBOXED+IcfCPrPnqrfss9FDiT1RunErErbJuFvhPpB2StaqoM7kBjTCJvrBRAZrFSNIKT2P
2VBEqKRBHu7hZxj3p1+feLT0IZSTuu7qddFx4M2NvurGI8AzshQyczw8SydbQzHqQ2nkBB29qwFU
otAlA2WBVPtJ+6ctFAgrwkVrEdBm5XoOyLHaw88X64ZSzcqK24CN+NrEbN7pfIK88+wgHm8sRySF
sdjJb8gQR6PCONj6UtDu2O9kT0rT69zSu2+8svg/MTHDStEdJShywBkxiR2KNBBSscaFnOWXfCnu
9+qjx21QPnQrq8dH071t8f4vOkA4ae40A9vJCz6rLoy5ChEYzAFI6iux25/P/ZNgUjlFNR2UlU43
iSAH2/wG89g8JNDFoBLflkC35UWZN0T8RUFoivBJlVUrIQzewV41X4TgFMnTL4xrdAJCGJIeNmv+
E8KAX5H1VyC5SuInji1ECth4qSW1nfaOlIIA2ON+/4WPNg8Xlu3buxUV++MW+oA6qpdUA4QB+suu
i/fwDDbk+rwIWBw+9jJXQAWPx3spxhHhf/6RVNZQjVWXaZjB2FTgEhsutmeChizvHuaj0TPxpgvZ
1C7Agm6UQDGCqCESRQPKhoanUvWLbPBOyt+kvJihgu2b+WV/v5VjzyqmOrlYNFVnwl8p3MDO++Rq
fOMwuZit33YzawiA395TH1v13ybNECQe3nB+jS+vtlPCmOoiJRXDv2SD5vYps/8vLSElEluBrqvV
kHXHuk34a76Iv+HARVhVG/mFu45CsYHELFHRLrnMvntLpMMX8yjlKYqk5f8Rr/xO9qoDZxGPNk7X
zegSyGrS7TqxJU0VbqsAh+FwdZnpVUNIaNQcyd854BFX1vdXu+odCV4eiY/BurpMYQ55Aqys/G38
XtgAbbcM3Y+NDCThSK03nKLxo3GDbdrzuGUaGow5wFEXsWL1gq7M4PIrUYDR2OP6PuCXzgOYw6rr
17w3vv9AXPiEP29l+6GgpHNfRnNjj6E5+a0OGkaaW8kK3gxyBSq07WH9SVjoaJJpphnb/XtTpItf
rTicWcnByCLQ6yps2G8TXHu267brpL8sxXsJE0LzR9mYZi7eftHB18D1vOrWIqyKchlrirxtaDpv
+o+X/jJMhCyNjXD1pKnCosibOYAkmMPV/fhovPg7vkt1RAPoUOPLxpFUIeER/RFQ18mEfRJH3iyU
xuPPd3/EaGnSTfsOnSZzLGBEARnTh2I79eBfkc4OXeDvmie2cy6tcKnhROoJuHf3geR9X1iXpOxp
98jLfSLV3yivSrzx98C7aG+fYfRFOB/mjgTrzYW2xX/vdPCLuyZb+SmBfCT4ljfMfpEFCC6AlNMv
CMiygQOIP0zHahplu+9db48aGC/Z8pU/SZGzN4Nvhd5MsuIo4qFNirfU95G9jEdbl2C05V7CXLBB
fR6trmuBOfgvG2LRfGRBKPC4/IYz0t9n9PajQA6m225Uv68Qa+UCcZH5iV4lqKvWJClI+C5lXh6w
udLNNok/UR+6N1UfUunq3BVhpvMtm8ewgPN9T2O0GcJrYPyhk5eG3TzJRkklaSSZAbSjHU2RSqoj
4Mdk+sX+gVL6rtKP5ZMzKz9ww7p6nbDDUtzUv08Zrv2MRCDPvKftsvvb2Ri2VBwh7vvgn6ZbwI95
q1AaB8ysT5wcrbjh8YWjegKAHt2CDOlbTizqDILA0cjjQ37N6bi2TpAUiKmO4NVxomPKeAtY3bUa
9luCljXfwgmeeNkdgrsIxLcoHZAKbK3AkjQ7CjTK7OD+BlyX9j5yOTSRwdOQPUWaja+2hgBenuYg
IDq0hsgT6t5Mz+Dy+y1YP1Cnz4YxzSQ9rJ5C60i+XY+FuGKxfysJnKeEqFpxwN98h3MX6o/7iwHg
t2D40bhocztNAJ7Xp+AlXRjTbz8yrJklg7l90FMkNMpash9i+uB9/uUayCxQW0KZzaIv4HNGhkzT
oqvr2UwQqER5O4UnSLPmGsk8MsmeAwovaq4Oe5SlqSHrP1O+OAb0XH7H3JaUIKvLH+FubU0j0DuM
bYc5aGvmRAWjI6C+x9ODbuew++4TxXbKnfk4Kp9/KGji0Kzfr636zWDNOWGXGQhEPcMNbuABkr5g
hQL7s1vwJmI9UkxFBYCFtl17eZ1f+igh8N07+FtGNg4hwDpB34Qvbm58Zki3MkD4zUCR/du45Nlj
K9Z9qpy5hql4hTgKlsVBtoCP3oPVNXmWjhJTyR2O0tpgCbuoMwEecV4lJ44gEFXvRRTIj/p2WZif
EAZxCMiAtLCJRBRb6qBADvxjIbkgVSEHaJBnyGBf5dk3Op6ad8hsN3lyvbmFofDVSADNMj4bBAEG
ZBrd3Xia2iMcelViVPwy6Yjb5gmz3sf5BKWAaXHABMjEZfASBZoHXqjv+I53p1APnWCI7oDwRpw3
u7p9N2CxzXHfXNgLHCfnUej8aVv5LvEmcWw0WooioWuRU2AbISEhkMlOps5IdfRHtnEjFciz6bvI
GTkLxeZiOFvV1HngShQ63vXKNEQORCrvXx/u9U8bdc+koKuOgl8eJXPhBlWF37ukD3/c/nRU1dLb
7p+RJVIR9sFsD4NYFhUMcNqIv5IytQbLxBgDQ68jA6Gqd/58QpNE8C7bpWH8YQkayXeiPUEJ++IS
ivQ9J9wYJU6vtGqe0kfcJ2P3DukJFhY8Q9/cmdSk3PlD4YFfmSRVetaBZY0Mj7EoZ/sK+iQ20xKU
ZqsWIDyOGM49y+p2Ronmurwfm0fND44Sh2UNTGUQOZZ01sMox1fzcUjbJ/g8gCOJzx6x0gUvdFkq
qbImnQ5urkSoX2Ek65UF7NR2DUKeg1jXLLXsGN4VLm46UBKrqGUHu4vaPktuCrRIpC0BpSCLhF56
LVVyDcwQVSPMUPoGGbVZJwZ5HGexcmAzKrfxyJxXUvL06zUuj0lyhDHX21mFw4IOqVe/G/j/QT+c
97GkJ/iEidKfBuuW4efdvJTYgmsU8RNd+zP2ZYmYZjl15HwOz+2V6M+Asoz2kWPtFI/Ty6WCjAR2
SpkbpwFCplTPYmC9p2qE1KCB2ToO9QeKu9voizaqEoCgUu2QBJQ+z2DQ+A4mvB07PP+mfVx1OUT+
dj+LPF1asAUy/+bQVU6NubJTLxCF+VXupskrcWQSsRNgqcJiNdMJVnpxcb2596L1JLcXhIaIGoK7
36+jVQ7NoGuaDRjvHmGCQeCFamfd3x6LGjepJWSE8+5v1UXdOUrVQFR2UOfwdNAdr6jWTE2a/nMM
X3DoYAvKlSwPdXVWK9Uo+LrS1cJy1qHPGW20r3+KumY1T2ycSRARo/uAXmUWfcFtTN5xQAqSqNDV
sVS+FMdMtvqdEWBG7wNJagCDoalaok4Zfq4o32MFM5h6kmICqBqZULt3YTYxuCmS4s83gPNvLDSc
GYhnffKFAXLEjAf/sW7RjvS/gzwNonwq00qRaMpTpVsgludM4HjLYbHsLJrsaKZFkknuqLQX/fXX
uf8bryyONuF2y4QHQivjpR3i4ON+2jUtCxT/n5/Ki+FkxEcuwI6VlXaie9E6BfKAirpB2ZT3df0k
hQitnLU2um6aJNq9uY2He28YKJ7QVYaB/1MXkjU/2I/4ZoLIwdEX9NHU1J19ld4aDaowROfYDIje
YiGfnoohofrlr2/3+IbKWIBfgrsUJ2hhpfqYXMhshJs9cD3WKMo96g/KrhHrtKq0MYperBXLMTD7
9cPJBTumbEZhfILV85+3cND9LYYftP288NBzVDMTmgy6XXPo/wSAmluGOYp20YNPz5Zs3GoY+lpk
pssY8p0AG3FFpstAnFPtduOQF/wWMF223AUNr1uWqLYgrvsARLuIAaqXy+BH89UZUxtnNgK9Axjh
4PBO9h12RqbJQli5syvwnzuS0D8bQlM/+D3+BVWIDNTSGkkO53XjB4xR2jsuylKO2yGL9YhsKu3A
5OwgCTvHEjnBAaX66MSoQbTlREyUpELUhbERazmQgY+Nfv2pisFT36phCBA2DqJK7pY4kJts3wGJ
AlkdhGjnpyeO69miFXuwWiSR3lyRIwNVNCkr6NBsqLYvvx/EsXGgz9RdwkiruGwrFIspZiRQHtUx
jitxK7L8Y197Xzf26TREmbPbhcX8kaf4jFyooYrbbdRDKkjVqA6xgAwJn+d9p3GSG3RyyrSOhjId
OuBtLdsfKJmjV6jTab7RJySYlXrJKVJqrMZap1PNpAPUcTeykBIoVrSh9EEpTev8kZ5eJMsZjxmS
O7MPdP/x8q1AmtwgcC2UIN8pf0nMpAlmz45Uq7GlFkEVsFDu9qaW26CJGBhXki47kqR7jktwg0EC
iRNyX3K8zFLt5g038VWvXATlgUygupHpv8CEyMFoqX+uLd9e1+S2bJoZA7czMwY91rYvreR3BPV1
39ZER8i6q6DVvuqgWikPkjfs8N+9ZlRcyswJ83xN5enkq5iEwBuuWIzw71FB2+ICnIjCOPVeBFU9
LFcxnYZVxdOFcMXB+gprjtFRv4kkysPzP5OewTraKnDy9HAKI0wQmYYo/FFQ1a6uOTMipkzhMmeP
9CmBYu4CzDs6AAad/YZWxP6IRfJNEZOhXHlLRpS4atLpqIxIthMnlTTQWVBYBgGnmUsLPHekxhpu
Ljfi/QjHcGT4+fM3GuydskAH2b+dElTIGKGkLHlCf0ffa5r8MmJhyk4ZbcaxJeH7+7hZ0fisnR+c
iH3mw/+d/XWJVJZfdL7DR/3XjUsMmuwjBmwDXZC1UXZHiUmltoxMfWfYFeoExlijduS/RWAW9MBu
+ELAPtGabBV1s4x3nfnoy0ntp+5DrGGmP1o4GQKnbmwvwq5Q1TtcnQFQlj5/Xw8stSvD4otOGhhu
iSZszTlyfYvapXpKRME/c91gp88bDj/IatNglMQsSrJYMvJOXn5sFof/cLB1zrrDjHgLUWfQClB4
AmENZA7w4NBKCczlSqWToJgrN29ZMOPmB7d/RAZi8kONIkgsjHV+Ouks+/UteBSLvCcSNrAOloIA
HxvawClDOPwUHqgYgJimW25Eq2MGdU6kPHw42dZV1pDyZn1x5KCI6Mh9IFT6yE3adLPbeoVxp7LG
lVb3j/segYGYyL9TkPhcDmab3HlBjVXMq/+oXGqE5WEZ955BNctdKdq4lY00wlgH0z8xnNHWjvvk
PuLcXyBaOFTxiLdpuPVA9RBgvb72zuiZ4E5Kck5U2l40Q9Q1OnHe4nFIqjL0u3neaUfxXP8MZy+V
UB4s1rgvpPthVFujGDIwbDF370qkry0iQyh4ljEkJB5P160j4tOjQZrop42N2xSG043yOODRkF9q
jJMAiikBFM3P2O2Z5TWCWkyYTjRewA3XChw8r4wyypmrMK1XcB2ivP5ITmQG+S1ftdEsULd4L/0y
DFyLhD0AD0kj26utloAGkbWjh2ssHwikaNXTFYgO2n7pbuEFXMLtCQpZUrFmETGeBQZhdanwYfET
WOpFO++4dyR68LclCOMPmrNEdVBGPmyiMwPmDSi9ySnuZmblk/fBHZ0ug9QdXHwUK3tT0SmKaaZq
w2WT0/2rQd5AAn8JOxaEJcVEGT24+S95Cr6dUcP9LlI1TUMdzQKU9SUN8GFJlcM5y5rgRr1ctEBs
10XfZfGEc0mseuw0e931Rwzh9kcDdaICnknpzPDZhp6a7bZV465GxKTZMzaO5+80XdTkXc9xhd65
WWf5fpHj2YXPDWXUrWbYdmfC/XHiy/5t2pFfmFZA8PJRrXHOEgk+1XR3DUPE/JEpPwAQBoppJ64Q
o6efujy9gxg1PuxyQhAUp9ZFgjKDR+fgj7CvjSWh7veK5SPD0F1LABS4wPfZ7wKXwKVtl4YJfxEA
15FzREvkZT5yJd2blqi/Ge616eWKJ608cFzTjr1H+XKCyicL0FJaHWFHAyim/K3UCnJeZX+L28Xl
VaY703Wtyf7EF4MQo5/dTWITYDS0seqnKcVvRKMPZKBlF3yWD9yayY663Tjb5fiO44+sk2ZMWEXq
Vo3z7t8vRypTh7ZGkLLiWf5pAJnKgSEEbtsqdBKxM7Y/KZZN7yT58Yedr+KWdp7sTrOW+lIpZowy
8QsRw6ncpzavD/eXpttjQyQuFHtXkKwPiN9sjmv2xQ7kPD8hzrExEyLX/+vy45G2dWNDyBeNJp3b
CRI7JKtbk0/AVKc+Uqvjl/yauX7Oh8ZiL+OEUlzt3PQ5IE3sgntHY8N/SfeNnZ+fQvM5x833/Bbc
Ooc2WRJNcles+fsEpoCj9623VmaTiY1f5z0O8D0bdUCFG+wdurF8w/0+1brBXdr1rKGAjyOcMMH5
+ZecG0Gnj+mHumcpGi6rfmVbH8SOu+YeDIZp9jI+l+YSAQYszhLiFH7CZ+JMxFeXjLQmjru6eJDY
bQvGfFHF20gNEUy/3gEDFGsFo/pA7gNsmV76KrJAhQlI+CHTWQ6OkA41iO2FUqgqbD7+gt0WpIBL
jXJMi5J5+ebKW4jgCfPWQxkxUUJosgzvD9mxsKcp/Y3npiibOIFgjR8TLnizVpfPtwMlMzkx4kir
NdCws8LqM/pTL9ooYfXtEeZuwV0W9ejYHRSeB3rvcJQr9n6KWrgs3fMgzbqCvGV9ChyJDT/BOM+b
j4ct3CAFRgCzyCOfgijcLWbA5kmbuHtqzkB+qKDcyMgOgUz/NHzIRW7M+a+czWRgbDUPOcbxuQg7
Lbyunv8Z2C/i3YgvzUNNB2p8TUEgZ87xHQ5nkskxVaYW4wB9YRwyFoLUE+nbXSNmVNRq9bFK4T4Z
Fh7N1nW1Zo5/xGG/2PbnE6H0YdeD+l9549Ixqwe9kCnyIsVcVYdJkwCinUmb4DNj2RouWBEAxcZM
tE8EXrCFmq/sp9DrT5OIilalOuUyi36jNJOvT/OCE0CoyhmMk32XTPUNwZQqsNhRTrQQBByGgZA2
UF3B0MMQW/K6hEv6gwcU3KQxielfxIAbwQwS40W2zpzcCmtelXxzidGLVSPAEAQTpFlT/4cPwrnJ
ayKwdYtYQ3tE7KdLfwDgMwdX/An2j0sqmiNf6bQ8K3bJwqo/6lP+VF29GVjYFvI+KVErXCbrR7ln
qeMv+D0vedvsW7g27OVdpdqfPZmZSXYTEZJFyRQ431e/EumC2ckLjs3RmrkVmxZ4juK6wrwRZM53
0bg5gxu83Q9LG0IhCgeX5+Rskk7s7U3s2ij/JVRe20QM3ZoF5ttvh9gh5MGrjOeJnwOz13Wkzy5T
C0Xd+EGepBReBpqYaMNZgBvgiQOZEi/XNCs2rjn1/huEO00D8knhhUxame3573gJAtuqGZ1s+VUe
+gGZCoe4ga84aLLKxbQOYzrMjzRng9jiRO7TtGpgGn8okp/Szu4QCJo9BTWNl1mm6/ueilPOHYob
c8/QbYbmFVpsff45knyPFal+vbXIxKVdipF5zhkorcFslaxDuUerNP6kNLH05qnTJww3TDkb7I7P
ja+BYy6ITW46NuV4MRqjFW9uznvAbU7+HuJuc3HwrctPei+lcbOh66pkYqfan8dCUTtK+ILvMRTx
H/CtFPgmV9aZG4qmBr4ociZjOMrCXQdnE+Ai/TONl3V/SAnBlNOEgUat5yDmvqDB+D2WEOKZkMdV
5Rfg5mRc7oy35yp2+SKuqnkIi1AjLhkzqek2dMSJopv7Mmgi3BrPs2vkeW6zxSjmjOmmCoFHgCeM
6BWIVf1TUz8/OomAMLR1R3YF4OleMd+9Nvc4cs+d8cvh8QgIpFaJiIWCPeC8njfJwSVnCHMw5XZe
PVWpZ/v4Zp5/3KO/FVJNQELWu1CXSesmY3AwyCzSU/MVnOoSFdUVheDRXIrOPrOB11JyP9vWLcUM
tkgZ25DeeiRlwnNyNemTi3HQjgRTj001RkbdMgf1iGRmX9xDMWwDSyAdOb8fnTYkygFWnYvTeSVg
vbL0EzwNlroq8FmQRTkrMpxHA0pX8jEkpbB/S03tpIxymrlS+CByoZbb4MOu7m2ed4TuqK7Zt30c
45UytEJnDu58OHFpTgK+Cyoon4iAJEemLbykSLsuP365AQOr008csNCrReshFqq+bNt+pImi4Nfu
c8b0y6gzK/lk7r04ovLtVVnFSjm8sFwhbx5lhkNhRYHQ7CY+R+xStHgV5A7oYhY1bG3qoA9OUrwW
/FRfL56I9ZpQwAeahwCeiZ6O0O97cMHdzzXFo/I8x0ppy65NYC4cz+oEOP0ra8tgWay+wN4W/DKd
WtmlFjR4BcSMZYouRYWllgezf69llF4PGMuO1hUE8+VzFHv9YC5hs0Lv+4Ts432ItLTOwFU2P5Up
VHrQgfR1gPihdFR1a32USB55SrzzFB2cN/p6zKG8ObiBFIrSQSgvr7E/etZrKGhJ6oRuv9HG4+00
gbNHqGzGtccDToRc8GtSNjsbQwgLjIoneqFwsDejguw/POD4iO5AauFbiqBtixcBMxNFled9z8OL
voTbs8y1ZdmgstyGC6xI9mwmPJlTjM/8WhnhFPRWkbGeJpitAXAoUz7Iq0VpIgfACVgourwbzeoi
m7FA4xPI4dUMpRgXZvQEpld9L8cEyUp0Mhl8q2u8NujJcJwsqEYasdXzjHWt5oLSUlXE/6QVKpU2
iYvhZPTawcaJmaWHfdpnbiMpnajwwBNXMbUAMRFl5VFcAFNm28sVDwYmk7BwEH/ddNqZQOnN+vS5
p8MXds1flRxbqEKshTc9LrNNdliBo9ezwFOsFBsxJysfabnB182h6nC2ODYMlAJgIn6AGGMqK7hb
U9vMiWk1SOk0+R4vYaaOFoS94bOK92PR1vkYO2YIYqQGR6KllpEAb8P3QpQsknWNS+UvZZBL8Q/m
Z187VYVftj2nMUHRnbFFiUDUFa+Nds2gtKZxmP3sr2Yndq28nQ7sFDxWa4obgctJG4VkepnAFVpW
I3P/r7gecKO+5Za98EMriDypjwTWP+K1D4FCVLd8zo0qQXFszlbvSvGRkNPMIsihnX59UMcM71oj
/wVo2gB9uX+nPtsC1161jmSoNPSUjF4mQAfVOGQqTaW5GQXmjAUjeOQc7IpA6fy3GxSksRjqLNBW
WPpmD6hhUtq51TSFHABpwCFihQb1MSE0HPSmf5PEPTkq+mY+SwCJuvSqHaPjHOpPy4dPqQlTMm84
L9xNWhGCxQW0EqddifA4LnZ9W40gUcc8rnb+8vutBQ8crSUTdw4w0VQzn8Z5BoIewskb5vcd+PNC
YnROBkTD7OZ1MVMt7FtGBXHELQiavRuT8mXlx0S8rA453OOGXAJRJx05/+fhcnCZnnTGraQJAgE2
fMuPv+f+JVBwc8Y4ao75YGL4MaMYxU+WBmJ4UFcstYLdLnzxVz6AcrGIxGP5PmGXbY+ZNUqYAOab
okfOmXh+vk3YmgfR+VN1Dt/8u4QWD/qdlBwzB9niwoZGc6gJdHB1s+UnOCQsck2WgLwUkQ1bzabB
zNtLykrUX0wMarIG++yLgomWDuvz2jtPbpcJoOeY4Ty4AiL5ziNal43ttDiIcauSa+ZPsSo3EA2B
sWkb+dIikcw9ELD+rQ+aVumzGOAE/Ef7Ti4qJO9QRshVMzuV0NR6TO+AjUIC4jdEO+IHwu1A6zxi
smdOqlwfIWsjQ4XRYaShvNwsDBcOkUOmNf2/WFTnrbyI5mSUH8kp0EYD0y/Z/kALQqgeG/MJvp3m
U+bBrcX/3T+sndcU+qwYApQi5S0vuhfLdlhtvwJN9r9OCWV5zGIXbN61pIkZO+Mj2xecuwUAUKGC
uFO16XFbRrn077MUXlXDhqdMQHvn5IJEw6qzRGPvVScuIaqkSxYPtQZO6hKY7Ik9xoLtpr3RCm8f
1WL9kdNlaQKCmWi7YYzNqRyywjeQX9QbrgfuXvQO8uHe2aiEqmIAEIEin820u/9wVtb4LDyGZlho
sOyn/YcSj5XM0/W7gNw2MR4dGKaSQxEh3sFnS9aiibbpl4y1jF+BCbLxaCcGuPT+XXvA7Wfdo8cm
2xFDb6hX+p68yzrEQizjFsn9F37Y5pvklqJNXEH4xahf+Sf07kIfWdQ8haOMDYMHLnmdXq27grvS
hJO8udqN2Wt5d71uoi+UU1Gp3umH1sjZDcMYAhxKU58PS3WRKOVkK0UUtInGZLtkuJ10GGwlUOhd
NxsbP/HHzWf8+VsUYxdzeCpFZ6MpRjFg3B1lk6lQ0+Ipuh0vIopdDDZwVhn4yL+skYoboJEj2+Lf
UfkNjwV4/FyOP8TatVM9aAZ7mi9tu7KYD8qZ1bN1qnT5GZ76oiyCJ6KxKYzAx5wIN06CZK9GIL+g
0QKVzB/CSsQAAbxSpEwo4YhOPp6ZTE3iETdDMWlOfaRCoNqt5gkGSO+ZvS2qonlS+ZIsik/gm2WR
nBeIA6LQBqXBofsfMNnfi3HREx2rG+XLaNvyTfj41X5bwIkvwKdTRskCL887y/ZC9I6aWJ+iBoq1
mhVsZAYQ/opk5/0yvzRMzb0K4OelkO/rxSj2NvogHuTfW74DIx/JhR4NSUFMjFDNl2/nSQnmQn0C
KiTiABIkKZf4i/KeBsV9m99C1E9pJd3dJOTeiUjp72GqhzRi2wlgrbDNAFviPFCDFT/c6H+l7qCQ
dHG5vTTVppZcPYwD2krR00tbktKg3PdSKRgZ9Vt6XuFrObsasZj7s5HU8WcvNba2K6Cc18bdu/Sr
gptatGFk7qb5Qil/zu5Eqx1jBmjX44BJMqQcwjPP05CNiOUFVlpyw8Q3NemULNP45DhahjSnA7AS
M30k4bOWIUyWbUem9OTTgEHKjJK4a8jSpPKvFmjrtmarvPz8ejRlUtKy0HmSDJQsxENWXeB1RhIu
p+Cec8f5uUDAZvs9OBwkqunZO7YNfvZNLBzOrtu1siSesBrqV9jwzSRC+8KUsdczUZkwnRTbYcuV
BsMnRnDc89vZ38iB0Zv+pVz2M418ELz/dCPZIsA5FcRTPtmdmVggEDu9YsPytwADKlZrbTS53dx4
nLCcfTt5yxOlePMGWQXve5gxw4wVlIHeef7o+fxoLmGQOzW8cgaiA8wY724Wx1EaQ6zcrdHC5MTd
xVuw1IEfskwZza7UYPjzIvbXY0lvvc9iUDhgZofGYQLl9crz6HZ7hKnG5nWPrR5OciH8dWNYNw0a
7dPh+YBe6OyHKSkp0BNZL0dWQliX+uvZ8l26Gnhw33VqpuXkIb9NEuCAbB2szXEs3QaY7Zs6+Djh
0ZbHDqxoIrFNF1OtaSZzAE7mCAXBJVT86EwQLZA2lI873JXYA5Sp/xfO96ZJm5gTlXmiaIWBo21U
vnXcdG7uZP8SY5QhhzsJRaICkNXNHCQVURVbF+F6PeyrM5WSASjMyMzXk8ClUZp5259O0y2sp2fI
0a1u2TdJ7qCTRUI4mylbPmihuViAaxP6XMgm2zDMfM/tp6k3fM3Yc78zfac8oJ28tKDn3LeGU/qy
ju5/nnKHUY+5U8u9qlQ3qQOTV3fK7Splxqb8EFpYQmA1KC3tzpan2eOxqbqoM0J5uiAmskEloGK4
zXrJueIjBnIJgJuJeYXnIjk/avW5q0TlT5iJLrrKa0Y2NcA3oqeRG21+siSgIPSgRHNrpjpR1d89
DXu2ecgklXC1X0qQzoZeNsaBPGNt+7hspCxBgaOpqJZlDvKpBU9iO8ocJBZFn1mUx//zte7oslh4
Kx18YQtG1CpAa1Q+SNcoWWh3cub7Dqn5uBVzQvbFL7P8YEdAocyobIV0bhZf4bLeN027ieRvX85i
kcHqcWP097u1JnFCIGT8OLKWaPF27eFcJ+kuj3bbCH5Km43tMlED1luT2kRqI2mKr1wdh8eOUHU0
M5I0hp9/oODNQjCUfnRV0pHt2bQUsNr1ebxmxbXh8B+8xBovVtlT0Q8bADMPNjthkGw9Ab55FiwO
KEAIrU466aEh3AgbOFs1scQR3m1pXUlIFiNN4i6ULLG0r7FGt3+0ZrcdHlDoxSlbGfLagz5S43PR
U2s6UhLg+KoJJZfW/tDJJn/jH4rHfEt5uNLYReHEIMZTgwtts3KavvspXzAJZIMEyENDUvGvC8VI
T8AkPw3K4vLnWbd57VCIetO5lxP0Oj9hW/oyMPo6N8emzrQtNo8xLE6MYirLZspnPM5MORJtAOx2
o+ASMQr/GIqIFBE6aAivCTsldXXBKvPyipdeRWdMTGTbM0FLz1fZSJfi+uSTNHUOUEGIS1DM8urD
mmuYFu2eTnUXJapuExx+UX2iaBbaMHltC4D0xjedKdvRA6edpk4jULWKMuJ5EmxCeHm9dzeaxXd0
n7Kp27MvXpnAfu3b6xzmv/G0Fq1ZbnlWba6CLOqBO2nuV1X/SjzJM56qtLm2WZG/Kx3ZghnEmi3W
Pdqltu6KEy09m0bwTDsOPwLDieRTUT4VRxbdBQxYDPZ5invbeaocO5SuMAjbuu51HumSFyuSSJUi
RrNXacVq61rl3GbYSbvKIbUmayYWPFbsB1yF025m+k4ZVkvvXHebeqo8Xq5mtsVh6RJocRRHS29R
YIZwk+vuLTZ5rXpt0aJoYZ5uTcxcj5u3RUQBdZpYJh6m+NHzLd6gP0fgn/UIaOS4Z4jcC9fSyfic
MSFCemjcHtazzDpD7HJQPdRw+yr3oaa65Mu3RCj1Vc2lBLXLc9U62yvRwTK/n8mL25ZUvBWYXY9C
YjWo1MKKqI1JWIBG6CGBqL4wvnb0Yzyw9e1w5auRCjtRvAEpvVthoYCQtqyAKBKsSMByW3FBCmH9
Lr/pjUu6y583O7W0mBK5TewsIDz6Mv5FWRp2dNcqY3fDdLSE+V13tvFTYrs28rI0kbiAqaoL/ht+
xHB1GICnQ1EiyRs2vzfkyAG3WS+kaSnTy376PBDoQodK6wOzCzvlUPcYl3mkRvS9xjt4zZaGTf7v
sr1OkmvfuMjSYGcCc2HDqfsZxXy7HcHXgqOW582dNXUNgxgDtnKDc3mclX50pWtJWdZSWhVQ5hM8
ZPyZeuDnt/xQXLCKrV3xiIjiEDJ0Z0E5qVMBM09pIqjJ+JheWTle8DRe5On49L2SPyECTPYTbgkO
KzYvGv3OyV8RVzPWB6ZwNbQGsNAnT/7NPlinzXyCJZCPeda0ME5mHNvDQNScqnKPJTaWDd8RJ3Xh
YYbdujnE9l326htNIFmyAEqZWaSgSmfl5cmAjXZj7EUOIMzrSWSGWoUSGh8f2bdI6p1sbquVznIa
48Yej9IMRo39rFwpk605exJ/ujNVGkySLl//Xte9Q4C7GSgvK0jwsIHWNBE21hmuq6m2w8Q0wP8F
hceyZe7P319oDQzD6JPZ5u3LLYSsI48p481fuZxDP/YF2yjglOKgEFrQ3JEzXmzy7chWYgZVbZm6
4QssfPAdBv12WBX5MWQhsh0RKtr6j2WZhsPCU2E2rtvdF1QG60L86B37exuPOY7EkGttdtbtYkZC
smF/f3+hmWyJ5izJn6RcG4uFcw9u1FI9LgBK0kG8Px3WfmJ4+bNJXxh47YsN2jMdvA0wODn1G3nX
0Gej80N7Y3bwR00Vtp01eilYD7oECd9h462JGmhCNcokeUzeH592NciUrGSOsMgOxSKWskQQYdbg
89ogRvlZhkgHmcC2XQkOd3zf/TObhY+hVnEjXAj6XdUhwnhhXaykGu+qMDtcGZEzNtzqNVlbrC3H
TLJbAjdHrqF7nTlyrh0RrlfFHsr62IBR7TStZ0OPiczA4q9/HJXFha0QiltNis8uofY9E9yTlCOU
78B0YPRTiV5/XsH2dlS7ekOFp2lTizdXRQDfneYwik5Tr0SKQ9/q1S2Vv2KLqoRsQ+ZOHzSv6G6Y
wz6gOpc2p0oSBbui3LOCNYq+o/XIHnj9y0uIzUGhVB0AG2IUGaq8vS88mAIfdJPiSAB/uqZsb5l6
ujXHKUoGi4e2XbRHJCyTB9STgL1kqHNr4MGBJeAFBmRaQe7SX/fPt4U5vBBCQPBIEhZSir+F6GN/
RjTQV6nCQIUIv9Il320PZi0JbixCpd03DhgzEKisp4B3MVUS7WqQZiXvM9ku1xPckOo/VEAlCqtM
e7+XpexK+0OchoRdfLyLAOXhkO9dr5cMsyg+1UOpi0mjXOWfOGkIggmNeivwxgWAGay+BNJdgJn1
FsBxS+ODmK7UcqdAowVasA+xArclus043uF20exJ9ALOm07A1oCjImmf6i0drmJ2qYJIKnL0i2VS
dyvL6Xbu1Cj3oMBLJ8SbupoY1Y0og9KfBe0X/Y21/VhEVxisQJRkxvP6HyA04Gm25fwnM075G23q
acpG8l+dBDD0YbPsbtBxOsDSa79MV4v8/9k9QhrnsL1kIjigvVTQ/uphJp9LIMK9VfZZ2YP+6rMD
KkPgEC2Fd6b+qJ09ewKD3o4b7tYqG9HFxEXV0vhScV4pgvJ4AzWSOzwlotb5YOBsCwyDfqLOX4jl
mxb395xtC/g3GtjHa0OMqqnoPjGQ8ECFFzGWHtLwyPhFWkMO4xFMySlO9SaczTmCazWXwifl+wOo
2W2uUCdiT7vK2OUYTueIqmZG7eK+lqDls2xOFdihS18Gu5BTYcIZrMB8L3/HwoENqHikpz9pn08M
uyz/WwozdyIXW7YqBSx/631MoJYJ3zTNCIPOpG6iQGYbchAkcIw+cnOUo8I7p2NnWZtvJ8FrxEqC
KdVLhBFNKl6QUf6xL9frLyhWJWtXYSsm9NaB5vjOdW6GRtFYqDhlSR6nUaNVZo3SSBBvxN5Z6hcB
DlOz1LlAp0XIKqiDcerSVGLLyP0OU5ysCbfDsPFVOzofvcmZd0MV0dWNB5ZQ8LumZzYo+KwsDNWR
itzWwwAT7kr1tp1LLlxiO3t7717tsaJMQMCR3dNy/iRS91PGZzAWUK5mt7xRAIfAL3qnF9nTE92N
08O/lrUWp7AGyDVXVtgyGPMUmDsX8T8wPPG5syMo7WU/mJ8pfsOdhGTZM3ZrWJTPu8v2iAFpYpJe
5F/s/Ev8T2NKIorLg7kFwgIsgGekYtoE6yeJdZMpTjTxQlHvz2RWRmJTTpMog5BCveNqdc1d2NK7
nZK/lt/DhEx9rJl2HvneGKXJ3b9m9+Fa/df2iYPYv6xm+d63KaDVaR0nF57wolUBCGsQqkA+RlPS
dGaE7zR6ZfBh5NmldqjjUnsOHhEBLZTAsOfTLcJeYshHcJRFsRZlUoWjqXSVG44cngFHhijRwyFg
DTJ8eXN6Zu4XMIKYhQHCs3u3JnF8NNNxq2BSw7cyjjhRT4SuYlo20/jyAIbPJYLTfHcGSQlK8GxG
G4zYpfu6jtJ22uHLZnWMvFi4L3songbpEWYkexGUl5G7ZfDWFWrMgCPVC5sfsDXf69aXIRSVN5xb
h6vArRYoT7HZdz7rfjOORVHTxPXb8Ry9gSYMUvxenryBGJpyEDQqybql2NGT/vQhcIBhiT6bZKul
Pd680p2kORDxBEbFCbi/IJNSN3DvspXjSvckOlxJSxytcLtwFTja5ODRq88epThGhAqVxIJbPFJZ
oT3ojQuNjjfGsc4B1xPoU1qWQN5Y8EWyYtNV9bJZWVgkXqHd1/B+cTFYjeT8BUKW5bnocVOKH8nE
r50K39d8eB24BfMjp9GpEb8OcCcYNsIZ8F9x5gbq5OLEo+L7iTU9gvd2+3e+wmAOF6rf77N4bpAn
nGkTPdX/PLkA6H6T5JCPTQXERiC3yrn196QVjc938NoLkqEvHiKRL1YZHur99xUBrLRW5kEK6RYL
7cbR9vFMUOWiHy4XBYpd/GBBV1R9+9lysGKN9a7CjZIOF5OyL48xwkmPCDmtQlTaBOBpdHcWno/n
1msG6TcJKssc3FjPTvuZsMuIyFDzTczNBLwRoqqJWCR9+RkDucYdFzlhF/Yt5phovvUZQ/O6AQ1s
C/lzwy5PRN1ROI6pyTiREPLtnHdGbkJV6Hl/cbrJd/p71AyrqWridfVjBhWbCdr2RRWZ6O7qMojl
X4RNi4QfhhytCNlSo8mkBBgEXF2SFccplacMpnYygnQH04gxqsXLvToRUuXzzoY3501sWN8oZGY4
WCk4N6v5cX171h9nB6TV/2RaTwOlLmaqF10l12GKnT29eIa+nivA5WhQs+gB45R0meLTJfZM8VxC
W8c/eTeVdW3lJgedb0h2ThDdVDyvz1lIySumfvFgVCwy70GJf0NhW8F7YYvD2hirLR/HAOx7T+E2
pUr4pKWC7dGQc3H6+/5sgPXBySvt7Gkxl477LSYVBY5f9z61PusFigLCsZXXokMxy8zfTbk0RdP8
nF/fxOsUYxqcikrYPBzTApuAb5ptpgaobPdkv16ypRVS52GhdEx6fh/ITRjPuWV7H3EklNFKaWtO
txtZyYeElGCDLe+cl6MYwkIIXtmzyr0RGPSE2PXUAv/1MHAYBTM7yIlZ0LQMtTMCqAjIs50SYzER
5p29IIIWSjVYVnv8Zt1zjmntbvK7PyvQLcDbXbXBiBmI/1ATK0m0kooTVQateGezACFFeabuGg1u
HHOy1ervSDj6EtmIzQoTfrkjuz7+tqo22lyu2V0+HHw1u0KRYwlRohhpewLmGpt6Df3iloU636U2
Izkkp1/ciQLwrMtQYRm87OXNukX9ikkDoXbeUy+v4glTt2xTcY2RjhngEyOaobD7kYHOTSxbgrgG
Agp5YTnxSJ2HEFofQPgJHssmiDKlqpvJKutJZ3cJKOrfTAcoL8oRq4bDNoQTsEIPB0U/4YoOQgEp
NjzGTT7miAXL7h+AQDcZ/LOO4qTqSq+2ExoKc+u4+1NXH5lA1hwqBicSF3KR1XYfFk61gkRhD4dJ
j+6QCma6dLyjzMkVuotV6WG84/4GvwJv0EACytEsLxF8T103281mk3lGloovg3TN8yDfulTRMjPi
qP4U166JaZX/ZMHNU3Ip05WCjAtFPlyeI43WyAvT7qQEpHUkcxWW7uawA6+0RSrI9vCyFVLoFbNI
XUF1XkNioseFTp++VAxZyYN7LsVgjQEUc0K32SEayj0i2A/osnh7EpbkeMBC+NQpv++eMrn7HZUQ
F4XBuoysqLuRnEs3n95nz9oGytdP+yZHZiaRfj7uwJ5UhO0uCPKmciz6uhzFhUWyw6c0SSbM4nQC
pWXdj2LGUCppQYQ6ZVh385rTlmH5E2NIOmzgHycQFrwW4l92GW9h1jMGjG93HvcnQEABVSFXGuyI
xMBGEIuD3DAiAFiLee6Fc+EzZqGLxtz1m7oYIeWdcXQLymvsLnK921u8E5bvy7IbbJbPSL6pOvtU
ZRFL8Yv3bWBXxiAaWz40PERLDfn/v1SGYccNmuB/wkOw9/87XY7C1M0Lrs8J90AthqKxTNC6KbSa
7RFNIB/sGWnCnsqTOghcjRhlcOsR6HiIPc/gRiCEbNZj53FWowfpg1O0aZmaBRAJfiuKdo8jcwQD
rqaOhpROCJ5tRlDX7OZAbr9uF7AhTabhx9Gy4uMTEIM2bA7TuocaZrBp0xM+Sbs9XqpFMP4Ac2eH
CcFkAamc01mpp8ogJvgoUf69FMSMsQ6F8Ovi8q8ymZJ7ixNt/ixEOgcK7tDZvNiNWbsAAl7603t9
FG+39ANF5boA3mRFw9pO+CL8vrrMBkfpG8gN+Rd8672btXI9bOOf+Woo+63tnyMCGLmZxBEsfvD2
AB4K8fMWAPtA6gjIeOrcEMdzK1sHj905XbDAZRWzUciPl5dchCHI/QHZ2P+xLyC1nzsU6ZP8ZrO9
rdPOqRKPFkyJ/mTCDz7oS1dYXhcwFj/cHicReWfUw6R1uAezKx7ucoNFLEUPs+UGEX1LWFKwjj2m
SW2o6Qn1z79JYfXq/OWG/ax+P74CQmIvUue/15UJrerlF/PFi/PBmrfOyEUBD6bwWAdeHcc4/S/H
AZWzC2H3UDc4QhNRUAa34iAvgrzSXqQqSs0SHBPHHTFs+71giS5wUhisS00YROteK0HDXpFqBNqn
rpyNRX7qNqz1g/pX8DiX1iw/vESEI69ZJx6PDi2aVd7eKj+UL4h1RrJVLMXAAtG9WfmWWjp692vz
lIczOrtswF/TEKB8vKi8+J+IPXh+TLTmVXYxSY8X3PPs+NXA7jNt4Iq544/mdv12I94S9xkPupVj
wKp3KV5gQ5roJPHgAfrnrSLhF8jUToxLZjWtm6/LeZfxGNM0/cOJA72jGoj/F9Vf/eHf8yvDmlJ+
iM+Xmqd8wYBNjILE8n8PYVEmyjHZ7dZ2U8h2FVs4mRFL06PPsBmT6loM1zbyVsyX1Zzg85vO0EUQ
9PkxSzzV8jlJSbfHugIO01oW6NpDMpKEVwQGWuGDqV22hx6QZq+8q4qRAJ0+gRX4WthIhwozjsx3
M+zEOlNDnU02rGe+P7ap63O6jF09M6cbqWTDwzgMNnykG6XGoSimTl3HWt9Wm5ogwqgvQ1OoD+mm
j6ogwXfdc+k60CimNd+5V7/6uBJKe2ypNb1vZeFSDkUl3bzN0RRl3Ah2HH7Jf6Iy7EBYorcraiST
zj2MPMFvXNtADvuXOBo0aff+7iCv19p8UQF7KQkn9NFsFWtiF1EnS/5+F1Cjsi+Anxa8Bnnn3Yx7
8/Z5fT9QWBEfp80VfNf1XdR2mKXuNTOwLIi3OB6vlDqopmycB/bb8xkucXFQfG93zHoW4Gcl4mF1
ityT6Zrbn5ICG7X1Js0k6dDBX2QybpVv3Cp6ZBbFe2l2BujDRI2X7vhEslWKhkg6wIsS1wOrqzuV
jtdMbsAbJ40nwwFi0Zs8FgN5K2j2MP3FTGrLMNfYZJd5jtnKiOuM4iJZ2pLiz28TS6nNjBKlHSTG
lxoWkEZI3CFnlunpN2p3tuVmF2kZHW5TyU1GNkMvc5Vqdk8U4eG2kXX9g2ElL529Ofiwu3l7jBB9
hfugO1O6kdAziuZrJUjdYSHMvFzODAhD7MZUQwxa9Kd2yKR7iYS43Y9v7NgrGUb8983hCV1T4sw2
uJf7gkcmaa4RbxzAk5NUIfS/yTXlurOkMKEew4tIgVyCaoOk4hRZA0Efnh0FL9AxaJhSVkOFti49
AZX53mfBfI7eShVJ5UP4JEXIGWjCRiy+tQmIzV8132ODvqmPtSHz+lVpLytrMQ04QUcYl5noTN/i
WjgmB9xzUnL3BUCU5Fw+RTxyz41qhxeH2Y3F4kSDskrxj1x82UIE4Jwb3JIcA7bo5vnfnQdu/j5O
Npe/cMz2m5Yw9GZ5X8wo9NxSY/Q+Sk/b0RejTyzzjozzTaB+gdSVC/5+KPvuBzGu2nTSghA5L3ls
Zh4dY/WgchLCS3q0sx9+N7DYgnuiu/PY1RWlxYJHpmZfsYV18HXysj50njUp6aNUaT3qAFEBfsDU
I9FvMW/VbRq2nxZ0l47cgfgTIvfCHrFPq3d2o6mAeVPv1lPfUpNvwNqp7HUd5abV5tbr9jIzzbbh
dXs2+U+bXhvvrwODZV4VWXId4/6WFXwqC8IX1gH/WJVllBjEm0q+z5aYoGsznUXlHyro23MOEVWw
oTGxEPACjgLUs5Zj2t5/UdULrtuVzMrR6g95T2PY9THZcShDrNTRH6kZP54NBI9XJqJuEz6eBWmO
TT3YRsGPQEKoR9qwZ5Hv08LbWtVpKzIoWQNW8Quvd8bHY1RM4B7KRHMPTx5fSPgytlHY3WDe+C6y
1wQta2QClUl1Wy6cO8ojLaeSy2J/CuWuLdoho40xHQTh7yK0J30pJ1T/gFB9GaYPBw7CfazQ28JR
pnoP6548OuVC9g3Mh/s9ZR3lo1fc76ITgDxiysc3kz0Gv2TbQ4c/oRbVjk7ipY5W3cVZNTcC72sA
JXN7aV4Fth8rtDxW3FA2FbErZoN3KVoNzzvHuLlYzIEfoJxNhKlQKwOoEvIN31fJnvjeH56R1Vjv
g5RLmhGAfEVDLbJWr6Hx77BcvCybqdEC5EthOL+Ilydaf/qP6il/1b//3bt+laOJK8SNoSpWdf+Z
q0Ix9zfGAi2YNRTrCKPSWMRHJBuFl1n7MJUQCqhIGo24jsZhogzJdp3F3PdYwbZ8wlO0QRDF/pZs
q05nTyz86WBiSNU0shAJvyFcXGSLk39OXwhV59cX+gJbhOEt5po0E9J+giCi5R1ZifsudqEYaa21
ah/UeuSz16bL/TPxeKoz0JmGmW99IPnam136MEnTHbhvF/34U+ybRAmqRnOTyLavuKmfwjNq/4AW
NS/prpLDUzFmfqliNmRInf5Z9cGcVeeQGScQSrz48wjRMopo2tAzFXHcIjAWdOqUbi2Epxg8vilP
ofKkDONcZAllxxn1EwCj5CKC4sSiUHLg7uOioBrb6Lrb9P6Xt42fewW3w5KPzXFcQYMePDW6eZqs
scPINJ8i8LtnqA1kSKZCTN84bohk56X/4Gj64deYWyk6qIymZ/42dKbVWPpxfROnShW6oYDZblFa
ZCXwZNRzzPlGUrTi3J3/LYAYK339A2PuItMRzFx8jr+NtzuKUGPtPSmp4jX3n2JR84e3x5zRYzFT
zH0uasBBs9znKSfpoS5w1EPssvi+0GGhvcXPpuHh8zWRV3yHR9q8PBQ2IsqPTxzk1WMC4FXi/8Aj
2emCH1KzD39JDASXiq+MWtpu4uE4Uc8/OiSsKrJ2XGQh6GFMhEDbui0RBU8kgoELIPfiioXPvItl
LWAIBFJ+VxI7Rc4ZFJkmz3RsF6MNVbs8Ohk4n0b7V1b7o2XXrD0IBVvXtFv6ywGweRMcNvW5LYa7
3udwE73puF3fP7BUi4Vet46wend7pa5ud1T7ndQy/zGO6ndXPQdHvUThTH+tuZVnRCbcbQWLh3UW
sOMszQR5XLokRrcQFtSZE2EVv4Y/OnYnWtXfAw0YXSBMwmCGSfaXnLsoMeyEHpYdN+ud3mzb0VDU
ibVlPCGKfloynDQc8ZaoBaEHOiVzMLwhy81VMM4bufPEteprYQ8GeSAs0T0bBDxq82hLmiUa+y4k
XtrvQyyFP+xc2WcANJqBmnRsr2EVA0y5HJTK5dejiehGFT6rH5uSKVyc7JvOi2+HWes7jtU8sn2i
uVSX4ED19HAQYiiJyE4SR8ufOyojYvPuqIiCiaA36O6wLuqYAcHpRTWL+6hR5OBsEybDjpTdnULU
QA2O+x2Xr8nm+O1R+fFAs505euuB8X4/hRrkF815HL6lnjrBlQOAOIoYy2FNCHQvLWyX/OxZ2BFq
i/NXgrAwjNIcaAz1q75y7VCFw8ZF3dl0FnQZNeN35FD28HKFJbEooBSFWSgLpRA4rMHPLsCN6hyu
XIJzEdTIBNV+Y51sN/vhFlTmJVpyRVPp5xYXYoAPijaOriak1+Exzsi0Nb/2hoY55DUsxme5W34M
/JUoA8+hn3XhUcepNj9ajq9lqBVbkpHfZFrtMFXssGKnd8sFP1J/mlvjH2iAVu3JOk3pP4orTHDQ
sQNEcPb0mGq+rWNLHKi970K234ZjveZZtkXTc0EJphWkMu/lUXFQ1p3l5VPjAt+nrNwBfI+t6aga
q9G/xfnr5mR8xyrU+nGnS4wAlCQ8CRJRTZeRIoBWknpJOMztj3NRK5RFtX30gLo9Ashp7V39qnBJ
HzXXMrrNhTs3LNI47Hw7nrV/Frsj9qNKNW9KhENuXgU5sqpLNeBrV5z5BsHV44v+pENmNnxKCBV7
WoFr596hOL0lRYzHr4enS/LGqlXaov0Mpqj5IEcZVxYjJFk16R+h2OLT83ISE1o+4GGYFGnhiSw1
KuOKz6kkvVVm3xi0QUupih2XwWnnkJ1t8Vkw/Ce+Ly5V2a56EujIfT8fljUVnjguzXzfpH/aI+aB
09+dne7mM1HT9SYon+yQi/6iz4AL7TYeBZ1lug0dZFv5/RypmqbgwLjvX60gtp2/rc6OcHA93Gfu
E2eFhRM+wSrMBpeMCdqxQgnOmQVqW+W8nbLSAL4/s0srWT/cvll/r6CxMSjWk+ji7LUdulga2gCZ
gO3/bSTW2pM+NWh3Yq+SORp+tn/gIVutw3r/qyQGFDgTTVdk7ea/G/8Cd7SVtJtSZEitDW4eAOb0
pTuk3rOhDC2T61A/LYbpmsK3pCmfKSWv1v5rAfLBhBI+5TuHeDftvLFxAnnAi490dcomheZbiSp2
CUSZGQ2rjrB68bG0stS5+3Gq5eunCHwmVCyzh64jXdjB7/1MfWd2syazCoL2CV/qe2Yak5NtdB5x
a4H9SYUXm4kDlLlMtE+nR0m93XaF46J0Rih8gpqtSsSs9rfWe0JFFonhsSLIwWTwLwGR8IyJwyc5
5exUlSgakNusmE+RW66ixiSOcEiNeLlVrVXm2SbOpuVa9MXMm1iT+wL+FnLSo+7QMay+uCeYp5gN
fLA2NCvvW7AAopzzmoouOrUKkZlPg5H3btIvOJ1Sz+WlfIeKYp6/Elu93A89wRKFpkyGG2zy1zSI
fLMqIk8Mx075H2bB3ecCeWAX47RPhOKNzp3Kqncb+FcLtgSUlrr/n48EZ/H+5XQ5DRv25whwe87i
yxVFsP+hM7WyM0DAGK+FV213MkLDlkAx6NO20jPXE0lPghmNwNRN1XIM8QJT/1WGrSg6AOm+APKj
SqoElIqPy6SYaCoo8t+KR3vfngQYRMuLFXAPR3XrDYzJvCF2k035y0YfP4UV/kifv26JVr+p5YL6
YxyF72LHErY3lQ8D68qPrgsFe8yxWbIPeYyL06fZBC9abVgqHtJzyLJVSpwV39IB9hFuxzgqS+9R
KrG3ppmr/ZBoiYeplAtfbSmJzrdGQTAA4UQFo7R6Zv2zGSukNz02CTeq0ELru/XQYMPTsbX9xrIT
4TN5VZs/8Gvq90cqQ1Xpp6WtOsVusYBKukMqPhYsdxFRDXyWib5Nt0czWi2S6jomT9M8QdGQuIY6
qrTChIGJyMc3lz+urFOFeG3K8FUJDaks0jtHVdP93cvxrVA3P/V4ys1SOhaCmh+fCd8QWOapWxR3
yRbaDRYvPCBK9MxK+QOnkuU+jPXsVypbUfMXq5UqAiz9Iu8ZlnfDiLfA9k1cNtun3S/2mRbxATn7
UL8QsT6CWRZ5wqstCxg6Fe4Oa41fZr1XEt7hZXnAAUktRd/vIBwokfBn6giSENPl8xThAUKSMrFP
3EEZrq2QUEfgrkQkQYm1RaegEqp+2blZHSCyLjUHr7z6RrB7o5bKX/Ky+9fYC3akwQkTL+J/+txl
yHJbgM+4g8/paF+fENT/R5Bvyyh2iPZEY8yePst9gbV8NH/9suiPMfBNBkiu9XjTQUAnvaCs2WjQ
2EQDX/lH3SyerNlWu9nrGIcu6RZ+xfhpCrZ2Il+vG14AJI8Pow5AeFXPib0WteErghSytEdmYEBs
kC7h5sJnaYzcEdvcwJTM2d+rapTp5c1m3x+8qf9behARIBE8ox/hysfTTuylr326koNmojDiMPvR
f9TJ5vQwBAzP6MgpSC0BesXm6danBgpAvW3q+qQ3WWqRLPuS7qtoKiwZXU911ZeQh4mfuzV3K7+8
1Hsh8dTC2sw4MP31cRnagYBt/g24J5hJLYosQgWiz6e0qAla0drg6tKVBH/raAgoFRaC9cGroiLK
9x1dhYiHwwVW7nFBfZwfeecwAlJcxGIU1Iq/X2zmATSpGU49i/rA5zE37W9rDsKkJVviQtK6+MKF
J++mN/OXF9rhsUzKq43+HWzlUEsyFuileqNF4BeKPzz8zt1S5J/nzycHFdjdXBBKHx6hoD1CmBW5
CtaXRU1eK53bdiC3bE2QW7rHbQurqmEPq+mR8gTt6Brp3CGK32FnLOQz99CINs5Bi7wA0K8hScUO
7pv0Ja6Tos0jvCdXb9QTnbrvEn1uTqvXhFzyFhPh5QYBOYF1ZxGVY5r5aV2PrOhP06gZNSbDh9DC
m4H6KboNBiBT6v1RNxX4F45cYBM8MfDTZDGiedQ7y0N1CAfvXQ5TWz1PHszHEEucnjiNdD/N3PjJ
dXdSqZPM9QYtukYkVUDSIndZZd6aj9y6Sv7eFQZ/2IgkfYHUMLJ2hGdxmkmXjUzn69VPG9F86h0s
/q4wUGSl/k3hTz8IWfGYSHeK5gLK2P5LxcwBi8IaGsTDexCqbCylJ6FRQc+JmXt8lHOYYJMnV2N1
aeUm8MzESUGtUGOseN3Bi9kIxKe8QdReMJblr3qDP2ywABKqf2/l8pNi5Zv6Qg6tQMpaccE6zkf7
p814s5DcJr8E91URk8eseIqyUGs4geJPlk5zb15BeaIs+WLwb4WRj5SNvQWe2uJyGwTwBSajM6S8
AFtzHQ5jhxbgYJiNVe1YPZOA4B1dJNEBbGVWTEwXgw5VItl0APUhtL81ibS/pusjFNs5s3BdNtAd
A9zEnkKA64DBOYdfPYtIWpLU3cam0VJVG1YbRHcRsVa8ABtcLSqwQVWpnO5DXIWYrgNHxJdu+g2/
6e9YnUQPAcO9zwt30dD8KgeCcy5Lm2nLk2lHDW87IEYBA74gD186tiA3rKOVKQboDMHBURxzHyZK
X0etJyATLKYJrrGDk+TezS+dUlQnqXNF8AIG7kG7ih3LziAUt7rlwYvsoUZq43YPHqVtjXa7ezQt
qr6uqF407hVcXpjNK3QdSb6kvPBjLcseUl2CkrmmDcY6pG5+X2fsV8xo7aYK7XuwA6EYfn6zTzZj
aT7fbz8ZVFN0vgBg8kr/YL/HxjfPD7N6puV6Klxhns7A5fua21qdlj0BZUxuLbGLdFjsPqn4Ia3l
2CWVsQvcfaeDpuKNZ6lHxiBlSH/A622MPZdCNnRru8xD5plzH1VU3o3BcOCmW91PBEviiqjIf3VV
1DwvspWrkiHcI7kXxegps/ponG1RFTTrUyyrfwYmByIF07PfXqICcp6PdM5E5XPSB11DZC+OIXCD
qP3qE4ScWWEcHA157V0bhiTu+Eo0abbECfYjqoWQMHSR4yAlfXv1EQROHv9MODkf2jGQOkPt64gC
LEILACj0PBPMNuDv2YdC1EnChROMCfyp3sCyxB2pd27ZLtrTWYEbjKd2CVItldSG0cNmeLUtN4Zz
ufVHc0RzRxnY0ZyTB9yUyBdCf0lGXY88aeBTJ9zMGNQ+6ryuY0AI8QsWjmnJ+n1Sk5YVRFMkXkHf
H5qqJKU0yuil0VipsmjAFB7BA2GBcjWYl5eeHL3kwIPHvfrqOr5li8BAI9MzWLe9DXuT9SwpXcjI
Q35u8yvXGgiFNKNsoyhn3XhoA8qhKDrQSGwVZB48aexHUWUmTauI0915lSwY0hya7ioutN1M3y8G
38nTVTuwG1TNftnX6lmE03FG0hXIaYwyFLn2XdGHpdu0dZxrmh6bp4J/VAmAF13T8Elbmr6+cL36
jM+E2GBrEaWNXvxAOuPLn+rlkvfHYq5o18YDDc07lXUQzfXuyIpo8l3jHLcmqpTqTP3ZRNVOZyEY
1XQ9DFB7uJX5/NGV3Dg5F6zf8ji9A/Vq86T3iUONueo5GXQHUUBxHVNeS3iyq/RnbnQFbbKlg+5n
6GXZe7jfnspJDxt4kOMDLiarTCXDZopXRNLXwfKFHJrT9F8egaCHZCnwo48MiwYkRdU9rIhMOucY
tmBMQbNyAIHWt7r5wxyljcTWXf59hJnelBkAcGtilVCR/N0jRMjoi3ZaEGJJMIoiOV6GwU7aP3PZ
dr4qB+6lE1Sjk1Z4vP4CPAjWFvktxoFb4BBQs9st4QG+OZhYobLk94SOOBECyGW/TprlY1fKuBAf
XKPy8K9rIwB0lLzwDG58y/53F6YABZVzcVLqirsp+1P2ME0CXBZ7qYtL2G6ooYDGSTy8GH6j6yag
odZu96JkWFXkbjywVsNkhh/ky0nG+VshMGg/dvQVnI0Yhda8vgLvu/ie1EHI7fE4J72iozCDjPoB
KssAW7a7HS462a4zKbVLxcBTKjSt5pzm+d0MsmJXaUSio9FCkUMyG5fb5ZUn+icWLBIdQGxDxVjK
DOPQGHqyilF8JxferI8P2EYCbYUUJhXQ8igJWcLWKjua8AaCkDCJGv2Q4m65GSvTr/r2sKn7SraO
/BwahJaOrYjzY4mD1In2i5PWTTMSS/sknIhzgzwRvFa7lzJxvC/Xqy7eaAvEOoM6UXb11SgmewlK
EuQusqDqskVjK3gMQX89ZgAkfuhg8AQDuJ11lNFlC8Xcuh810BZC4RITdID4sL7fK6p/RNPf0BRL
qXbByv9UoDuMGjCwU5w0DJshR6BFZjBsSHeqITNmuqwHbFX5dtEKkdSj41XBr87LfMk9ldrRsW2y
PrCuofh+MdPG2G3CdlkYUpeOZV17KyLU+jGQGRCnSi9QErNr1RutqtpTikfQIEF5UAdckoIRgUKD
tMTl+MyDqpd4yDw+pO7+6MLHq1X5JhJOF2a4cGv2IxxotnbH3it6NZ1kFS/hi2mQ8kVgF8fldNSF
mHcUXZMugphvtGxmaVaKrCix24M3w/+VnIHgU2V2FCTGwCsQ/WaBruxDsHtgMExS4XModJrcCMI4
cewdv6u57CImn/H+c4qR00aNSAFAktf0MpmruvoAx7b8+FOAJsSPsjYLTc7IDHbL5rIIcC3xfrmZ
UC3C689fa6RSwqcVfSGBPKhcoWzICP2uMrMMYBnwv7WFTdHttDzU9136EoR5mI/i7G1SO7TYIYQg
T8AyTVZNbOgNT3jQFLC27PwtG3IYjy6OFrHRxXSdV01AuMeg6FAT1md73i0B9R1+Jwf8tEuG7pbG
+qy15xRBooX/IDAELIUuuZNmwCTzAwzbz/tbSaPOLD41J2wOLAQsfdI1DmIl5iHjmSnlMGjhBbck
XhgIpnFvVfwDGXfW7ZjV6EzsDfIKcGtti5w1OT/YVcDqKVt9uxHWZB9pHRegidPmcBPiVdvipOzx
lAHZDSv5EErnXH90eSe7Ejz7yU3gHmYt75nL67f061Nb1zKr4htoHa5e7qQcFZgXhdPMfVcJi0KD
3cDYG7THWuZL4EO8v1MqEECjC8g5jt9amWeAwE/AWf0XS5P5ODJ8m4jSH8Z2U7CM0j3mX79Ix42B
h2/wC5Fa2EwSDucVx6SFTtqk5nOuSs/f67eabKzf+r/tQ5QdkXgE2y7PsiYQ99f9K0yCgo7L50S5
oMfi7dua2KBpvLoAUQ5pGlfDxxAS4wd5tfAKsNHOympiTeJx9fraKGHz2QKXgh8YnPiLteA9+Zvc
BLJEhCuP5IM80u7Tsq3DfYeEx8q1hYZfq4T+CiEbVspiAFGGUqCh9W6+ld+9eVwJa2pa0eJ9SXVW
22+069mkutvdGtl/Im14uYis/gNT0xKmHvEuUb0aBxZlRnO8glLCGG1R5xkKP9L2R2Zdru2+EC7M
9Je7v+luLWtXivVxRZ7IniNcnjXQZmliJIDZcYpg+yP6Wj64HX6c0866RJHqXLNaMIAe/sK7L71L
gyfddhZYfFI782JpMnLrlMfJVYlBvbsrs7LXW/c6SxQctTHbtrz4L3ZrFSWsASqZOW+DdgZP3CTi
qjQ+OpYeLJRuAD0NkiGsE7uFLup+KEsfp1a8RPGx50EtrSBL0gSYuo/YiXQOMCGDWrJBMYdoakBA
D1OEm5ClYy6OTlMJx+/Y4IcNclMffVSSMev22ILIFhrExuEozB6qEw57ZXgGzWJtk12cdX8t+fOh
yCFJB+oVli8coKs6IShjssgompeyj2nowNBEVPRhtR2N0Rp/Qh/GRS/jhJDvNChSU50NT2ki5BHc
PKxglceWEdbA962RdW4bm+2bZZNSGC/iniJ90rD2UUa8Pb4uF5z4USOV4GEZDZc3pcrGCV0BgsMW
u/Hc42LErpmRzgPQ53Q9/gCAhCvWU4J3JQQn4qRwDa0+W5FbtzwFLQGV8+ARyVx9BVyiD+NqP/2o
lnCFWrItH/9JYcD5ysToKHIh5YmtkWXzGeUh/bkuHAIiVjTtNSK7nwUapuDCItiynWsUuec4NCCT
KMCOAS1SsOyBVXWKTBHKQyqG9qfDDkF60arGvgYPi+UND5KhTLlJjGPgzaj4NvmPKazpVVi81GnT
KuV8h910fULGFirOSSeRxwff1hzD4FAvkRP+P9bwVu0IvHzdlLrTjIFsUOe4B63MJyZyFuKsr4XV
NoUu/xuYuH2fd0IqPW4Y0cAq5ndbhT5VYVtEkvlGt5uC/sPVy4/4uU7UWvtxOIGXwN2KLECZNF9p
myL4F2v61qcK7KIGbn7V538039OqO3c23tPqImdVkOQC6IGMVS/mkDU3FrkinwPVmc5TWvmEVOuG
LkZ42CxzGWZVDqTcY/1av7WL3iKt6ceX2iGBigKWJ7EaXEfkRDtrO6XTMR9WOTeL25hJ3T/JWa96
sk2eBf1Boqaw8dq3NP9gV4RQGYIZ+HrZ8BEVhDtZHxK1ykQ5OyXR5X9IloamJHC7IvDq5e5FaELv
RjdEXHs1vyffG4PDVJN3LVRaBW5n4goUbx9VVBK2bACDRg5Q9YW8Fl5BaEBuKgoa0+Z2TkAjC3f3
r2gCrL3mQht9oN3BkhVySykyVeeeKyvtBLWh8KLvJ/88FBxO58BinOAd3PKi7gIcEUSDKI46Ogox
ZLWCPu0pBBNNnYmA5GGoFV8AI8P83IqvvmUSdVdMOZ/G9kYG9Mf+rPGrDafM0ECGHxHM0Aps+AqD
RCLWJauGrv9BM/SL4oM6hxLj6afh3WVWXFzbTFMhuFC1Y3mCEZnWbEyxCwcN3F/Qg1wp56KJrnZF
XGsOsOfsGwxvS1FwlX7dVKROj60SpS4gkSWB9DvHndZSOjiw6jDz/pxtFzSd7g35zFi1P0hZyjjT
sNS2CUpAYbvluKbzCdAu9NWNIPMk5MdVJ9SlgBxnSiThyDDnqf3Tku2QKC7KMJmlJNFQTL/+W0Eb
HgvhkP7EaHs4Kb+Z7fWnwr7i/TZNRS1Hv7U9Wyy3UXxtHcYo8FbJyj0VTPdzNdCXFsbC6KEQUnAs
RwabgX4YfeOeThl2qG80RUBsDuoCbdu7mXydqS6+zqKd/lOF4glqAdMpCV+Vg9k4vAicEUwOUrtM
d/4vh8si5VTM6RGDlxrSAtavcdWSmrsw3+DgvMLeHo+phLd7+YL28qpa0EZC2Ko6EsWIORSxJklU
52oLGgMotxNW43jK8TJoa40Q+WjmWjyTWgpGsB22bqLYGv54HBK3JT5FvZryIlHIvzDazEKKvDiA
Akn4AEAcGR3IkVAkpPvT67bpRv3iGP+Ku+BfNjR9tb5HtkkfVnRxQ+i2wNFTNiAzZKEJVKAVf2vT
RLkIVG8GEx2QT57fjlixKZ+vNgB82xStgrJNDeMB5a8lgrSvDulmuVTYJ/hn/TApqaOkL7VXcdw1
e9jUnaoOI9RazZgsbQct7KU6PvPFXtQ3+6ROH0uOk8bZM2JwRPVYzPJVop5JmDbtCNdqVl9S4WOt
sh+wOrWNScA5Hz0IMJc2D3i3A5gOpco7POr4FoCFc5D271QPSpp4lvwlmIdyWhkJjdoExC9yGMmu
L3opf9TLUAUtPsUBFOfOrHhR0gfFE93ofHpRsCFI+NW4+E9lGoUyCnXEOY2ppm8PkvHtVBzN7u+T
juouWV2yqqmhhSb+aSNO63nyaQg63ByfRE+Be7Xp6v7oEaVIFbwSc+WNsvTaqsnDJVqrWnu5etI2
0WXX5ChzP4iE+8GxvFzR6zhynHylODynB0UtSp7zu8u8/pTx0G5TIt3I68wy1GSpsuXWnI5FgYRo
Q/qPN0m0AJlzU45JutfDl+aAE/obmJNrbEsfwz2JiXcrAGR4ArLHhRr80WEb3HRNjWUQjimWKVTE
8ZO58LtYwsEPuz85OxTJhWl6QS0WluVBEwysVwrCcCjozGEFtlY5/rdN6SsMVEc93gf2N9a7K6OI
0pzg7UtxeLrRQUsaMeYMuU/MvaZE1cUTiAArnurgQKTwoZaicFUGoH/orB2508IAszihKdYccU+9
gxzbtrk0cm0guAUtAWP5bhYj29OQTkcOvrcqg4Q91sgNJXx4Mdwp/bZTUBGsxhIueeRWYIon/pVA
MjEbwrDxrECWBqXdrdRevQUENl/hfMvQnbEIrGvozM26AeJJuqfD5Iwy5c4weJCStBPZvOCTSZFv
xmhXchurOePPWRdGeQGxAGN5tq/tLDc15mZBTnrQDIvVeWAXNJmu0izp7RaTgEc4DDU5+2A3pVHV
cFc0wjGvNdnPEQWHmstMEiAAQDJrk6VWyWZIMvt+jVUg/tuoUoMUfaUKTcr0r0YcF6iZNi+psucu
kpstNqJ20VdqYGrEBO0LrZl6vXTfzZeAdH40+nvUv9hIKvLMuaueWwnbhAq9fmCnVIx/UIMBh0E+
0M6srPnOrcXCeMOO+SFTCbRwhd+HipdPft5Lw+8Qr09ndQaAkkvta3Hsn6CnXkQyEcGvY1RJtgEO
rcUjPMTE91+9A9cZdeOMDLyw4BAmsvYKJscj0XjPG9xlWS6avZvJvoiFTcZpd95r00Mx7Nrozam+
VljWo/w+7mcGkz6D7f1fO9fcWFsyEu7tDjN3sKCjYbmyJSCepzxeFiRvtgFhQ+8s0Y8uK6juBdam
qc22IklYwsEU9W6z91KPpPRncMJGAfJc+tLf2aIj3y5Mx2bAcQg2JRaAQehkEFzYi6AK+lQjkVEX
aXnBbWV5V7w28rPedRtmp8hLpxr5f1qCjduUAE2rChs0enwYC22FDPyU6YYegyxZZb1tHQDJzvG4
98U3xXfOAGpvaUtLRAxntefxBH7LHGySArJU+8v2M15T7QVflbc7yufhpuDDLFrNMEADuDX8ptS8
cZtl+BVdXSJtxUmhTI1SBfH5hbXEs9hxuaqD2lntxz6nI/ER99DB6WEjhXPhCrx9xyiPIud2TYRZ
d4CS+h9rITGRQfAaS//O9tkQjd65DOFVVRadObygo03eaYxGMw3/yVECXr2GvSeOreu1Kf32dMew
g6cW62ZbWojsTeU7xRI1azxHes8LsvmFRVz5sTScG4a/91SkFBCROOd0U7F1tAoTA3u0tDGA2y+h
N/7VFlWBIBaRLpXpE2lZo9Hq4WN7rb57vkfJc3WQCzV8YvSaZFWOZAd3AEBQ1YKs0+XOv84NuW5e
qx03FeZVOsX9WkHZ6LZfnVC5t142y5M3/gEcOpT7XNQeSNC8J5ncCEizhUr+vzovEdxWmhe4N/zY
y2n4FKz+CqYXuEZ/bTNQhfnoSdRcYxPd+jEUKmP1NDx2nu1OsKIer5UrdHLbIC1iXun+9gyfqz18
7EKUWSEqhMmQOgYQ7aiLqYSAPZG5AnsXwepIx6jm6DPDIaXVD24CXq5U/WmJHpIIsRImmLPMngbA
2jugf2CmDVmbKErcNqZm7ufXgpEMaUal0CrOvtjJw8SkVJQ6kpUC0Hzc+MlJrTA3ZOiRkD/0Vy+Z
NfBdG+/U/TVqm72F+8DKaRAAak6Ba3Yt8M9yyDVcr8x2xnjuaKs1b6ZA7RngTBFgK/sPBKLCBA79
GulAvqacefw0B8nlfL6FY8Djap9Dy4VODxMTV4a9D0BxDbNywFu7PYE+WApwDXTA9UcobGcpIubb
UPVsx+NChcCMdAjbeZO5gtOYNrVa7aXZTHP/x9Nu0VK1LZMhXBO2h/AaCvGP7eZJVBy16hOrfJR0
n6eqHx09VyhIid+L50QQe2OCl3NGv7W/qG5smmDGl5VEe6kJZdFZ4kbtdHekpyHqMRwdM4HjES1W
RrxD8sqI/jZve6Kjmfb9xyc01pb51cGaI77EFQlM37TvPv+hWnI6v9s4J0HwUr+4ZoA249EdRv3C
JZEc8iYiplF8ZKIkNQXGXgl4LjTZXCmpzYoJI5E87Z/X4gLSzoqPWDgGG18b6w8SxW7U/2gSct7w
YFSavNmqzanhkMQVpFw/CmOy05Z9jRsQCEdEk9b1G9TFEJo+SBKZa9M1V2BXAwBP3h9Dv6hXwG0P
BPylQ+a7pJuoYiLRQiL46Ts8Mzbglg99q9da/Bf+jyDWYA5r9tZW0SGrh1RCk+xhq5rXjpn2GNkF
4tzk3mKPmvubO1W/LFbmS7C5I6pOHaEJltUEKGkyErKDn/zf1tnkbh4n29Xt51v6SFm7NCcn23tI
2cwoZBuBV70OHlnIjRqqtQAcXW8n2aSetOLXo8W7GVFxF8o805AsNfwP9G63uDtMPVo3EZF7K0go
mt7S0soXGk60ksrTwVtfpJS0cWlV//OV0QlgheVnF12EhPV6dDYqHH3ybJJ0SS1R81522KV+u9PX
cJXaV4l+njNOpICoa5mrzVmdmzRySd1PHEiUFCPPbJDKSkpKzfWq8mHd/3AEaPqYpRWl4sWajSe8
bJKzQnIXJCYthDer3PU7Dsv3JReg8mbOeKYP+fBJc7I7mjM2tc4Um6+q0HCn2SdmsB0W81+5wmg1
VuXx2pep+lMTJ0yMwAiviz4iXTJzmeaY6OwHeP2ifujpQK2p7+OboVw2xv1nDChi5g8mwdBCXCzU
BvpOMaosIHLojNptD8rI3Qz7c30FxuAHibTkivui3wRxRcgZwLEreRnxsQKAiq3FYyr+2pgdaeti
KvhswrI9zb5WlxPBg6jqD73au/wKMuko3zCSY6z2UOFrTWzHbLVis/NBdkbMqqfi2RuTJ547ikm/
lBYAWesr0W3JyBk2ne1CnNwoVPYhnz20cWA/dfBfEiq7ef5AHk3VLgWsp+jByB/iqgCLHyFxjeRt
NXpBDF+rzw9LQL4Y7Ks7QSpF52rb+UKaUHACPtpL/JtTC+lZ3FpN3DVVKmSKNx69ENrlnguxLXjc
VsUMVzrQzSEIhY34Xl6MYagzrvVJyC8UqpwSWu4D5QT6IgN3/nmJ1h7I31xzR2j62Mf+nTsX/aQh
Wlz0ZPEEnmmssosvPCbFBh7Ogrry3dxsf7TgHXJNL1LA6SyZZZVTrTojVfHxLVX1/Sahdf9lHBk7
TsKeCDNwsdPxOdoUkSZkFQC+IFoy4sjDGAwosSXJrAVuKPeC3LZqk+mhpijyMoDIxluiw3AZXljw
k0jzs5TxWJNjQxX3vM++/EK73a9+Hx0qrTo4eYeZ8HX6i3xvmZnxpLphG7B30N/Ds6lazqvejucv
bQgkRjDIJ+c+1HFBxolboY1l5EM/zn1nK92SSD/DEQGvH+Q/hCrLDuFHe+VYCGAIgAHmzVBMIRee
oYexLlVaKFvBZFDyYc0GWSTzvYisMWxXOZHXlLTnEpwasg9keT993F3OUi58yf9C3QCKpj31LCCi
jRQhSg5YGygYchANabPDJV2JsWtoAAuJZHuHStAbLrfRrtzVPlUaia4rN+fmdxqeKeoMyqThdbTz
sanD24NnrW8TyJdjeIfG+Db1Dt0oRYLY9oJ/ausLomXQlJlajZeKH7K4bdaUdSX6+5g0ArXwc+XL
x/ldTPKbJssPXEWcGmt8WnrbcufD1UGr1xNpb+eW+5tv2gLmmMk2zQjzw86oLhRgKz72hlsH06jl
o8IokG8hBP9KHL9+Aw7hENyF/ldDYATDL6E50gw5kqjsBuCr4A5aiS0ZXFz2R8FFJ/Sy+A1ucrEY
GwjPlkaFCob0nMF6R4Rs3Qv4lHwqy8puBWh9YTwwqWv5l7nc45NW0+uQFR74fsqCRPRkYOhjqoLi
ak1qkaR4fSWVIFr45XpQ5mUWvzpnY3PSjv09VtKCy8Rz/WR7bcv/JUkgbS/lYYKC3xA/JTbqlBP3
hDEmUqxiVsxuKTQop6n+LTt4SuV4qjInyQv9Z1zkPPFIa4zwtnKB4D7gtaNK74T/t7j5agaRlAAr
q+kh40JY14cGs8FVyqjcIV/CFwhm3Fbe1R+jxVuRle/WK0c9ZCfhfEK6Gx3RiyB5P09XV1Ohx8tU
QDIpNWLxMI1Oqc1PENT/GnMLFjX2ejkMPziDRk5lE7lK7kNgrV6WDmR+YL7EVfVZWc3KnZCpj4Nk
/he9ahQRdyyudK1I7GnMvjp2npVNZWWTy+cs3ieYIsbOWGAjMxNSKZMzlUqSC6fDiBsNj7TpZXsY
pRutGGd/oR4P1NYarO4QBTAnEZBtYuDdlKrwpw1Lnb47Vw42DRf2JLzpFWCrGrxV+KRGSvPkuDEj
cam3T+ztqv5I9oVJeNAmR2Fn7RjpiWcqUPnVIT05QsXpalqEVaWyapRMBgdDJ806Nr6WO7YlDxJ1
t+oumPh+xegSUydItwT47BPNwd/9PXZ5ynP9d3HZ7rZsdq4qhFoqyz5MHlSew9AgiZAvFP2Q1xZH
2sF9mWZw9nW+ML6yarUS0ilei4w/2kEjIu+2YGPTYs9jpfCRQ3NztqN30UWvz1SPdsyKPI7GPV4s
zJvLkSSVvAJrYXguT6xavXac5qJOFYDn5KvtJC2uYwIL8Nib8w14CtOM+ZIW7+dq9mG1nUp0mEcT
71Y4uYG5IhDQU8wWFdGEHTYEI+B4ygCCke5JCLiOR9+dZofAPkguuEWrFlqeczR0nrSfMVngdG88
bGtNQyt+VpQEfwcTL+TNjvHB/gDUfXqQ8fPKCptWQvt3NjqIrmE3G8bNSKEWaifEMhJnoRgtnWat
LpqMUm7Xy0/yNXBC2b5Fza3pX1qGnpobFzZW1LiSf1YxETl9dkhRY0qnIiYw8h4oIRLH5TEnHSkR
NqP37S+gvO2s/Iu/2+/f7nS0KvaCuypgpHhv3TVvD0ch6I+DoJwRFszJlK+k+fO5l5TgIV5HiZZD
3j1X2+3I/8FTUMk+MNi6Ti9bz0csQ+6dn5YuUvGAXhZARKLLXGXJnVhUSvB0+16C64Ys2vLFcAFC
sXyQXbNe34aqE0e2eVfPc2bRwzoZPehkNOJzoej2lbMyvDzMD+iMi3wRPUiXmvU121SCKGzzlKag
W9gh2IRwI6TOJGTqm4txPuJ9GZH48/0YeMA3RZ5jukDBofQ3SW02Rhwz6JZaBjFHzFiXyG7EewSQ
1iLZR3onTV7hneV+TiwU/sTejG9YCF9ZrlLU/C4/tIVUlmCdA3cwN7pg3sVM1cRW8XTqPLQOEkjk
N0MuZF8CReE85Dle5HikkkpKoMrfa/3kEmSztjxgjgDS1ZKyP2Zjf1WyTo0Ui5HTeM2FpX3WmKal
WWbFuTrsvUAxGXZ+DLSo+ADlD9Vq6sKcTyWQAQNt3KA8FNkflsQrCaLbxDH9vV7AKEUy/p3kyKeI
BzP8k36WxgsaBdExyFO1nixWHULjC3iuL1CzH1fmGZ72nklMmeZG/xnBp65Geu++2YlA2qix60Ez
zCbyrPt3qniwMSNcE00gIoSrl9Sf6qqCc6cOgOz+dXBpSp222W1xaoFtg1vEMZ4XZLA5xSOyfkAs
8+4YAGOmGC4lIkutZVOcYmL82XyxFyT9PGmZzbhhnK3hIAaEOTtAczZImJqh7O6t58xZnxVtioad
5BiiJJclPYU9hZWLxfAUH1asgRkEiIvTBqBwavecqTJbWym7Mt29P7BnLIC99VoFdH6L3uQS5eOf
Dooev5A/jdpE3Gi+DLs8NT3kfXve4ILFL169gXIPexEuGWFd+iKeaRRQ0BZszbexiWhF0w/ET9Kt
Tg6d0I3YgblP24+607EHOyoXfUFE/rU40HYmUDwXu1QeBsE4ThLaDuoZS/vqoWGsb0OboioiydJN
Cpq1b0ZiCM+wwm0EdNn6E3DXUYYX0lo17O++oABwPUwEbh9u3fPGiz9zUfgemjlaX9Rwy+TwUNRR
lfDIupRgvIqiXu9Kg0Vv0bC8nK6XLyoR8P73qHdUdKYRhtuc+0eUR3dwMBRIHr7dfZReu7Ntc1xv
Plkxdz4UVaj/66YUrrg7PqsgZXlx66giFXU6VCFZijL4vTuvmSVkDvUHyWwM2ms0GdQDR8zC3aTS
HMfrEmNYzpkR5FAzX+Rg7y9czlxJ689GiRPRX4MOtaxC7QjLF+rlaO7qNDgd/y4iTA5IV1BAXZ0u
quj9OWQJyYnJ8L6z6vpXuXBJAGol1H79IT29PhVS7Cn6AaIYef43qq7YlRiLMDY2gluiZ4Kx3Jai
XLG/gFLOO0YUmB7+2X71WVsdWIQhM1Z76kHTjIbSCSe25j24U5/8wBTmXJgbt1gIbewPV8ZOQcmh
/y+437yvucDDp0nqnDzQKtrQeUdrGc3N3p7GN7W2ds9Qym+Iwa7+c4CS1QyfuX1DPbUmbdLxYEuO
nqBoyXrtCsoov5XqC61JBEZLAtoO+n1AlQCg1K6VoeOgUVwGV92HogVMPpGz611jbhiaOjgdoAI1
vKlVbyvu/yHET5yvrX/Gj9Y1lqEboPm12U5VkQBSF57W8pfdNQ46xMW9av9WH+h1RbgpPNdr9TEd
DRnlok3RXEjf3LIbF19qia4M1HCY1nKtMa/KNl5WtXQtTtOAWYlD76ZFDDJbKBgZD6FyREn0DXEX
PNC8vgvqa2vSrsZjcXf0IfgeibNDwSuum7tpApjmPJhbT1CsuZLOQmt/kmHKYEtqj5S2h/R1UJIr
yL7fMyx6+BRymupwZkK0cifd5uwtPbwyL9wKAZztjeIZHWJuOoyc1H01h1GC1khx/H5B5O94wqPu
o+f9XA6JlFPT9rs5Mwu+nMmEWBlyKkMUKfU78CD6hEwM69TkRCfGnsRcleZRkYs4qNFyct6EjeFz
aUPuxrGPYgwfAdDDZap2AiUbSXjyM9QP/QVo9DU9i+aHZk4jPQmMhqyU1Np18Du67DVb8mWS6T5Z
EcYwuWTMadzDoArG1uM+yj5LnuM7qIop4a6eFuIZ6gioq7I18r2IvSGG9uc59yNVaHzKriZeuUbH
QnhmKtmTP8lxvEuYhSzLjJiiW7pYeJr1NpYT5uEQcl5YaND9OzdWIyYj3fKBvUbSGOfNr82pjQtZ
3SF+p/0kTumUFRycny34oEArtM3U3pzZYMDySspo/6yjVyTQ7fn0+nn8BT7kKQ13S2CMNuyQ6Mch
BC3YVOu5wXtyv2RLOVtvOc+Ny4yVvgHLwaB/mgrMp5pWHLXNa46u9JuQyoYbvBNACAerLPu0yNfN
S+sw8gCsupy21f4JkQf3xqjUHL9IOevFAvE+dZsONcxGgk9LMY/Lgo11p0cEDoq2skX949zrBPd1
lmoCTv0PxVyLpy81yJlI7rqe6W8NnSXNGZ+QynQV/bB7EPk+IQpWrQyR3fAQmEomOTBy+Hgs+VVB
gezUSYPLt6kgnUDH5WW/Sa1JoNrFNc7rWS+dtUOcnOQJAF34FOCTLR6dFrHZAjXZ5ADa7eaMSX+l
G5BT2I2BSi/leTI/Q3Hilg+WnZPPv0KCwrDVjCtLpKY8PFpFuiMd6fOCj4vJMMtIudgIu2vwX5lh
cBOKVLeig7NlNnmof4IQHTHQVqr5Wm6L/b4RxM/6e7RHCOxwYAnHgAb+pP4B9R+o95bXwMXH6yQ9
OIBwMpGFA4Beoptdv6rrdjKtLo2iuq1blm94YyAUsR28qcyZD6yE+5eEOu7bk6ogvBBTgsKvrJcA
XIM3abtIpVkY+xHzVUCLpHaHMkxvI8gXojUnJunfoI0d0aLS7+9OrfnDCAb50ckrJ5djj1nyghI6
CWRivWV511szDGoHK7zRjRoLaytw/QZwxZ4FNG46nrUhH7XkxFA4a74QdV/r6eDncs2lWTSHxF7F
KJJS9rMXmijolD66ei9ie/VyG1VLTuaJl9Hv0IGmy93UDqEwuhiUM4hWNMQ3E9+GzTJdSH6EvGKf
Qc0QkEUK0+sQPU2noBRqScel+Fz3xaYPiXw58gHYmxFCOxOXw9XIJGRb0l6ePUsy0zGziYh5SJbd
neNRZkN5sfYu7sL86NqfmNhtzGJ8O8KjH4TpOV3PLV3TOwjHOAn+hskStYpWGbX4CneiKbCx0BMx
aRHUFClc2+6QIeOoMY9d2q+lQHWvBSx9ivtZe/UbtBLVM31JiIJOQ3eAgbIa5oM4oM4X5K6lT0D6
RgUndYLUV/tYcmPCCqTPXjrCFD2f4VzcrwQIidx1G0q5nAzWPgk3jbR53gcVLUlLj6oDBLSY+YTc
ICTAh4b+yTPLwV6nQkiTUyIkiMeMEt/A+ORMbK/BHozN7T9qpeO9Crc9lLrB2kp/+6jLYSx/aRPx
QKBjA8MvpejXJHFPI7G20bJ8k1uAcwRWnHE8OCt0pIzfJeKAEmlghOotv5RA7YUSrT4LoVXOtktS
2Tdpehx/UfGQef5CJXnhsC5pQVGEU20kxqWUKCdPpP+1Vd/u/V+5p/MMweVb4+3fcN1c3UTx93eq
TQ3TiJpL0EgMgh5Ybj6Z02cFtQA1iYZkUKkuWvV4037RWv/6bQyPqE2syV1mHsh+fFKp4EKlvmnm
XKy2/FuKpmriWaA9xrRNkgQljxXFV4EfBXbMdPwlk8N4cQdwz2Bvijs3NlIKY0ZZfwCc6k3agIkj
IvCVVmeWlRPHtd8ImcoIb0dRe+MRa/2go6dwoQatQYoV2u5ud1vIIMl9xg1xT8EEiNnOXv94MSNJ
XhEHdT3GMJfgwt87xgAODiSXPzhdQLThkwmsL2zeAa/eRHHwabKMlQrqBcfzm60v3fD5liC53FBH
RSOwSC+NDTPFiwsVnY5Ls9wmuHOzKGq2FyBlm32SUCJVfoyvr89FLHyPZbYLBpkyRlarZN6lmrhh
BQ5hS8+vaTTMBfjuLxlYdgKni9CVCzWQaXB6rNPiP9Zgqo+WORpdOt25+veoC+5cdW2uRBrzJxVL
ljKQLVPsctsfmZ6c1RGL2jOyalRhtN2ZeWlQkykWukyj5sMmV/9LyMBy/AKxfFNyCkpm+PabKIT2
n4hALAyKy9XD9lTtVFPNYkxT7H/UfImZWrRm9cWLB+8gKTW+NU78jpavhP9IRxGbN+/54KcnxQuK
7DeKyTzRiRV98y/IFQppSYRnXarke31lSar7d3ry+NOcWZvNLLWzqbipU6asK+7wBRNnvO3n8jVc
rj5l3Ry2XrhW9nN7uOEXZ/ITkJRbaF/Wr1XdHBCi1ZcJ/NrfTOylnS61IOT+tXJ61DyHgvMj1ZR9
TO2mN8LySAOG/Z3CnyXwEuR26PujaZH8IaSNAH4IA3FDB3NA5jNkBcC0+H+r1FR9y0s0Y+4809hW
klk/NObvYMrkn6TQknUohtFOf+YUGVPqN0+Wn3yyvfWbabgDAz+uURTQCT+7d4DcmNy6Kl8VhViw
NRK9P6AR6sP6PJD0OXfTnmtPwdejIngXb9sq1R2IAoadDLKISL6xcjvqeQz+Qj+Xi729bd8oWvJL
aNfhHCuHWPoj6/nB1NCVnkP/Mg4EqnIDgyZq2V+pzhH4PUX2Kij2dvTxBUHXyWLW76E3OVPWBtWg
k4iiag7LlAlfMlz6ZpdfBCT5wBBVZQCY61c3IDVDXa+AGhisB827JWzXZqcajnZpNRaSLHBkso3l
93f4O6nML32TwddeUW7BvFWCPN7QzNjpUYFVqkzDIk4Eoh/iSoz97aVkWboq+qFt+F/yl9vnaLkc
FcAH240dbkvMyBGFS7D2pvJyKfGSG1rkfaoujjcWNz0va3/9JQyv9yCzBGk/oklwMQb/o3ox6qNx
jbRKrT/6LC8JJoin4pj7b9VtD9eIJrJffFiPAS9jK+2WR5aEWr1kteKAhn3R/xBZFxsy+zulRnfB
yYrK0n4ZEaRP2pvBxgiBkZ0QynfsVUppYJKnlDErZHv/drQtRCZbnhL+CLzHBEunJjKN+bUKLf5B
OvCAoQIoELi75vB3FoxQqqEYlmryswy8b7V3DHFABw0kjID+Aatdq70wqGqVikNtnTglQ1tG0+1v
PWBsFZQ1DcduYsTjcrDwUtgTJFLEq6ShX0RyXM7ksXRWgpqFNmqaYC8UoLQ5gJAtW/Xn5PdmxH9M
c3Acp2pYgh12JiJF8f67fDbiAoEtl5j0HAowmW8S25h6ZU1PCz81ghjKKJaUochDgZp2scQw9Nvu
S0r1qyKUdznJmmWmyDRrz8/QKyPzt3eBA6Edrf4ZbKrSsNIw6CCAscRmi+m1Mi005khw0vYeRPk3
XTmgTP49ZL0Rt9lxNFzqBjvsx4GdZIRuXeNGaH4H86e+Z7t9Iql7f93TwLBphln7aDgR1kBMUhdG
dl43sDpxydMi+fhPNY+yqpSCssqCGEtmAvcDsUu56ssuAENu3mtbiUmVfZNNMjDezLOys+HYwYZw
VSfUgyFqvazZaP7uvh8v5Lz42Uyl4+AqQI3q2p4aG/6ExUCarE0/5ioacJKwqBCmm5wSo2jlr0Xx
mRML7yNaD4g8sY5TmZvruxW+cVA94S7+AHf7QV0ClXiwMDipwjSzJT9gJavMmEJ5DhV6nRHlJGPQ
1Evwxav8KndMfNzdRPJAAVQmsh8yJAlYHzHQB0Wb1fyUgeSZ7l3grbg+xiKuyotoPXnYLqx4VybI
o3hHxCJKp9ODFOh/QSeiBO2C471cf4oFfm/BVhy9GwqlEWickv5jch9WPYP7GQj3b50HKz/ycLsN
HJsF+xO7pclbhOiajMZjfnftKKugwwVFBwahkj0gwYDypvOYv4/afveV76mbNxQyZVkWBGXYa0q2
2fZksSVJ/EdGKMo9j0GarwI4bGSHGG8UDJOQu+ufUIVLU33VfhzgjbhZMagxiF3JNE3TO49Wcrxa
YslgXBVvgY+KyPvy0HvAWfCPQv3AHyeIWRTel2D+WRXVlyC6L3zsOOikR0G+GH4CXguXfcFT40kg
XuLvQ/mnwdDxVTvrMAXoWnY4MySAAbhd/aiW8OagkaL4CrID6uP6Dsomg9lEpH5VJgW6R03AR76c
720utpPzkGF5O4JiINvlDezZRtJ1QLPa23bhqsgD+6/5/56oVQWi+y9WGFrCA+RM390Uc2kaf2gC
MJumZZ0I+ToKtjbldbdgkBk30jqYZjN2Q6/LvoY3M3+4JO4dGmusl68zVg/SGWe5nU43z0a+h/hc
HIXzglY23RHp2DjSmfqymoRQjiiO/nO/1DmRy7ElB+HKnBPZ2f0xGXVzfZMNwsWzcFqMmBzzQITQ
06xQMT3a/Q37WEkV3n5gV6+frpVxi6vCzRtDwcTvVOOUz3gKckLJhMtwjguUHE7Hdj2bKVWGiov/
s+QsWA/tQfcR6zCqHIqAuTdK8iYczfUxEUkRSYV/sYtpYbK2qBn/nPnMDEsiHTgnCkuhCu0qBFWY
BW4a2OK+t6ENkFItm+aQWVH0JeCMsUGCni5bkf14+LmfOcfBYo+ysicMR+Mv3nim+KF/YPZi4k2J
y33EG+UOlb+2VBqArSYoBfXchxjHfZszWITpTLN+9eq+dX2VPYlUX7pgHDc4B6EVXRDzLoymrGcT
HVdnNmbyr8krCS/ArfKJIayUmqvmux92yTc3wjxwUeRTC20BI6bssK0mWeS3tGHqZdDgJ2qPwJiT
rRmndQgnMKNkRstS8w+IpXfQq4U5gGHa6YlrCDiUk0jNxj7l49bruQnov/9TMBVNo7Gsw7RfXtxz
JH82XWRFY0L+rTSi5KhYWtJCsijVf5KegcC2cEK998bAxa315zfzyY9B6KOmWoIODcZe9jkJKkhd
B5TFoIC90pGrRRZxrmzQCLXQgABXNLzTBzUTZrIVQW/Tws9bmYSGG0koDsiJKov0bvc+yuNe1hI8
Chq256LMDinpQHKWg3NBt/Moc+43qRrqA260DOEo+m3BcmMVXUAnHuBsJ5+ADmBZuQT2cRPcf0AQ
u9o3OskXfrD+C/n1SVdseLX0O7Sy07sVMpiCM2K2re7Rz6ovsF4QkEY8qd/GHa3AEoQROyoCe0cE
VUR5dp90LCwXXckVtL/Pbj/Bxqhbayx97CHEe6K2Ul5Edz6kjSaIlpTzmic2WE5CDGugzJtqFGSk
AFwkGV0vXIANfmXl/9ftcpSQrQY3nuL0kuHPdj4PF1NTU5+1wvQ/qwFvOb7OSunguOeCg+DKbfw/
2wSQpm2/Uunkt1d//wy9Mz27rMqkkRfbcU1pwp3XVdmhVkNgJYjyTD2pJ1MCRH2gmnoG0m2ceuLs
LDbjIkZMMItF4Bng6/2G3yjwngsegQCVfzkrThKG+EeafsibQWwj1ZnDFwVPhcwckpk+vjfhLZnb
eUmtZ4qIl1+UZJ0v/65A39ZtPfQFzG5DN0a+JQvJRdozQFL8t+TgjB8B/XiZ+VppX9M7M5dEvqMn
4rNzYrHc0japHS1v36B7WODT8wE+DhPmFAK6OwNq8WS6MiFVhTNyLcSkBjsfP5pnSyFcvZXRJBV8
3EV8SkYFBUo2REVmJSlfyK+WHeVEbLfy3oJE+h6ajWqrwVf/YWMt3c7hIAijbK660fAZpFJvNnV7
bLCPM4b+fzoq6iWziZMsEenmV/XHAg8xjn9gXx7j8k9Rs2XQXp/6KxwhTT/5MfochmBMEsjsVjmC
xICf37mIBigzafItaNMqP4fT3VLQ9CZRleqphHCNI1AKcuuABoNsCxVvl1cNuQElpdEGczwh9pwS
dK44SI+XM2OgCOSI36ljQ3LV5vjrqGsiMsxcC9EJAW45LXWsi+2iARi6/h1iWmcb+oZspMF8nJjM
dNbO4xpSrYMoEMN7rVB5z+JMiQ5k5SsQkV773Xuu6SZLTaYe9X70LWtgZsMcEcWs65PUCnkOprsv
lL87cNDNnoGiopvr8Wbfqf2aOXjv2Sji/Ct7YSt7aoTeFH+wEjFN+htJgjr7SyorH+/1derErEza
5v32Fuzyutd/RC0K724RC1J8/raDv+9WYuRNUAflnD79sOQOMASx5bAm9W6MV+nL2IcxwP08mX4o
6zVYRcFcbvK/DYUNoKfYOq+IpZSwU+cavpmE9by+A6K93DllI7TXoklBGZKKnA08ZtqiiX6SA9PM
ZXAgcgfa9dB0Ox4Rr0sd4G0cfGPsV4FOmAO9B86lZQg2ioY6v8p6OhHvpaaRZIKIjkU8LcyxUq5X
oQfXJ+UNWYAzvYFl24V2UuaKc1Pip6fvASZ1pv3+otByBuDA0xKAcC4YPbqPTwJ+uTXXBSxCQLl+
R2hQg8eWzChgFGsBkcrFc/VdmOS5omRh7hbr3fzMCsQmeOdbodU64wTkKXIwiUNXiYteSwoJ+ofa
X1Dl9E+4pGRMvmKA6jf/1fjrDAR6mC169B3KVjqfoB3x5UyvXYPOGFyVZoPNrjzoklrflPFsYX2D
FvwjPNCmF88t2gxi1Ehj3R+L6bw4urw1A97BTSDip+FeyedMvtXjG5BoJma2qCYGPM9zSaHpPIMc
T+7cp1N/mioL84NCCjoC9IPQZREyRq0W0kvMoI0LbLYLTU80viMXSpJJgFqn8ySqFLbWSk9yjNVZ
1HDOsbZqRfpSfn46Iwq5jEEApfUkW9k5dK15zsCjEu5WbtdWGpYk5wllCLR2nx3qG7VgaPv9JpDC
Y6Xl+4hKyo2Ww8plawaKXvX0X8s5TXrm3yKqfLwR4LP8lLVow4/9XfjRiJIhQt/MMhPKcQnhCotf
aP5Xuj5ZEJk5Vs7Ma/Nw8nUcKq6f76f2cVt8gOysMaGATS6Fi44TghHf6tV6Iqw5rt/LozSOzZ9G
1YKUtgZP3LwcHXCL0GFC184qJFGeYECmQe3EnWr1KNg+R8u+mL0nMFYJ+Tua2tvu++NfLh9l4UlZ
s1s6ouomfH/PCj5SO5fK9JLO5HS4hX1zB8XsdkWkN+jG9mYLy2LfYkpP6WqDzUuTsllH9btTNdPn
ZhDxG1VEStEJLmYCS417jqMtF1Ot7NkTuF2M1ABzdVFjWOwGq5bG8M+UaIYSJosg3iK47zGaZVFt
E6N5maBo0KmevSmeXRsZ5/uROp8T6bO6LAezmcHtbPb5EMs7+XvWtdGR8YKLvtuxz5y8hMuzjmox
UbwCVM2vXUjBZn5T97Rnqyya8v/DtBVIF7JM6w7UBHdlOfdfnupeJI12g/+gHSG5yEaGUwN3uHTz
qGIy94Oan8OptPKVntb+FJrpJ/O4K6Wox2WSIGop1YWMoKV1YS0+brzK+KYv5gQ8pXaO3P0cPSZV
8oDPNQPbR6cf0/jdCr90yMP1kGENs8evUavj1phs9Kg1sPmJDRaJ69Y1MyhApu1zLhGuj1NF9qRd
TVapL6uDkckvFUGik1wxXQLTGGO/DaMATuYANtpoFlfSPKKc7n6t+I7jxH7TVr9r0e/wWCyysMO4
vCK0EVuQRbSUTYWZHvlG5blgbMLTp29BlBoDmALOD/lTJ3fTo0xVdFckFA5Xm6Zn90uv/wkQRBnM
Bd4xUIEON9Qf6t3tiDb0nc8O5h8co4m1w/MkNp1R7vJgsm92FDM2tfEcI3ctVGAYGsFxDyttRuV0
bNK+cIFasqhihf2ycz2lT5xD9Qnn0p0yQXp7K3fMxg8lCeGYrgrJ5mzea1LLlEQEh6iJjh+otHur
XXNmaPpNoB6LtyW+XtgpvthNeFO9+n+R4fTBJvnUTYyW4sc6vCR6aAyQT/QkfEb5yzEDNXQ++km9
PtWkgHp7+exgWxWFzYnFanoGEWUatFhJhWgC1VBjSEeclwIdevof5YCsMKmoMQjxwzlsBsfWAyIn
nHXklEBR9LknNPrfH4CkJrzc8vEzNW7t5xdeF7LaCbbaBMl9alXRxPGezjDUGQ3HW3JXQspvVDVm
Kk5Jqi6a52PiVH3SiO6wfvE4frypdSHqIjtYdlWJiHWawZWpFYTtBZ3O1vlsWtz+TwdouYcgY+TZ
cvGr+QTOb1GFCt3CiA80TSSfqJNM32+FRBvXaSoyozIwKnOuJDbFdpTqkVwJ/wknlyrE04PWTHQU
SSTZ3C4O4d375eSrSyFrK4yuSIGjCmu4auUksMkdVfBmfAPSl4viLrzRTLAu0/J/yakaMyF4CBR/
UZfF18Dsk1k8sr0r2kxbnFwaRvdyDcGyi6l3Q8EO0JSBsbwfI3nzBYx7SzLusoRKbOx+5B4qLUEw
C3RoVaBIqrtcSxkxKR9M1J5sGnCgUZNpvzrd8cbrzGohm2xHpos26uYZi7Pz0tlm/fJWdghTeKVH
FUCtrcmLau0wbQJRRDu9yl66ai61beEBDb0mh6aYFn2UScBhVGXqfCJkBfcu9e8guUAyJcl7XJOa
kOJVbrqa9ZUP2SMspvpPye84S2xt1thKIMf+An9NpF3gwe2Boza1ZbERuVCuuuGA5xNScz9vm/Di
KqGnlPQeG6IRmMA2GE8YcUBgdrk4SzmEm8RXA+2tcl3EFJP9rFOZz68gfRk7ESJ5KeimCl14bKOJ
NV3sKrEmUl3JLJvLaC3pyrl3eNmMiYgZHOa7A/Njx5GWH+/z0LjYYI1MvPJ6GEQeaVJ0szfIjzrs
Eq3fCwjaO9eWoqVSe04mk1g0nH3LS9bXzDoT7M+oZKvZd1A/1DD+dSoq0ZXFgYUR7nBUljO2IONt
m7+ilF1ZXmOHK1DAEaAs2khKjy8hQ64LBw0suuJB2bK1qrEPelj2+l3oBSGzvKmP9+xTys+Ja9Z1
hREx1MSCzVEOszQ/TZJOFyxhR4kI+CAsG45sPb3cdjpJeh55nc2p4FTYvuB0knQjsdwb8Oo7qzla
nhcpS++COy3COVkhyAAMJBaUQH182KXQ850fdyZKm9D4fkxcLB7ls35z0xTN8AC5nkF+aoy1cJcM
HksqyOBUUeRtEvPkx/n5PX6tO7itLWE/s/agh5/CnzYYkGlc6ODvYG0mWVce8L3/l5/zvNruYxI3
rfkPPpJBknIMcngEaMlLf8o6gRZ6MUeRQzR8vx4VUKnZNuH3QFxawihjN/SFE5MrjdCuJxAqyDmw
ApEmEqiYFZthxGMWZ9SL7FR8WWJ/DHEfovmx5obmnUQ+1rivbqkoyuxDSKVDAmRa2XjkEeITE2nR
AGM4Cevp5pYpvuSkFG8uySx0aYXw36hxU8j4rsNgzt0mqXuoZlBxFm0Fgo3M1iLCUhjQ7aNJay0/
qDTlulocWOAc8dtj9LKKW5iJX+Ux6/99SkMyOczxu+p6LQJfRY8S0YN7pSLgYH8eOteNyivlAM+R
VOOEP2+8tt574SdOd9UL5gHaN1tBpPW5VKR+8fE7P2qA8RrMqsekWruiqXlH9mA0PCpmbTjbEGVx
2xLLRXPNrzR/6L9rKrV+ZJbb8RKiNVyslShNKiFXo6OGdk88UXRkl4mOxW29sX9ipnLjYXSMNlIn
3iAOOJDVknRnLQOSjB3vjA+Mq+8hSZm5Tp6Hb+y25Pdn4rUAaebKojthEvPIaoSJ4bEIvWdzZTm5
z6Vf5utHMjzunKQ1w6omM4ITj1kXTF9r75nHHp6xAgoEOHHjMMMlUnCET+KY5joIpu8EjXHHab11
CFLG/Z4DbOZzg0HOi6h8SwfbBkq2Z7/JGOKr4H+pdX8U0hnhtJ+S5oyYXJGNu6yFL84ENzWNQkKe
YJeqeJRXrZxL280sWlIXwMfWdW3fPhOrIwIt/pts2+XfayUFn7Fbjh99iHSsQ7uZjScMrhiWa/79
fgRCPR31VuMQii2HA2LPB56f7Wvaumh/Dn0v3Huutxnyls4mGP27C1Ca7kz9yE00C2zFlLkBdse7
WuUA6Dl9xB4Nwj2hAiPIiMK3oPtCpF7ZB2bo7y8NbMP9z9oa1LaMzwu3L90jlGguNVYj66p90qbw
Koh25htx1L3UtHwJUI97nYRN9QH+RLMiLx//CNuIyD41Wox0WL3Ss5/1UytL4edzXT7jRAuNQd6O
Ij9ufYAEfeJ09fsgl4jSWGwjN3WOUz0uupHhnJl0w4JpKNk9Ejp0yZDHgt+wSkWbcsYoFgj/L9jk
SZ9sY/wNm9yjINvOuSgAZ76V5IYNgOnXttfypFwqlxoIYJm0QrXZjyvovdCk8qt5yVwLRFhzF+R0
Td8Q779uEBfYo7qXGiDAcEt+KkT0jWSDquJYwRa9ME+xth20hg24e10PBFiiWu1xewPZB/feBGOr
+qODGoxKyxhAaajoEwYsf5BP9O3E+Ja7CEIwo3UiZw/lYROqazsyObhaHxaxzCJRz8hgrD6XVjYa
gveItZYLg9+dqDSAacWDVCRNDGHaAJc6daMzpI7OzP1dqXELA+eks/nd4KE2bBKL06xn7iW6N2c8
BIE6IB0EY70Fa+9lIPSXNMQ0ZOUxCtx4IjATe/eAbypluYTdIit+1a+PqobKqwWqc703/SsjASSV
M2UJkP2fuLMF7pJ7U60fxE8Tm9zNtJHOsGJj/8TjjcfNqeTYOEY1TrpUByIrjSVSdhEjWkruLZLu
eDZN9ydLorAsQIEjHO/gDJGF+sDGcV3xKbqCHwHKUek8Zz1OfWW7XFyR8junQzRtHrOUltjFxXPO
qZP1uQDfGbyXrhUm8LCWz4Pew6eCt91bxRTBvl+8MY9LR7ExNay0yubwPmkBJjLN4p2DKBKJf8sh
QSctoOjJYqhF3kgyJQbdbxbbXGbiPWsLgtv1WxSrGx+AcoouPOl7+Z2ap+glwvMf05KARxwD3/Vw
swSK2BjjhV4hNGZTBUhDOr9vWf6Qddic8+2A6hG+UCAPC+TYCbSi1i4HYJH0olI50pHMsPUCSh76
Ir1SbPmqsFAmuzP3FdGYeGmRz7R5W0idpRAWh3+QdXp082VB8SphYM5IdZlyjjEAs8Z2Thiv0735
nfBTxPExaqHCPQOY13FpH17jXDKlprREl5okQXae+Je0Hqg8qYOE0bIPBZuHQ9TFTCqhLtHVfihf
7RTaDQZh9HlNLMyk+Vkum+YL+CwSgaAazRarLHVBwSkecPefi/FD7cSFAIXXqrp/WjIFIc71cJTP
PuxURm5AaEuJU3pajjO6siFyexYjeDtQQRrezHGlLzf4+z5+/zVCntUNcBkUcQFuvmvGdXjpAAAu
gELc3Ybu9S2OJ0BuBj8nhmrH1AoDlY5NsqBMqx2fhA6Bfecn9ZmCphW1iNXMSxBdd3zw9RifNBfd
FHyzCPwW99fi6OlEE/jq4ABpFFuHKWgbyzQQhlm9AAuW3NpuAK9pMoLYngGhg1AWMUWA2+nPQpsv
lv1C5g1dRuqv9vJpcWEhhMffGGK8oW2DrqiFhD6PlVI0owsQaOsUUkCcrYHPtOD+PIGQfw4io3wX
76ypRwPbg7HdHzAfZ2wPNPz5zOqobha+pR/xszrFFh1n+mHT7Yhzy7OACMmBcbREtVxZBCoUbGyW
GiX9GUgWBDNvSwwB7kQVkmFrG8RS7E+LqcTnziePQaMXZH12dtQ982xecQgzEGXbdu+lK/v6/MX0
lLA2Kn+k7S2wBmNHuLEOcny+AhxgRwvthZ1Qe2ueswCVxrXeunvFPa2HMyz2qVLogElkSHNT9CE+
2qpIXKY2RLJ7getbpE3wh1rBghPOjx+X16Uvh3gwuCOxlCnEs1skyZMO70uenmpAf4JQxfAYZGX8
u+Wvst/eof0yJ161hognSifsfLIypco2THq+JeG2MOVFmXZq/MIhISc+fX7//H99xGu+6OMTOct2
b0QYu3hqTGDlAvPIdTVU6YsRZJhnrIOxvL7JCojXVB8xPuvSHYWlsUiGBLoj18KHtubRc/e++Cmi
4LG9CLbjLPky+PUn2Bx+Ah+e0mRAAzzhqr2YT0hjqwmoEEnuyvSH/dZh8DIhbfPlTneBRufDKiIw
h3rV16q0jH4IZNa+/45Zfeq5RN4HSlevboCw9sgfwnKped11NHKGhjnfrxhjduz4CNbmYFoTewMO
bVFqQ8E8bNY1GWBQVT+vLSHJTcSX0LTJOVYY6kKD6+IYw6i0TOY+m/KrOuu89BrlGjfdEYZwPuCu
PMcphDPZr7CuaxLece1FQ1HVMwJpuFiJAEXafnwQu8ByP0BMI4P9B+nfLTX7KdQOTpaHMDj2jn0G
HSU2bso8CnBx/9rA95tfP275VJMdbyhSOxqd4boVJ96WGd/7djGbKVGU5A1JIFsITxa+01ADcf0B
EduEDzgQHip5vi6OtlU+MZxsEg/5DDdqu7lHLY70rGbH9t1BuBHUxw1LyibNT158cK+AragBlMd2
k7/atg8Wrj/ERygsMAXG7sibMC7c7YVg+75A0G1AWamHj1BX69vlXqXWj8yi+W9p4L4tHBK3Kqkq
Bh+SGHhY0W06DmdzOEH61KqTUe+qJ/TjksZ3ImgoI+/SEm/vuHCSairUvivmKWVo59hxhIltqAeM
carYExwIMxwJuZouS2E6/J2G1N17qILwSueg529PKxZp5Gc3Mm7kWmm1sNQHC42ELCvljUqcDKJW
2cE365TDvfHpmZN56BVVNebLaPjkLRy/kASddjcFtVjglwPvGdZMUfJIjse0q5VLtJVAbD0MMB10
dxjAz6GFXgMYCnRWAG6Z6SZNSqD81mY6yloq0SVhwEWfh299TUfLMrD7tsMSXokJQitSTKmXGSZp
x5a9yBkYrqwHdzyuI6a8WZRLYqwx6w+jmGCOhZz2zQDrJwlWbbaJSIRvXQRDfQLPLjpcRkCeAPVS
Jeo1UmGQ2yi0q4jTfmDMEy+Lhv+sSmnYGj1nqlB8TNp89FrKYf5U63EghVG0vzrQ1UbmOLlddxmY
Y5ZHPcOHSF0dLZz/+DkNEP86EUxocEQDnWZUugySpbI0On4QSQVLXp4uhKbeeji+gMfvy/qvS491
RcjvAMLhpJTzbBTWMU28dPa++7cHlpLkMq3Vt02Ka4qdttwOn+/YLbNEf3Qm1KjB126bv7/YOKvZ
tYVXUSP7QVroJKuwfjo0K+SNRWo5VJOkPIx7YRijSmp1qD3SzpSC+0vWjQ/SGJvMLkx5cloJy+i1
B9GKGvoCyWYJx/iloj+Olq5Fo0JyglxGuvJ5ttw6f2wy/fGrKJI4eiFZVGvd/KLPb9GRhCFrRXN5
6UxOzki5kxNcdnKTZS1PwxwaUFIk4t0IcHaqLJiqPKJV+TtttagmbItc4CGhpzWd06ewaBt6YNGa
2B9CS3kkY9OWvhmsmpDlHiXdinFCzuPsfX+pn9oaRn9sqek2b5N3dk3b/J3aErJOfzJX/CTgfl3T
zd7eD6yt/VUZCvKPxANeMKuhyCXzsuazwKplM7lv5U8Y/BkKx2ilNuO0TwznOxg7HDAgAWvYnGjz
jaflrCzIuWuzoIla1AL43WxQwNPKkz5+RPpJ66wi6GANv5rveV8hA5R06jGJh34kzISJ9lVWk9bv
oRzcqkUM1lSr3hIpFpg5XErOiQ06Ad4+NUbIKmwkNXIxoCvjQhS43zizd4x7QvOwKxXgvVB/FYjy
w5xEFThml1JZ5EQhva8zW8VBVfnOxpeJbQXPoDY5osK455fVnWIPqtWeGxrax1XFZLVdnuagF6FD
H7KktbZR0+JGZ4N5u0uDjWiRibVqoZFMy0o7oItb2p12EfGbP+7OjXov24C+gXb3nF39IJTw3rc1
H5u9e4zk2jzM7kT1C2ucjelsTfV6/mYU3NRQS0KQnaCnCLAZcUY/ptNz6pWsmeunlRvSBRJuelEd
mGjCxzMqKGjMD0Omjsb27knw9QA6ldnQhu6QpuyBKWVgNxpUiKoJvjSr2ksgT3dA4QT/i9FNuUKW
QFrs1XaUFckq3OK+brQVHUVtQZqjsjQ5CNJ3h1U+1GMKS4yPLCsFUH0xFR43URobfUGZpZIloyAr
KHyy9S2JPRgWHYnIoQKLBMbdHgkvugg8aKnJf8zqBGdVFItZL3JQ9svv18jga220FDReBXjDqot/
JW8CpQTdZjJzfyjjJfPjNa55ptHXKAOTqZdH5lYQMc4lYNAfsZn7aRlHLrHM5y1oar4sEMa7MbL0
YvymYApTKmVRMl2NHkw/MFxk6SGBVB/XGVChda1qYhSH0kj2zK/u3tIvES5gJwOCmsg7Q+pQ8sB0
SLTRd4rqXS3/6EIuEEpZd3TlfgJuYSIdVWkcxPyhd3zOFNTitK5Sv104cI8HlOmNK2LDCLdArn0x
UgToMXTlIiFoab4qola9Or5lgu3oOMKA0Vvd+tm2mitNjo2dw+M9dyZRSxkhgBEZYocvfws6mBMh
r5B96sjxDJOBzCOUN75VE2rwF45aAuOno15Ln/KL3i+k3M20KxrCMNb+e8KIPmtD7Yz24V7Zgt/4
/OUWBAW+/wjvY5/XtOpXO9NNkrNf4QjcVOWTUWGLhGZ89o+o7RdBf5VEis0Pe8fUBH8E+tPHghj6
7JUjS5f8qMlCi1D95PL3FOw6QBdeprS2RySx7ICEpKAIp1qMONijA9AtsgGX9rI21GRhQtVy5WJL
xMApPwoHCXg8B0MKbSO/uUT9aA8hoqJEC8451V7eTp7Xpz/mQkSbe7BgPTM78evoo/vTD/qsk73H
jEz10wNKaedN6/BXVPdFCENMGIiYjCWE3tqno+4zdGfOHFaHRd6c2jluMRX3U0gJ3kvba6zqQf4T
VmAWCtzwoHfzjn8nzoJAwwaof33vKkdTRi5Igj57SWnlMIiQUzZF7OoYoukC2H7H/sJ/sltKRa94
Tt7kp+7DVPns/s6HT0ASs61ZdQF45GOTvXnV4WWKoC42e0O1u9Hz5n3P4Kk3EghLmirInoQySaLs
LAo/4vQXpBjwgV39L/H7ui10m0yzDnEO1oNF6+7CGQAPjYJSDl7LTmkOfZn/Ox4QQsl/VRVfddzl
b+5gn6JYvEIFg+jDodRUYH1zc7HMoAmzho3934AwHFlhaLWSncoKQ/pASb0zxNyzPUi/vy9x9yvB
H4LH/l/AbwxrAG7vgugOQlhc8Qpcx5hvjcx50slQZjGltj9EnQRiQFytFZo92z1iiFgZufsv/2OF
Lpc5SYdTYgwAOujEdnBM4SwTRphKDsjPj0nbftHD+GIdcDOggMIyDmFZtRFRlpr3pXlRHGefPEjJ
KVq2GgGw8OrvSpTMK7vqDkc/e3SvZAYBFlg0K3RXXzTctocQucROdt9iSI4M9fJqGoDla0qpZt2w
C9wEHzkiHaKDzwGUsUcucVW3R7e6v936wq7HgsMCZnEhSHtcsh72XtuSnsLr2fqhF5MjqnPTheji
whjZ6Ri5oATAtNbKuhU+flkW7uNTPc8d7NuYW2I6pmPdF3kcjkZqKvp9NpaZM2uTk56F2+7WY+TM
ta8RmMTeZFIm8VfYDhu6ydclA2ep3S7PwTm8/9kLBhPnv4gpbp4McwTR3di0ovBLoZhkiGvc4bgZ
pwUwIMF4PMlDzdb9FjbdOQEYYFiMlxyFqdnZgBqTZ1rV8z9qkwn+gTZw0AIIfg8jq8izxxuUyseQ
4WS5Q5waLJNOtB6TU0aC8v4W2VV6T+xDQoZOaz2PqTUQtDtMnuhA5jEobtYVoHsj1q2faHAIpVyX
Ku6s0qwqJJTJwJtvyy3vFPzbsp19cuPDTBDcE0APTYDh00PqtGeGTb5mk5GDKc2zIRR90ja322lC
fhREflj0fzSTI5xBXdwCEDrnXNVJW33N+Cbpe4ljwKTQ9rQSzTlz6Ib2oqh6A2Pv3/4l0bVpW0zn
mkD9Apo5ymvM250a7YxHbgaE7MF1YXsnWmixqzlKDvwcIrAXHymkW5H7ESvLiuLuOqZLHL4mqjlA
ZB2NtDgdRaLY4d+25cwdkLmMrDb3GAYtT/uBx47JBauDfWN/EQKYTllilbrMCroEa1OYehkxXRP4
fFgZc+zqibwZqaD1PnAZH+Al526TVFZQriVVS3CQsh0HctMlD/uFl11iLCEnvm/0mhYGA74No8ZO
+JQm8EnaN9sUfpbolcGtjEvz5KOmFre5VufnabHcf3M1nboEgrvLjTOJ4FSo8y5ZbQv2zWxD4rL2
yk0Q6J+FrenjpARE32KHOXq2jLmKFSTrw1AkDPQgnChZujfa4Iayq50Qm9qig++DP+eLW5l0Im9J
OEgwAxoKlLjCfhEYl6cCjByt+icrKcO+DzlmOt7fwI3FnSJdG5RNgQyyMEXZezScJXmMZqPKQPDZ
uSgpmzlv9hKg4QAYDC99sd3T234SAnoEeKLnkbEQwtBW+jjJnhu6EUsa8Eqcd3J4jSegC2O/tsqD
LFfMnSslVjIMHpGNc6phfPginbTRFMke9C7wNvlP4Pni+KlAI5zgxsJleKHHtm3SQ+xv+NqDQ7yF
0M5YLuToq74u1KvYr2Jh1kBUO4cCka9/3+yqqICPElnIvtfZo0ou1dVmy4k73VQunSwds8EMGHve
WmqkcW87qnNkAopy+bKiJwtLmQvsg9uYcl/0Tr7RtdyzGsU7dICd5H0kXZPVeZumWIderImRT7Ky
lezp1PkjhN+5YaoS4YXO8duHKxK9aIUU00KkOVX94hlqBAQYLNdLUpUZNrtRJxDjRMfyTiBxx2KX
gVjjxmqlpZAKwsa3V35HHHlSW+hm+CzLd1vCngxlu6T6uhvoazEwZXonfL6jP+t7cutyl0hvF1iX
ZFpy+2/It1FuyFX4vwiKSKDnd9cL3jahevO1i+O0xqNSUjRE91lF5aO7BVFLZfj85mDvs2CdEyV4
M6TEO1Xe4XdB0AzdWT+KDyPZ7Rs+q8ahJT74NGWc58orL1jw8dA01fJb1rTw+X4QBrd1+pmfNg3e
/x1KjuhJczzOHtAS52Jv/rneD3K/abWo6u2ZtsFrTs4m6e6Zg05U05hoSQNJgkMPsPNpharDzxr2
L5l4+avTJmabOyonpQrNburP2Grbt7NgMAtJfIqtyXCJFqlIdMAoVoF5hCc1WaZn70EKqvwC07ms
GX07rHf8rEnSeTl5cDwrlLC35u7E3XT8VSj70GbpEkfQf2sYz/YO+XybCKpxYuijEnmppE3z2boL
iwopRdz3yY/PGfcV1nMPFx2mqir+b/jgc21IO7ffiJY42NStk9oF/uiuJgWA8jPmVAJLfCO2wzax
6+zMyE16h9LCGwHcXHfy+pxOsI5erJJZVs3JlCxiJzDUkf2F/ltExLuzTVwqnRVuat9Xd7l0+XYw
skY5yr87pejGM+gnxEJu4d6Inkvk4CMr2fG8BB8b8Q3gglkiv9424AIUq+a1dtjXZ0TEZ3RmuXLr
YbjG9yDO9WiwsloBQNvAV35HX6Wlr0GNNzlA3Fl8PpfP0Pf88XRFMttEe6A0YR2biad8E3B/IW+b
pKnv9tOKywW0CfjPC10IM1RhFMCaaEqKlepd/mJzqtTxPIiMAnrt5MVxy767B2sKl1YbLISv6keD
yeaL+BQmPXjWroEgl97qfhqSHPfrEtEUGai9eCACqakoy9EoYRoCvip6jAUTZ6g446G4aYlAO5gA
+tez6E6SRcPG17kJWkUVxX64G0dWBUkYtRkXtsrXMqIpPcpCO3akKStGrMs+aDkkgMaLWMcL0xMv
t7Ttrpp9MyNq+2YtqJ2iv543EyXXeQo8fVGK4WbmlfExogh9q8lFnLmkGp2LuyBoV9gbR3c/sWrq
7hdnbTCxq1UTXPk4Dbtg8cxa7yjmyLF2RkXCz/8zv70r/dK+Vl8ufEH2pjdyLVWZOWWsigg2UYnf
MQvRDTZZlt5YeEx3BCbN1IbK3n5Y6AALwDXrivBvnlNza+z5Ex48ZNbczo4CH0nF9N8tDNmBvu2a
9aiU+VbzggMWVix1+ODTt2rQN4XIyPcm1qSm9q5OH71AMAA7OlmXkRYsRs3VKweoL3YTFgvFPhGd
DDoea/gkHHCSASQf/91MjO+Oy4JibMESO1zijhQD2szyb4E4+gLutMZggiG3K4f9OY0aqm0rEMJb
e35WStVfykzZqpJikUhXI4lwttGYLNptm7Ijwg0ZyVAaQtIjuXhTOflL4Pll2cd7OORnahiaRqa6
cPwtVEEgSpAaR+5LanKINu+YyUSRcwCZT0iNUedPRes3TjF1LqhDyyl/yTdLA/qzzLjAgG0s8WWE
nZcQkULMeC3BkRCJhWTtnyhYfkwkd54UMYl0ehJFDEoBRTDIFYahJ/QDk+ysf0A1pmnzYGHpg7MD
EUEXug0rU1dbdPuFl3vqO1mmU7NwifWLXI44embLyydaLuSgqAueZEgcLv6W+2i+bkqt34Kjj8IT
ACujmxkqOwdJLSvcVxNHjSUhqYFRDreUkXt+Fwyj55DmFCKuz+00e9mfb4xCIHAjVMfsGTJge1AL
2SmelpE0YAyBFCNzWQSmoI3x0SJc9Z9B5c4ony4ahb+rxKGTp9jlw2Qg2T5gpgar49mTtpoz7j9R
wi4Xm31+qZtMB2Sd27lST7vWI6vk9S8yJSVPRRWH1ldJ8P0yMkRgG+CDbUdSnGgnlSoI9z8gVYsv
dLddU5bv0y3iYkgTln6Fed6AHY+w/oK7h7Ki/DRrQE/R7UW6iFGNY0W0Gkb43Ig5ANn9daqlCyLO
5M+OykDVJf5S0qgpCslBoGjc89Cs1mS92irQYR6yFQ/o0B6b1lI7Dj9ot2fSQbvsV9UwFnfmvpXy
gwLlRULkIdqgkArdMd6WpPiaz4vjg3hK/XwKfCtjGNlslVRHveYLkfA1rZzMtApn5r41Nt3m9Klw
OmjtCLeGuJYG8zoBMFwUOZn3CTOOC4n3GWIkFD/VeQ8P9ANUHB3QqMSKZ03nTBnJ6e8UZ974mpPb
S3n9ej35OO297FZhm9QPBwfi8YdR7NK0Jf2WmZHAmj41imf9JYB2Gi5OSjwVMAbP4xaahymZhGEn
+ADg5xG1etQdTT4PfYV0x/ebdKpyzieHdCxEgmLNAkdQ/htDeSF2BWy2c9qVGBt5so8plAlRI+6Z
6z5mqtPFpE/z0P7P6VY9C/Huptw28Ba9tC7DpHldnXW2gAVRRwqePpj911V+Q0CQ0I5wolNvyQTZ
byRDYSBCwXCzbOI3/s1YGbiO9jhqkuje5/kVqe9o1MPbVx3i9bSrE/PFqQco24FeUjL9mqJU/B8y
t44IQR2fc7QqXKFYCfPWPJN9GpcYYtHfhPv5sXifjva8bzYZ68eNeZ1g1aI0taXP3Q45WCxQJfOw
PDlmqvIKXpgpXL5FDj2Bp1fVZAEzfaPlBymGEoTA08JeV3G+FsA89Fjy/8hvKmcAFhuElv7GSRIR
3pz81FuBgx+94rkoGQa1Hn0HI13eGL7PeFmjiGTyR2jzgS3XeOlgYtx1APbNfTAg4d06Wgj4suRl
a5zmsIP9Q9EhWk5NReZUEkU9dLCxpPevueYmnOsiynjrjxkKIZB4KkuHeX9hyB6WWIrFg9UnVsmy
aEWI5XP8g345PU3BLidEHCFu0yMK7GBRMtApwbKvdASn23RwRCc1yHBdqiYFsHB4xIPvNKAJ1VyG
CvfZXyZx+xLlUtrGOSus2RCs9AHM0qYbvLhDvi5J+URMXJrpXYOdEa2b8NWGnuNYJ3SDXnpWL5o+
MfRV8RToWtA53BxyquRwut2JqRQN/R71A+8U4rq0CbTpQj/aoWuVjngRyatFuWYtOlK38m8UqY1j
q6i5NpVpll6fpUoK8s3XpyEVX/y5RxT0vUcC8zZlQPyZjTZeVZHBFtg1vVdVZxYNekUCcCNJcc6D
iXe5MlRElk+1w0h/g4O42S7J2uG1/A3tEvrAE8tGOrT7IgFONk+OUWshV1YpArvmmq0PwvoDWdmC
mJL+tsT3G/mcHdXePwvMprTeTU0DZsm1/d2jbn1iMrOgWXQDJUDgcN4F3dBGcgLq0iTLdjtSS18c
Vm1AxMBmk06vUn7kJVtW0coc4LinPWFomAgJlgz3Mc3eiM/+M8P7iZxkTFDlYMKRYsOriFRmhAEq
axP+t57A3xIsXFgpLJ12OWra6LaSzKV98zRxVEXBzZWp4T554DuSH4APOAWOQpc9zQlOioNWLrbO
xvA27SP+Vc8fxwBrCfK3IXAjjrGqYUPqBFm+GD7IB2L0DFupd3JpGY17okipqOQY34d/Ijta7ko0
l8IqjtPO3Z+CF//PMEtB/EEoBLefJzUj3/pd+H3uZVfnHkF4w7XHph6xhWCSEQbkPMDEoASUQAvW
nL81c4uAVDrQhxrQA+x4PYVi8NaOUvmGgSr/ZrbL95N1HPwwFlaPHoQoI0YVWqyyzdWt7jSwbS5L
ED7+DRDEDHtGlWMrKNzS6eGVdsLRW+PgQC0H08nAz0w99FGYStKWUvqjXGv5x+XdCkxdlFbYl0sM
4I1IU5ISUnER6NuCE3l9+r3VTaJ9bMJv08pj5ncTKkP28Me7XJOR/Xk5cLvTZ7N1mONvLd5u0VZB
wTQAIrFlMxEuqKQ3AZnyW8sIxd/9wYUYApK7iyyITAG/TxCLmKx8MOwrSt8gaAG0BxAHb+KU8DY/
5kAMAd8PUlz5JgMSpewo3+/uqGHAoy/M6Sd4qvd7Lvv0IVxUdOIoSKGFTqBhnb+fmMg6fHmqdifG
G1HsNS/n+763BowBzUyz6IgfryC8Dma4YZCVd+5N71x2khpXKRvmEmAqHJiifs0U+JnAIuhy3jBi
I083ge+TZsCzInV25VAMiLBWwWrKmTb7YkN29COkLETC6a8EGrVNVsAqmXW5iCjAalLHzLc0Twtj
/klEAaVAfce8S2wrfmEdUThxgZmB3uyq1gSx3VwDkdivJodm0H1rrZVlhDrI45kZJmeGAGjJ2F9F
jgWw+xGLPg8DNPr7FTffMIsyVLXLTbtTRZ8xDjlOTdydROfHdO1TQ9kgds0FB4CNNR5wMWE/v8mP
mFEC8v3EhboXq2zQZXR4UniwmhK28ujHi5+dc9F/kYYaFbnSUMw2gDwLd1tf3H38+FAgidcTZq9+
XvgsZ3wGhbVT74rXpOLHRY9+wyAYL/75J1AnXApgqFqRfwpKuH8Zj0jxeqlqeqog+F8FcrBmVrgA
2pUdL3/9yhv7lefwXRH6YsVYx96FpCCAj0rAC8HJWsjTqOV4xRFMK1IOlBaU46VbFAPpGBg1SznF
j2okKaWMNlhCjMa4tfAUDbqf49ybIfhFFBr2+tns44NICqo+WN1+hRR/W0YOi/hSIWdAXauWtIxT
3EE0vvdqlG1O2YOyPtUeH5nwvYOn1CM6fcVqYMPeBy8luQRKm7NL+c6JGuWuzf7Ydij4JlA6syTc
je9cNH3+g6GDOFa54ReYCsFO0GbA6FxzAuR8gscUH0IfrbHDkdrhhQU57AEBAHBnEmIapNb2+6rF
0FfFY8ymue1ktojvF1dC3HlMnEf2t3T3PdnEKntPX79CN+yi9/uH9xH2uVyG2VjvVI33KDD0rF+5
/iYSnAXb7v5IDIQkRxO40r2Vw/0Hn8yN0GuXB6Lgd6mmBB/pvgCVTaRNewU8pAadZZqJ1g3KROot
ix4m/7U2Yv8+L7ZOx5BuElnCf/e6a1J9PqWg2FVgKpTnElRoC3snoNfk7cKL/TWG3cwZ5VGITy9j
7Ya0LiSmT/vj5gA89T+L9pr/AX6kDQ5g9CDoJsQjkP7/atHwGTGeYivYbWJXHR4+9n4H8eYpJb+X
gmpLzodp6SoPTKEeZATybtlTKscCqvnOUSmYraDs4/KHyZCUwuKwR1ll/Z6/hU8PNemlHimjWC7w
X+VIUy+tWA8sCgNIQZPf8G99FdqS1fhpFJifhNXHDzkNaXanhPwdPoy7jEZ2hxzEOVdB3MLzdi2Q
fjLtSIjv6XAOXIrrvU2QYbbEqwOKND/vFZFbgSpJcNG0QFe2Ij7EQK5XS0lgJKyrvETX/f6/Ilqt
7qNJJ0+TO6vc+HgHXlL+0Vv28T+0nyUjtXVrdP90Bmhue60w18N656j+Ed5/SM4hX6diHsEhzB/h
D+WB2SPAAPFInSML+LTI3l3m3H3demQIQbPstqd8s/wi90Hyhafp/s2nnZknf7F+oJd+UYhnE34z
fGd+SA1a4fI0AduEkZpSIEdjdliMmh6Cr8WCPpFddKZQ9gRCMyh4IERG9VdIUGbZIjsXzho5bSA3
O+tYNbNFy6NJ0MUhK0VgwY1jZHfmrhmgAMVoPqdJbpceM/JJc3nlEs0bU8nwiJYxo0OxgYVKST3B
ig3rbFNqLITLXXSZKxOMMJIhoQijStPXFkX2JEeJ8R1wa8p6n+NFVXBqezH8qawHWXgYHuzunCv+
OJQi1zbo5yoD0Md2OQOKL5bWS7Mf0fe/feL3jqzg75QoMNP6Y5YPHCSK9oULqQ1txOAHx0iwsja8
u4npFiR5938Uz0gy9JiTNVS7HFiEzLrBacPr6b0DQPqtKQnY6TJDgF2seZZ4jfRfhJyh9cS8IFz4
tX/ewmXwgyNaPEjkM8zGB4gMWZQXUY9dr219BPWL+IC8CzzF236BazdyL6LE0q6Odqk0ljc+jg+h
vW+W+ZODaEIPD5ZyMDlsH9RkdeBGv+Q74ONZ+/4d3+9WdKYuttvRBNjysHHgNbZQ7xEthjaoACaQ
X0hJv25tnSqzeEl6+qAR0q9wx8Wu0BuxKWiXc6SXor1PLYVIOluh0K62JwU7XBeMaogQzLGQ27Sj
BgJaBmPRWnFSdBMmEv3fr7Lawam6eVm7sBGpZfRCY4C6s9TKdA/HSemAjvwlKseUE8O9GICDFqSq
Xn9Ul0nx8zNHgG0MlyuyziPlBkquv7jT8ZXGnSvAGCFV8mpbg+0DnANMbRnTYKS2l4IJ50hl6wNo
eBtBQUN1nSvuYIrxEnjv9J0WyOJTQDMYH4n++Hb7cKqTSBCZgvOsPILUXr2GD+5bLywKxixGAKcI
lznpr5qtOJBNSZeoJQSdE6N+dMkrfrG4+WNDhPImP6XMIAac3N77O7MSLf/8AvIqk91GlR0PXlwm
ehqcicmsOw3UHsQOrkTAHaTSDLTIARN63MCz5SrmRjB+L8tN5XEMyFdtbKT05X1uaP8E1w/ygt6k
65T6e0AdEz43EbGLbEWajDUEUqsbSsDDrz2beiLCXcuGjPrv3GUQX4+JTM9suAZ1QxuxThrh9kmd
3tRfrcCLgkV1rFbNQWs6tsLvZ85rPfMRqwQZ4tRDEewmp2biz+YIHxGNtBr5bJUwa6Bhm5KI9QI2
TPSQvimiedI1WA3Ill90eqbWqqAGRWPSK0sskOBZYgbQjyRwlTD9roafoiiwiD8Fu+bP9X72fhOR
DveTumJGqXj8CKXR7TuNVban3Z+XcopbfpJhHmTKzTr5N/d4s9JxnaRN9OfzoSjXfWC4SLoIxiPS
zA6efKXVET729fUy6pXXeGHTojfqURcKoFOne4LgXou0woIFAvZ6Yh0vjYYpvU7F/h9qalr1YWL3
pq+m8mpML3+U6Xepk/HRs7QIdnDCembsoaMyo7YiuF7rDXS0CUJ88wHwlGA8Csq3VQS3LT1MMhaM
nDNKIpcP/AwxhWQ68KFkZ1AkYstyZ1fWp7gQjSAt/DNdfR/o3brZpx2w/lB3KC2melU1W2HOc5/M
wDYzwq7/Tqa/D98izL1dtTfuOwxrpG6gIqA2nynAAA2IjK1bexrExDPs4Qc3KR7K0D9AdQE1knKZ
YupD+54ZnmGp1Xd3ypHEtbA+WkfmtiOhsS9Wl4pxlLiV+/Byoy6m+Gmx95l+gv/W12tQtmsBk4ij
BozWuFL+9Y307Q0vRKNOkMDAlwQIzFFN/P2U07nF3qH8S4mgp0lktFjWpCw0oL0VyhiqNDhXl8w6
O50u5DaiNU6ZqQ0E+EFBTGgG6tLBf/VmHqnLZEfs3DWoUzJlvcwfFwkAbProZgaevr3PHl+TFwsY
RvaD1So2naYSCro4Ye9j4sct13c3HoNhd1fJbg/uBZBdeHM/aH66J4kaycEhGKPUd0vHkwPsFn7z
Xz0f2eGMZL5s/I8j7r8P1XuXtZFxQrwa8BQrdUSOU/laF9bwP0QU9lAuAMdSqVx7+dIDcAvWO08l
hs2Vp5EKoeKfBNx9SUZ8pkx9//WNi5Rbnr4SN8f3Y0kFtqXUrOWii7l13on/T6B7KraqNx7BuLc6
cYArzrSxHr0N0eI6qomho5VYYeu2NGzNRn7g95vZMRpCb9eGlLKrzwjJ6EgvzbB+/R8KENWtGa6X
1BwqpIslpRhkIzKAGclQaAD3L/ZGD0p666x6nnwqFCj5ALVhi748rRiR5rwh1eKM68eODEE+yXlL
ubX2tWmNAJ3WS8k0lx9B7GGlKa+Fc+awCvjXgMHchwdjT5E5LwDZvBI1DMKsctHSEzoblerm0fXx
Tnjy1FJX2oNczBMiXB39eFTQ3mAaJScODbFOf/xwCLZDjPNT/yKCuRD+tRx4YWXb39gY/wCSucq7
5fw/72brm3BKFRWgKtns8xEOL8v7zePsbpIVM2qcW10H0KPFAR0KVykW5Jd+OsyIfwzK2+oT5pe0
KGOUNfOuLkGcVmH4KT3BR6jBkL1yj10rBN6g/ClbOfum+hGX6/hyoo9LiOq+bOUljVvzFRVrK3Ys
CBjYobs/7gqTayRx++bRiIkshRwKt5+RNRYFdLMmIxY21jVm0+DPqmCC1yahKzvH++tymD2dExRO
NjPXnnkGpJii4PoHgiF56NCRjil6jm0/Tw8YnLYVHGkQ80MJHT2z4rkP64kwF/VbbNbskLh94rt8
nC/BUKovC0rykIIpCZf4A/4HP4OPC/Li2TTQqeNEujd1t+bXjB55shoNvPst5Yz/gbC1m0WvfQKU
nifWuDRVj2kSHdWGeoWZ9GujtA7kG6uzTWFg/FHxvybVXLP7EDJoJfcPI08qOC9qW0CpQvz59tgL
0evfgG8XdySSflq0LiiDGSckAElagcH0KsexYZ3PpfYWb3w8+uu3hcUFs3o4iUBSm4jZolaXe1+1
+Q11OXBkH9iDPftlHdoArKYboJmAwBa5v18yMw/ecH9YeDA+dXnSQhs2MBFdfqTJ4K+6jhfCj2XK
pmLslvKhysmmOSYhj1FTBmyZP2awiY0C8P4D+6hAIGrpW3lEW5oWkUeuwrY+B7sPkXHMovC6f883
IgbGHzrwYy1fKf3JP1aGnbB+8Lj0rGEctmETYNGOkPrYRt4ddb0sBlhgqoQzsvWtY6twqaPhAU1y
nQFKu16lYj1KA7kaKqs2SmzjF1LxUzx0GR05CxGGpChjXTDhIEKXASH0kgjKAR/lXZzd3nD+z0sf
uvXMfSfG2shUVn0BIKxS/LVl3iSl98MFprEn5Edl5r3s6z5OCCIFIPNAC1Hl9XW8D/XEv3Tj1H/W
m65R0aEkWyX3Fkub7mn+DA248L3ORxJ5u1Zkkya4WfiFp96CAV8T9YstMJRONeaCzTKAzA4T2hML
71vk0DufXpBp63hm4u1J2xz9ZepJ4fqkQdjbaCP0o2GbNk/0Od9eTd9dXiUaAJPC/H1tloSXTMET
JW2gar4O1wqlbTV1Vf1OYmiwdFYyPYVwEN+m5ypC8r6J2sjj5cYiPxz6wIWXoNGWWz8WbRqMld4K
XceTDVGBFc3Buofr1E689lGmRKlyLucadvdOKf/0VKdTevyxEaJhja+tB8xLHl7k32cbVkZjZZy8
nBt+g9QminmAzcGoqBy5q1CJGwXnavJBUf20y28exeKutKcEmIVADXtsaa5mrdv7uWy8JejtL8Qi
akrq8lnTSiCTgFz+EqJIi+1QLClWuP8hMCcNN/5mq9RK5IMzz36Wd6Qrw9MCsgPLcoWoto5J+sgD
572mBlyQJ+ijeT9oXqdTvwF3X+t2btiMeVKSHKRUqnJfBMTTSZGWDf5URpzHqNidOB22mk4MwTGc
o8vTVS9gdppucgboflyo51Sv9J1QGlxzLAXPXn05/ycBp641v15FwO9P+oC1Ji9eO2DcmmfyoP5B
/QCkF2fSYxDM1iWFJjbyTGAb0X929uxm1Wrswr1TpvbHMWReoOQxRFXeI+JGlYuTr23yMwHGRUMh
9jPjqLEfgCHRKOd2Alfkd2OZ6oUH57pHtI5WrN7rTQA0QJOM0OSp6url+byN5RSzUZwWT5Zecw78
EkOdxLqoNV5+wShKctD/BVtHtUEamXqmoOBECrVpkhA5SxwxIl72SSxvHsBh97SuOCRbqQ3+89gK
oVTFSySZ4nNCX5MnonXMtmookDZ1If9b5rOTHzGsECNQYDJkKJBaTY1s5BvfpGeINmzc58PyosIZ
tNfcMneUowNzKJoitCBOAPx0NVJQ51oCGLZwPi5lUlKlXvRItx+/XuagLOMHlWPog57C/gSc2ejm
JQ+vlrQ9gmdvsrJFvImAIKf/TY7YTfKoeytXDtVnT5AGr0HLfB5LmkbRnY/AjNylXgKsir5wDAPs
ihCW4NOoiVPRzITpF0qMfnQbnyDo/vGu0y5BFnJum7deklIPe6jGP1EcmDq9RztRxZbPmMBkieEC
VtcnCnVtNWlNodXOhOvfzkSfRsIY63EHIxCOnB8/wk7VAmB0uO10N0/zsbbWzgv3LPd1V6D/AFLW
9NHe6aDnC9wCOeIjRXIHolAw8pzU+e2gvmA61XOPRiCgF367ghXq301rf6psOvIHz+kmc9kN+dl3
GQhdDgsd6dYtPdqeJtsvhlqzjyABYB33qIKJQjyVQ+jxKVxOMz60M9RAblelFoJrrh+SAqPrzGUa
zxjAtMIQwrmze4Rx/GYIgReYa2Hnw0hc9AWb9zBVlR9Kr3Rjr5LrMwENJ+dOqr+eoTzPePlX/vny
AWfmt2Bil0+FbnYbSDUcOb4HLIMBmlbIlKHWNnQ6PVZgaZeSWCDbBtTWAqbYSLMbHX+RgHoQ9DIK
YGUL7m9fWHG+wZlFihgGA4T607kUAMVq/cgVFYn3vqk44rg0RZ/iwaqsa8h0NrvHc3Fbw9rb66+1
iHaFQXI+52NatpQ/YAWM6hkNEQFlTdJDGDJPRbpxUv7GI+Dr0IEmVUCSOxULn8a7YOW5pUJOz8xp
MJBGV0zgL9u+IWLnkLb8wyNLZojBsh8IX2jqJbo9aXP9q0Y+ojxPbhG8bDo0TDuwk3JV2+Flt0n1
DXY8Uf+fELUYWo8l/wd2bHZEjCXhobtVpaLJI6jbjnYR7CSxp9/2LKVaaSQVXG5ebTuZmwCL6alv
0/gukqz+vRKCyoi9retlMXusU99ATGKr8brEpifg1oCt7X8wQ84mowfYimzCR9Npsh8KtseCkQYO
OqspayKcMMi1U4mH+gq7Vn6cbhcJW7Ohsw7g42nD9C0WJf9/yCWhx0x0jYqqDGd6wmBVcBKwJQdU
uch+J21yBsjnpeVSVm5beShpU6KAFpusciOIRxDzTvCpcAVLcYzUCbE4kF72FRDrf6ZNuxmKAbEQ
3Pev/6OqGpYcdydWexX6ady8kLPZEvDoKJj7inYp4+nVKNUPFhocxg42uy0lRFi9CG3FTUWSDRrN
7rGrgqBoxyQJe0+kh352RJP1Dz022gNXOs/HuRAH90D0m0DphZ+X+Z28DWdumUZzNataKuDP3ywp
/jtzZmCN67BlrfHUld2DE4EIAqow217ewwxqqCpCbfWdzaFF4KZ4pTE8tYNe4+OCZWlnA4jdPpWc
rGX7oi6LRxpgnsmrHYk7j7zRSuUfRdDKuNLqQqFGklTSNIIkW76Ce9Jqshf82geZNeSzdt0ojG7p
1XCjgYvY/sTMs39lm+FlBW2rI1wL1ftsODj1bU6A02pwkERBnd0wMRKad+e1RbO4yI0uWTE+FLeJ
tjcX2PgGNrCQkrUi5uSpO09vbbp41u/MwlotZCxST3IUSxgl11Y9UBqWW+HcUrCDebWcHWwvWv8t
z76hexDs5ViYsEcN96c/zAtvWep24y1MxpIzNmG8s2PdBNeK9MmYMkQxo7QzHHiywaeajEk2cLm1
d4nGn36jJ5DksxhraUjwsHWSfx2NY65Y8tIXcVodiI9Uhgv6+E8DDKI4OHv/aOBkcdxwP1/YrVMc
vwzzkRgvKdoIp26frXVve3CbcJZ8OBWaLZpxflA76/W8NkWSZw9IpGVlPw/E2Q3ECy3QY9O3wItZ
C/agP8tKiF2WTO+1CjGljFNY/hBeyANKGI9aNXLQAttMPT6aqw7GljUwF/8Qa7FfeisxjJ7Vg/Gc
WFgn1dXUern0su2MZkpYAm2Jv2NPFttCbW1n1QEpECdcpacxIcYTOwR4RoHzNm3HLf4cU/5gzBdN
Ife+kdiaxZqY9xHMJms6M76XhqtH0Lngk8kpMxZP1GapBmx3FlQs5VqAvXSw1qK3KRAz0KLrOm7M
rc8STEXXmuXd0KfbmU/19dIV59X6ddAa/siuwHt3Ol1n0p0bDGEyJXmMXTfo7J04WU33Xiqsbwvu
xpfLKD3n1YWxzswFGYT/EnLjq/XSt/QoT1MBfXxEcPraVzNtQj9vTi08v1Zrpo/6scQMM/oX9N6r
s9ElWjETvTcBRq+S717JjmodwWDbrF6VvxrrQymBXvowSr8VNcRJjrWurglkxM4Hh791FZ57pENd
R0ULWVOkM719Y8ELlX73nTbaCy/bGAz2f4LEMLIzN2wM9Y73uFqYNivjDRbujMTic8yPJRBm/Mts
2oIWVvmLx43r+YYtzEgl+GjHdMrLYBd35yjo54K4B5tbZ7zg+8lInn265s4CZj80COX5F+V9fQqr
AcvDoq4/yWV3rsqKhWUt37uV3DahJU3vGFZ1TCT9Ke0sn2czpvzEMvSt5MN8GxnGneltEFS/OA4x
Ih65xeT8SGwUOcfMkNw4sMShSDpOprsafjcfwcXP0/HxiBNt+KiICoOU3XrGtNOoYZODnx9+cYEi
3D1urqdANAuFlFsQIPvwhoMqQVf7gX8ZUK63upemQNdALqwsyXZlAqwdEzQskK416QKObHamEcIK
rfWIJvpUwE4pjno9DiBu45/994MctLX2VyoWnTEVUXUoEqJAJ9d4CU58LcYVg1Ru9Wfdkp42Td+w
oDW0sdUG/IVmJNcguOkoqpqZXZpoAUtGmiA4GtQiChPCEs5GOH1aTDUzdJIVbW3GWSvDMj2yIwDp
CfFFr0RfcrTiuYmZm1HNbR2OnZlm/+rcM6pckPu4UtDmOJUkxAxFnyjuUXQprSEKCgq/JsMxa+U4
LI51AmmLKEYMPCYAEa3YecxWuA136QCoBcfCCTLww/DcImTyW57tQwXRYxbdYhFYn/ajuICKdGIp
sONrScYjB6KeHjwvNPHxNuGKKlzLHZb4Xas4BdUQdUYmNHcKIkz9SICzIG673wwcTOZeTZPBKVDN
Oirria7SdaILqt+rmFn6794fE/ETcxSRY6T7V+rlVxXI9hjXadG4aJAWFsl745mWO5BOLbC9fMtc
abemFWJn5uWwM6d/yOg3m6PUYgFTBZ/AtaxMZpud9j0Xp9P7FGsvwfKqXgfktBP96PLtDMAY6tkF
kwRnI0E4yLPKNbQqUvCP9Uoaz7AusACOmGHiaWWYhJmOwdBn8dHWcWbkAn0CmoLjLvVY3aNQWfIR
6fxcFcdnTaR+Rp5DvnRjr4xCbKcuKZP761Yiy/XbRnR6Ohh4fAsNoj19mX/OqjM+mCiwK0Mu6aiL
2PvkdjlVtEVZG9TXDCdIAcuKA6mTfrND6oLen25A0oTSK4YalbpxzpmMtndqo7BykKDa4NpPG3qQ
L8Sb3zaaA4FNr3e7fp+rm7sVKeKn7bd9qrXfZ5oUZwaZZ8bM8fBFuBXLcLzjW++Pc+IJZEUTpoqO
ozSQ99HpVGip/DyFrLAh+ZR0j79xECfPXZeJPYFmXeN/WfOgHSwPGM/NnvXiB6cIGY/Xhuw2yPEx
DI0161jl6RmkslGxMiI5UcwRNmfwtxE1pncnDRelDw6LD4tKbnB41u5tVU8PY+r/yU7arjhOL976
GiAzUg2dm97LUDo3tXSpDF7muRPmo9Y5y6g6ZjATVtpZkYLzSiO4yYqA76142zNPypyHi1qY9Nmh
uCbUjAANMp/ioRkKj38vvGW/K2f6OyTd7v5U9VbdtOzBxJUDrOT5e7fb9itqR+1qjSdODxh01Z4F
MHDZ59E4FUjrHokSr6NqrgjMFslVfMq9qaDTS/VXWYhOxP0fQ5B5UlkmHDNzK/t/sx6yYw9O+HqP
9sVCrQrcjdgVVcWom9p6NANYy6KC6infvnie6yxthJiDgwshkEoph+Umyi7AXMcFPENigO+KD4tY
qnaVKgDuKuDGPHk8rr2y4D1lnqyc3TH93zB0cQNs4qDrYQKMYmHv6WokknnFQBy6aC3TOj5Fgp9O
zXQRApuvMYpBAflYoDZLLbTUAkzJ+rHTRpJjFbE3YpGnFfMPfzeED02oJLjPc8i08Nw8AOypRxP4
2nfVmflVFx6Dy3Kna4P7cC+V+w5fcma+dY0GEn0UQ15w08ZAL/5oyY96heyArL+Jok70IzGb3Wz4
75fC02/kf+iiZ+R1CpNhdSlheJqRv40ytUda+1dU8qgT+r/bEt+RhYMLF/f9DNdxKTeub8Pin2oW
38QfhCh8wwMkC570kuoUFoBqZ29jF7SafZ01AX6voTTG5aSZGEY3lgSLBozBWvRlg2NOrqptytuD
0HUARDI8pFJhStxCwT7IbbEUfLmULFJEq9WHZNShasMsJZG9JDVtECm3bHhz8nW1qw07UUuu1B1t
qF2tRtGuuwsFwvvka8+YUIIhHOLrGHtucqp/g2wQFtWQHaxe7s1/5DW9Ev2dLv579lrIllZSJE+l
wYcUZq5AvjagXQToIy4HjaMLhqxtAy1c1fz/2Z8EHw0MXWFlP+0ocL898sY+qotgmwoDQVs+nIq4
WydUGkocgCdVCog0lAx8f9GPJbst/uZq+KrQIt6HT26pWreG+DPLS8eMaW0BZmMv9SQ1LkoRog9n
90GGw+o4sfRbV2ZSI7U3jDpv746PQc5ivAaR+B73tRVP2v6YAk+5kMCQ7x+qoXBwpyIaZKuuy7Z9
R7dqrXeojgXJyzAvyG9QzBAp29p1ETHO10nG++JwvaQoudjZW8u/aGnKFkqemIqEetbLfn8oTMTa
dYmUW907Uojddf5x1OR+89N2Jsfn5AO9eWCLfqWRHpuEoSmebcqJ9yWUCMrdPjiLokFlmYlwjzsP
uBDl/6zilQ3td/hNeWT4UdUjK6Vyq/My6MDbqT4OV88VI7QKWZd71ity62A3em94n61ym3nWjbSJ
11Hw//RSxEz+EVNWv2S4rvqiQZPCbOLyJQrG1L7ld/uu1+V7W4Yv5WDVANfcHlp3f/kPquxowzve
T05cdbv77vWVr5RXHP5NnvhUegAofWm1tWBq2ojL17brmQjpMxUobevB36wF1FxjZlPvpbccsiXd
PFj5jMrhWDBD65MNacYtTUV3PeeQkc8eqf7MEutJFd4cH/L493Ki6H6TMMWjicyAFy5CO6irLC99
WC7LhdYGZzer9N9r2z7vMk5y8mxacf6AmqoEnWi9XSqHlc6NYhAGGR9OeenWjsCDTq9pEehRE3yD
3VNBuLdLnR+1ME0WqGQ2TJlZc3rVXzVcIurBg6bxNLI9ilpkHWBnVULcb1pmt8BevCmYinja5i3N
Mo/cRH/UMHsnLbebtdywIU4BMxIRLAmQevjVkzhCVWHtA9aLFWpeR5pwQdEDl5nd7b92UiJZHmRb
nYqr3q5lRewu0aHgUqo+dYZvdYyXnOxI4YC/ZYbFTVsnOOzFtSx8gN6r5zUjrqVl7lEJFlh/RV0H
c+yB+Nk6Lysa8FVQcuD0g0en/ND0g7QoX4I+OoqRmDTecRzGQpHoC43yhmaiw7dDQorRviHA/boM
kqiPVDJNB+DfNhm2lpxQXUaPNa7eP+4SeAWXuM9KRFWcmJecebBW0C/BQdxnhNL7MMXCEeZ98Vhl
/Sp2zchv2R8peZ/rBDUkH1MmEGW1GeowMIuANrEcO02JW4kWOtk4tVc7Bd0hEFmjiIRR3Aibfcp0
2j4EsUZwATrtpfQHzwO3hPNQVbFYXDJhooG8majbO6zNdqBJKBxxlS1FdVI8BTC0MvQjOYuDMbTe
zrs9r9VFroBVPl5uiLlmbRBIKwQTnhvd5FALanSwHu0SlZRqisMU0vZngU67p+AHpoNGwHa2Fu2e
6Vd6pTuAqcJbx5+jAweFv6LF85S5K026HfCxRi0hcLXXTRD50vECMt3YcqyvApvuJ8BtmxEx861R
1kd1hVzYwK10Z8TJn5DR0fd9yfEGi1IkTGV1bcsj4cxmnOByUOa0OnYfKE3MqKz6yd225WufnONz
1opOKUd6WQKW1Mdg9+N/uH6vymdLjlsOkxGAisjaLgj0irrzcZwn7CPX+2lI81+Dh3tHNXL+zX39
o4Hir1HpUMCjojkakrencaf2Ue9dfUAasPjyA+D9cLN51JdV8/yoPfiz/lV6JJRLwBNki3niB/+S
b8BVQRkGxrgc2ZTyySjc2HjzGsi77z3rcQuAGHCUQw80i3l7LDDDeckczV04JWJraxV9Lj9c7Mo3
xTuVmxpWEjnAfX/+EknYvW5saQjiA1r+/pfjz5kLJXb4jOBPa1K20PqmWM62Xf7+xTZKaS5rtaIT
X+NUUUJUojTt9naPoa94U6bZ7Erd9Umf3+6mDWC97Eb/NYKenTdW1W3/yLeA45xziQ+UFJwj7+d6
XuNfYJsFXEsmneuDnpTVdrAlBAX705MXnje3VrgpNjnjEFOkOFfvCoESgkJ3D7NU4RNNtycIj2PW
RBkgDEzqOYSduHGDIfBelluVmgfv1Td2nRYEnrKDbzbwqpZS1SuLMs/HICyg/FlpgLBjay9YDiKd
ga86MRSomXY1nmiZynrnoBnz5z9hdD+ey0Yxg5xf9mgrAGZ6VLev2xzfIJLvS/XmIS7MORVe1LiN
qJb5HSMLYDW4t53mi+py1aOCSz1CRP6UX5RLrpYmJQMZiCKxLFmrKfbMShSN+ALi3ITvGAwiief6
TLyguSX0OSZQbeTxipC0/B846vBxXr3YVltM46Ji/htE1C2m7L70aGM0xOCVZr2yD8K11PErUdwu
76SuZ//7YoS+S7RmDGBFZ+fAso7QsEuJvjB5LlbhJfKhAi2a7FVwY8WZfD3VWrI72u2b1apZOEgj
jsILg+v8PgHdGSxA1HoGHGbtuCy45bg9AEUI+i9H07y0ik+/TBwQfFqNPwy3FYtT8rWPytbh7qlB
WRCSaLZnQl1hlrx5pzbdLImRu/7yGZSRLjjony+WFpl1a/dyW8akhUnZXDfVQ00HwKHoTi3wOJXm
qJk6yPPmnAyfARaN1m40N1m+ciq53ovNrDIQX8Q0a8eGk59dARB39BV4Nt3oHc4QscxqfLbwBsYu
CCi89UU7jg6PTFaxUhDrgbECN/wckkZe4GsPPFuIMWpNR5+BF1Pp0BvFGYWKalyC1oENzpNhVY5S
arCZ8GR11CWLF01GxFDHPPn4SlGmZNV5JvSEAKyupkmQahBz0rjpUNkmVmtj5xHuyBc5V67WuWcb
B2S9RTKxeZo8vaiJUPR1b9h9mPbGaCiyEu8HJQcoO30lDgrfJuTraRX59dusjvubYxtFApUb8TiH
YxDWmC+WbKNS90qhwni1KC7ipchWDpJdC1QzgqjL2fKK3YgWOYSgIoDdaoO57tQ5D3WyCGWOB26b
P0wSs2WUHUlP4NzhKbrf3XKutdfnENWBgaE0cmXCro9R8FYE3FiM67hL+XbOVF417eF9uXIQBAre
GYUoXduZFkK0sKdvMZebfoODdmJbd1e+ZalLykO6KBNYaEysFWkrINDE16umDWVOfoQZmcmvxkSw
RHlKLyCQP8nD/KzxIl/eKbQYue0zLNX/nQruu0FU1ArIIPiYmvR4YXOgwYFZQL7AsUysn2uip02+
nOltPbnnYS4gTo8N1TD7Rry9vsvpv3KNHal1Xg68E2q6UmxXNvCNvp5beJDpu8eaPPBxH995O82p
WjuuVGHuc4qKxqipOALrQ3h0u8hjlCcNxtsFORJPbugm2SK95qdequmgGcHr31/1Fyn1KIP0doWE
hxFPJ5ENlayCzMer3wkRRJropi2F41ZOiype6f3WFUM9EaB+QW9P0QyruAXKDhUINbCqcKSccbBm
ggbOun+jNAMtC5/Ogrzk1b6/7+/2ej35OLN4y6djMK7Lot+EmmaZKNz6qE9sg7ZUbF4yZF64YugA
Y3eSP3+JnlQzMhfGFlGl0rE8NKo2dm2TDpdWo+7WxNi867WMqwZtT5MgaSGRQwEEVjsdmAMErpvC
NSbBcgmPyQottr03hnmDcEHMwtk82sxKyFh4M62V4vzsRUjsi+TZ9ioFCoTlfj8CqfVY/udsZYE4
GtV5BYy8ivd3oaF5bZAQxkZYpdtYM2SjA8/lE/ilSn0Y2gomTQc9+rKNbQnaHfm0lOnM/aGYVWEI
hDi9B/oog/rwq+KybZCr57a5tqwr21B0xd0iiW2l6wYKuEM+EajJQyUZaHYVsWwkPBk5uQUBEkg8
bZNh0CrpCdlILzurh3BMalI8vsNpyLmaP+4o1507t3fjlS6m8+cfO+8zLQOk2CNO99mYXAoQsrIU
BXceJjzkS07t3yge8zuH5/xcd6ut7yqxmuZT+1YVp4AOcXBHcC/ROLnkFhDQbMJ//PU6kqCG6WNG
zNkrVU5S1q5TchMWFNJCuAbaHinx5uzjeWl43XqXeEoMkj7BzO9QLFdMqSiC0Sw5SnY/cT2iH60C
RqGmL7fOerZ9dTwwpz6Un/xOPN/dEbS8/SNBoAftBZcsymRFGRsev9ei2mkNdwpx5lU/oiLeeTCy
Jn2JOXSiEJ4duOTxHW7h+C+shnltbHMD7K8R7AHTRefMq9QFRjut8+lTCBlA7skEkEfb6wpHsRtJ
VFHWWjx5ZCjTNAks+sqklX4fJDapx2CNg4/HI0Z1xmkdGO4shBTscjTcavBmFDkIvSpRZ143f+Ip
pNNXXYctp3yDRGfOIx3bY3VnWsG6/B4WWHcL74EizFYhGu/w6qBeVLV0gP3RwGH48yF+lIks95gM
kd8O2wnnfCcn30FOw06oFmjxL2gMri9IRvAkcDLO53xTYPlmrx54s+NJEBUzyH72gxDyXCF/zsnm
BkYr2Cp/Hj9j8HMUzH2eVYgLFkIvPJKnjGmnSRPE2bMAIFurZofkGlCQStM63l63kBPrVsi7n00v
+kxsVWjR/KkFHHjya5pT7KEkSVIuQ5rVMT7wNZcE+BgX0GzRLnh3CqJRLCLH9nIKiJHiXB/fGRFp
2Gpeh7T+PdoDBd4H7R6ZowgoqzTnkvX3wlwFjcoa3S8zXdZAd2A00I29ruW48gnuSlZX0bhBeWpa
lNcAkbr1oTiJhEg0MVc0Tc/HNbHf0KaFScY0TyckSGs+zNbqMPAJ+3q0dQ+a+bEBoTSB+XD3syum
tCbd+6sU5vPVYs8UeNaZ1wH2sdQ6H8ylHj7xZZ3RWYuQFML2zSjHCikkWlxeAjO4ygXq1c+4LBMz
1GTdmCN2svzDcFZrV66wWjcGmj+uJJE5h8itoX2N1pu7kbUVheDv/n4XnxdxnPg7EveI8f+XGMY1
l+lJsRRy88UbHJIYtXMfSRvXWRwm//tLAG5I/vjoklbiWdNFWeJlFrGmuxkVDgSzGIfciyM6lHvP
oobVDzsJEWkrCsAHXRWzgy51PUo6BX0gaK3kberlaJxoi0nl+rnwfbGEPboAoOSrb3iOBilEyAYx
qUVcGy+hKGcINXN5DsPCCOy+2NVdvoSk43tNDSZ8pL+9FWrVa3BAXiOCDXqfEk21Hwe0VTNhSB2D
bgxS+n+u4pIAcDVnnP9pX2yU6d7h87EzsKPr3lbKzyHIM0uMDuVzOBGsxcmeOA2SYK2lNNjn5/6X
TWhSx0UXmU8FOFDkCpkqrf3mvXA3lNuj63QVFAt9tZk+81lFdZzaLRiaLANDrcc36doUJDihgtBn
WcU/+tsZqUa5jBeIPMjrgVRkQk3g0c23Zabv4DfIOf6daVn2FVEPj6HYU0aZQ5RNifBX1p2MVR8D
QbH21rDuIXxENpPg0BxT47MvjkzFS6grtZ6nAkfIG54BdZ+hY2uWj6H8mH5c9OwEks2YqU1RvRBP
88Rag54Myh4s7+kxbUG+xwxohxDGIryhPqvK1czuqwGAbai00lyXTZAQ6GrBzRjoEw8DMzrXwTh4
/biW+OkBZNWvP9WQVPVF7AYwSNXYG6vtH9Usjl95M8xR+UoZGC6aZizNISNTinrUg8Dw7gMA4qbC
OXQGHHp86twPB3hClR2ybnmXb766w5r0DQjlGUw/3Yk0uQPHZoTKFNxwEp04+v5HCitDr2PSyRSk
IX7BwziYZct0ojCEMMnG/qdwkBT6eZcFT+7KdsKN5X/xOR3I2dlu3GzeWNDyVe+uUkzHQ7Nls6ou
954IsGMtRRYp8ZTlgVOEfkhTX7jXm0lb+9bsca3ZEsghVdYyKLobpt89zaQqOQf69yxyJNN67dXw
CTUq9riotvQJAkqY9Tw5mGtB8HGmqLhwA+HKSpimlh8QGeK4UMbhLf+EJPyJtYTB+GGfvOHCIrvb
FcUt5xqhdhFJ0mubeypb7Dfnfqz0K8lzvdpf0Hq6Z7QMFxhAsnkhIcKtmGaOZkfNkh6d3iyhC7qV
Al3yJvJsYFfO6RjXoYLPFHM0eNZOWcTIDUFJ9/1VDNbXfN8J4sNHFCr7F4E9AYmdv5Gs513Zy5vU
K+rQgEMfb0iXuytiobYzZyJ0Zj2SWk5KF6VyU8hYgOPWZrNNiDor8gGTtHBEvmanZnvQMAbYQtNk
7GzzixQNPIfJ+OjNYqIip2KSWCWxnwERkMtFncrtLN945CS25o62Np/DbWr+NTQ1KAvGttQKoDIA
IKP4KyfAVsz7xPPponcawPl+PO14qrhpGQKBw0i6TbRMe3o93iTepyoFdpk3VZCRz0wIqkA3i1Aq
JuOwt64dszV5MMgWq1yW/AQ+SvGYpM5ywlgJ5jDhOVhzQO40aqpqEHftle6ILm6I8uxGWcZVQrSZ
Vj97s/lb1NovcrOZKfsMngkTaJ5KLSQJQYcXmjMQsNc6mZlQqq/GYkMj6ExAQ3kfAv/n3T1S7XM6
gemL4mCuyJhBKuyv22ICYauG4Mr+TbaKXxS2juUv6e7SPyreoYEYsWBA2G5Z6KlSUjqehTVf+qD7
/CU2pEV6Tz7cihF+jo9zrcSZ4TXJiUMqNskf8P6dM8H9WxQcPYWXidMb6dknjMgeGaUur5AzyIcS
Bmof1ULVCchH0/BqSG0HRl4Xb5zEPNiEZRYzug1K7n2TZV2J2Bf/6ITERU6xkPq+kgbivIMGkhEW
wIxNX36Xs1+PFgp0jFPOh9dFPwmTcMfX7mYKJoLcLb3Lka3oAuY/kd7trVT7BAxhxM9G63bAU+2y
mcTyCOAioHljbP/7RQ8mB1fCVnBdl5cj7+T6nAXptEjnz/jWM2xz3xkQTmH515ubnQuFHmNYHlKx
EBloHSEIZyJlMLRnxpTOWOkgwuAKoz2S4QLq+b2CFocoP1wrAMMJfUGj+GMWdKxGGsZbIX9zcl4k
tp9RH3mZm+o8xaoJlQLrxzUWfAolv63pLVUMiuNIPrpLPDr4tM4JY275Ik/GHSwz4CjNusG3KQNe
g65o2IktciW26wP+a0A8Bi2KZ+r6ZihmqfseOp8oa1IlcPypbGw10bU0tXIqiHuxcGJEGjMsDZv+
gAyXk1hMLHKn8v/eQZKJkLFUb6mHgTVACD4y5+f33Gz1BdR/pdXbH9nvmPQXELUIlXguqzBaUZkj
3l7U0+ekp7HYUiX3K9G2ku10LuEwnGPqGx7xbIrWzYWoAbTzETzKdQ+UDvGUfWmJRlwNJaiqpns1
irhjToV25FXp+SQNj08dqX4UiwxK0YWrFBRP5QGE8U3oYfmBWBCiY1ipEN/8E/24ZzLBurHB/B56
qQRyiUYQ4/oQ/v1Ke9xOmvUDAYL8QH0PsnU7ojfvf5PW8ZbTOOQvTbX2DHEG9SvVRYL/j08TPRgN
SyAfvizex/UG77MMAOJ6kPzrTTpcrrW6HI/mXNGOWAzQwQVi5GCSLK7b8ixeFsa1cMLKfThUM/9c
m12vCoeaJWm9U1vS+eRahi1CnBDOMuEtUNAnQBs4XrXE54mqwlU8p2xssoHADLJu3/BzxLwZweKy
SClgQNu9l5P2DocT+HcPqpoe8hJmY1f1NfKwV40s8Y8fdVNaQuso8zKi9syvG5d8ih409nNtb3/n
0qfXnyNzOrW5QDhsePB7eShLXGcr1Q+LKF4Dc7n1yr2rCwsa23pXTjk5/vRSW8I6FhfEWgn0juAw
AlvaIhAltg/Sxssr+a/8Syt973ml5WCAwntFzTxIJlhBitgrTUTauZcEAGsXZqc4WFA4M5yGbcb+
blBApdHuz/AEWpFeCBAsa4i19JXX172RWfqk+LCy6R8JWezx2EPC51llCaSYTWFQqvH7ZyQXStFd
TPwUfEU9t+d76F8MhooW0LHetBbNQapsLyk9Ol+cqfXOySvx2SQyYTqIH4AyjzkFuAw7AvZVaYMg
i9YtSMQhY1EygunHL1rF0QtHDaLPfFXHMdlHEHtd2IJOe95c3SQN38OdDbQDOjfmqblchBBx+VWo
cNRpSAr6MBVvBkZx7mBqFUgiQbB2uAng/KF1ixkJLSHk2qSWF2jLvfVB3uaputF1cMFGcUms/oD0
6KdORKxC3ODTSjQTOVocXBh5GOgdPMQXWNOeGI+16Jcx9M29RxHsJ+W6baCrWeb4YRKdwPE6drgA
1ea00WMxzB8hk6CwoiL+VnF8K7QgG4NILce12+2mAlDMOjCV3T1twK0b96rl+vzo0L1uukdzK5B/
RgduyaXUqwyZ/H5VoHOLNjkkSbCs8pucSj+j3mts/FQ65wp078LbZabw9+k4HN9py6gabxkfw/MC
MHYzt7OoDZjIVoziAB4FPygUvC7aPK6/J8fkFBtpM7G5mUqWbFAnSGvGZTCyV+J9nZrg3TDLj3HD
f+J70wMn31/ArJZ+7QlyFKX3JloJ4szqELQQxyWqStm5H3whhLPZZrh6Nmf0nP18YBzFou+w+ETF
wFD1CHC2PuQv9uNMf2/BdUgjeb7o+FElH6P5RMSd0YqNXBdJ5F+Kyaibn4H/q6n46MZsYubJRPY0
9u2U9EKHtN/Fr2EnkPgOpw6CYeEsYpKkR66yX/dKFzwdZuOgHIJAa7ozaU4bEcXSXW5VplphvgIC
lZRATqtx+317eGbiWKzKaNRy1wMODXWuVYY9KO9haAWBa8ulYZU4qUn/32zY1s9bIYKaD5M84+Ll
BMfkoeSfnKr4eysy3Ap92JD3tVQbmAfcER0lsag+AMhF+VD5cYtUD4WBfhgYcMtouhG0bLFXmbon
kva0PbmOimoKBGaZ82fLAtZEfzq3zprm+s3rVGQBuit4AcAldnph/OZGx6GkhJLFhQ969eEM73rt
xPCEn45VL3E/q4CPJ6vgLACxvyrt076mCKtSPdd+XSKaF8O71q5TVUypDKLpjYyTpaq+xbD3Fvdv
B7dohA1HyTEYDA4dZ8ihzYqqnAesK/V+dv1WEDN0JSTDZ5hm9zZ4jctrJTOzZtdhNZEsYm+xl5d4
RDhWvdduCQ/K5qsrY7ns3j5jh2/jp4sHzEva5Ujq4Bn14zEK4/hSEZjecYYi7BQAyFuMHADsTNw4
5AkSpmUwJvODLyDdZdWT8c+b/8iVTEOgBu7hxDgCcbEPmqcKvmnxXLKWBlb5ZIfLTF9rAcePUaHF
azOPKFZYD5opn78zURUZI8trGqXiF0ew0+f7wpG6L6q2l9ErbnG2zYvMwc0o7GoNM9IAwDTYhg5m
an06kSMTSvenNit3Le7dwOZjMfr9CuebO5yZRUdYtWYqXcxQLx+eKta3M9fIx26Zw/VSXV9gGOko
U7dqNqh9zFR68LIVQG/NzqmHL5i0K5zrUzwcQdD15PS+gRIj6n5wQ/mvsEp+K74WqC1jERfoe68n
I09W6xl8EN34cGEG91AhAIxzCp5rzsWU9j0Cz/WAh2B5lF3PuXPji7YzHGR2WkvOvzk8cJ6q0/x7
17Q9uoD76i8OWV6y3ATXtzE1wiBbbAGvxKlH71atE38y8jhNPv6tKiYQyppOUwVPwXtrc9XnAHoG
L7YMLzDy5Sfc60YJBd1fjOYFkXPD5xjjt3ozvX+8BnLfU/py6IjtTyySRkJSPy0DVdFw+NQD4LYE
T4bem2li+3S15o1/Z4dF3EtpPZCH+M0WY9IiRNM7tKEDZu76PSyNb+e0XlvUvnOPA4t6cYywa26c
M9ikLb/txF0faNmpaYPRB5x0AP9OzbROcESRw0A8yUiY9h8Q0Hk0mi5EVwrfE6op4LXfpc7lMiY/
a8rMy2BzgQ7qjbqBrLr9t033YOjuYMySMfaPl7rMGyQ/eew4FHPqBSe0lgm8BjHK9mNs9prwLlPL
dZYgli/ndKeV6olu4Fdzqg3YzJ7NWEaiP6YfC9Ij3kpF35wUnNzbGmvqW6zFWw5xak6WWbROwuRE
b6FY0NOJr5fgJ4gDAUovxQcFZ6HmZIG/VykAhAFXTIXYCUAu8M2k9bWLBqpbqJ1ymxfNb1PSQe2A
gaSaxGFQRLypqAT+K4NStwPpycej2BzkqRaumokwxkLC/z0Nr6fjN1Mjf5q6vPW8NYo4JwR5exE4
d8NqfpftdFQzzF2te2zwwlsKyfP995nrHedGJhArjkyX1dhYbOQw+GvKxZo2bVtdi9jRGFeNqL4e
n+MnR3tVDqSJ3N4otaS9Tc9lWYft5mJnCM0LSWRYGjKqngBaxJC+CLBwHugWQ/lxnlx1ELwUyHjd
pd2EsHSnlWhfHt3IAiepUi6DTWKAqWPhNdwhy9RGMXdPzHnNNe020UsL45/jaQS5X/hplpGTzKSh
b7Qs+KMHKY4Zc+6w1hyMBILAFOqyW9KRRYe2qnhMX08GJqFD94Ox3O7mHZsmRcknvy+X/OVghFBx
XugJVG8xnIgWOXgTpYP90xaO7JYLZC1ST/hXr04J6AvKoUfMIw0oIN7QV9kwlEZMxt2y20jnA34Z
wVOEe3IXKAgE2DHdcJ2rXkU5Iwh6Twl/Y75RDekyiV0K6PMekXlWwiU3NuT7c9OA99YslsVPrw1n
p2htjYUNvclvzLpCEbgvwowVR/oTK6arpuFBnWCERu3KngYlEuZ/WWyQt83iRpy934+0YYUrifo5
vrdpb5gJAbdJ8lknZeqk1QaeB0ttcbjSD88mc1Vba2kKzjFLNnOr5ZUs5DlmG38+LSTi9z2rALrl
gufT7B91JcPdigsTVoamRvDfsoE3SXAVqPsIDn41ZNFbkFmE4BQyoa/75tQsYqvaj/yYk2eZ9lD6
QmfXuJDBw6YEQ66PkSJW+qX9Y5cKPRTkGz89C1adLm+p/X5rF3TauuhQecNLj1SLhS2D1jadYg24
Ayg7HrtxKVF9Z2LTqyhD8VtWCTsR5gJSy6MnhC2s9zhVg6e5uRwTlhMuJYFCNME9vlpiDm8bHBdj
rwelrh1Ms0gXSVQzRnLtLLX6DtJQu8xHsU3XfNkwN0Ie9exlxaO2bTEh2G9rlylVuVkwh3SSyfpK
Yfjlc5F/HfeOS0lczxn1r7cLT9NtvJ1Z1t4vDrd22/R1p6n/05LKa3jiUiHCpRT5EswCeLQISnVN
MOBzFTZaJgDwdLD71fcEOBgWw+oiYMOml2w0Q5L7cZKEysE4gkRbm1C03G1WtIceIJW7qVJBPrbf
ICP7uVLOoDApVBMzm6CbMXmIumBaVy3F/kKtCj9zRliTZ4M+1EruMMcWGD8/W5UWih/YsUGCYIMP
rhsG1aFm561oBA9U4o6kklVdLGEeIlb1NAo1/1jTRWwwXWgctMfFTM0QsvRp/TbsWirjptUcRnrw
dsX3HCRNE+TnjymVGdbbhTD6u4EEFFEtskfHmwDfho7nkaZoBbMR/RBoOnT5pLxGiFaWN8jGw9oM
fsYbaj+GXvoExraIoko6evVeTbVkgQz4zOQwsut6+fej1andoE2tP1GLHRFthuCVJzj1rm7+ErxF
okxHDQxgr81hYkmvXDw7NkCbQ4IiSVCXlNe5E98phJAezbXvRrVq0efJ5uePHk3dBPaD8AFCw3yu
aJpuNQP56kVf6dPsAmXBru3YRTjo6dNWig9XGI9RQfwstyN62Ex6a3aJ1J/M8Yw2if2/KFXKvmE+
6RPvdJD8lqXyalyLKwjsQY/oOVALTMAljwFQ0JzZwnDGjX1BE5p+6cXSyeHcQGXj5OrR3U83/Dk2
QwCRDRrTZ5fjF2AQDjoB0svjl8YIzI6n5tC7Rf68Rkof0whXlpMlqgzKznoQHRhiphpmLQym8cYP
IuEXFA+E3lPd6c+5Mv0t+zbVfVEhkKBGSINJmXJvq71L1qC56cBKXqwxEqvcNzA+/jdamzo5hYEL
CQuWy0gdLse3im+tgPjPxBsKDasyNHoOVVGCxPP0w9PBGTdff0fAo65HLYUpinbiK6QIYMUPBMe4
GPeUc4BtIet6WQ+oBcr0AaZfqUqaT095PnDqqWp01ISk5v3SYWTi0+hLuWskNbvWsjlMKI2vKea3
pyIY97ya+bWGsOX4ChKMsRXqe1Gt1/XpusYu9Uqu0YIHYiqu2ddHOb7GKDe0bZJyRSmNkG4Xo0nW
DHlsSDqb0HxoN4SRTiRJJYfG3ZJuUT3HDsuzeeJrj9yr/kC8CiSKaMfqx+ANBNw9trkV2Ls+olTw
Jmi9CQTPIRPe2N2lCWl1fY5h06hXmUf0NR4DRNosuKGdhzxr1Ajel5MKRod8r3tXmWAGM8uA/Jk0
IbNCBH21xbGVvyKUgQmMO0Je33VhLb4KPqo8KY1WmDHiJWGF0btgf3ADASXJQNWXIugxzUqBIvZS
Fb+8C172cTxRm1fj5Dipo5PXmIkiEb0kwfO0CYS2AxDR8Vpoh9o96GGwkq1X0zjzZChpJY2Zeqh9
mXl2j1lF1Jo413bMJX7DI9jjD1YShpbBT/6nIJGcQiGChhzLjqU/o1v64nl0qmen5zRPZ1hCJV+5
vub4X7NOUxMR3cdHVP/kHGPfS6uYksDe600e0drHniEs7l5K0kdWitG01R+vw9T3+6fi1Xf3GCKG
U89t8XYoq1ZYIxcbnNQNkKbbUsJGuteGa5mL3lHpP6uNBBa/myqYoUZgPgH3xUATuGrjhRp03HkO
mVTH8YyvcDEymWpY2xtrAVYChDn1EYfZwWB2KYlgCIQJbxNochIxeQlLQyO8HSQt59YdrIZW/beT
QjrGuSGR5fbbFttT1+89bLdygQ+irWm86CG7ACcgDPDPdz3r8kUA0MDhNZs/16224n6M+OqQq9od
89yTifkG0mG9Vhed7CtcxZ6n7wiICWO35YkCmz6mHr1fuCb6tuxMd47DDU/BGY6vvrIPIIQzsAHN
9nm1wtJLJSkdoSM4wqsUQ1OT0L01opqU1WRK0YGX7+YysLC3gcB6f1LUVJwAZx9Z11fD0MIavm5N
mgoM7szW+lxRvo2+mCK5+OcU4XuLS1XV0bMziQ1oOwJ0wPeangFYGY3DkYoyEyrXoDJGsLdwSm96
/MNFJ3WhpHtMl2+UOv30j/7ds3ibD+tX35QBTQpk2Wu20RTAMZzudHRbQoZVjxWuLCCZc3j3pm3L
egCYgJq58FLxV397ZasEu8xpO572Vq02ymwRO7zlTUH/zKqFHdLwrNgBc6BUX4DcUi27VCoWfANo
jwvc+bL0VlaepkCLHpyqlrYUE+EFYQ8+ewPrE3NumbcxyYqxAwCC/nhlNTLijuQaHhSxQkGzR8bK
LwizyAcMC7NTDDUj1U9BuVrmiVvFnbbxwY1U8E+O5NBuAYGsj3BKdBi5MtXU0n33LtOUP1Oe1St0
RtIb6eIWgoqm1U0UZ32LCAaBGWdwHMpY6mF8lG0ugSRnfVK7P4k9pzhfoCezVDXruDid2WE8Mtf6
wLXxCfes8/OpukxPvgOZXgDjiGN2xzErNROzDr+dtMwaZK5imVGkhi+gsY+k3qtE2zzEiBFn+nQG
FrSVxX5AEgr90qTORptUb09w/h8Uet3YwB4a1yu4BCY69dyq0jdj0Us/t/wS1PVPcMCrD55NyJ9g
8RS4FrUM9mFYry+DVh4J9S8e7yDKXYxWJmU7eDBIc40TPGHlvDk73EyQkVtgW8ibzlfqbU1PQ9NZ
X5IPL8Ledalj7qdVBeXShAfxP9P+fM8K72BIdXnJwgyYsAbO3NVh/7y1kHQQ0NxpL97iA1CepS98
/SgHXcV2wGCLCiAJ7pJJTGUlq4m36s4tjphMIFJZUo+2t8eobqbDUXNTY7PMogE1hq0zb0aQ/vIk
mNV8s7olbjR6W96q4dmmAvlLEqp6zMDhfp/nec73DXHZQpDpKrw2rCnfoV+RZL/t5Z3lj5xdi49H
aHguzUvITxOT59yRIsiZxnz2Xfo+46Mop1lV6SZuz1aViXiV/u0lt3VQE/DCClfGA+sA4sjxhPV+
f8TIZCYnUenAJJlBxClr6TMMYfEyh7pVNlID6xD84kiqR4pkHloKGccVB3YQqoNqy9eW/tsBvoQx
fmAXIfhR9S4th9s8QrZVIylYnfZ5THVysJDnth7lwW8MaLqV9AsYxOQ+RO4kzxYuxaEp65XtLQjv
H7LojUc010XVwW9VTiAtbQpeImZ84rjm3RSTc6k0QlkaKiCWoyDso/8/AZ3NUvMuqFKuNlH8a2D0
lR4EPA4+2Z/jPKyoN24J1Ahhj9//YaqAumIIPj1CEj54uCoeqssU1SiN8VSaKv8iViQsmfb+NhMp
CvPVT6cU4XABlitWQGsN0+RKwK7tNkRREk2Cu2A7IJFDPiuOxVSREPg6tzp+rAh5toNrYsdFSNAx
P4/Ja1M2x15/0MYZkrI9LBv6hQ6aj1yZ8hlvqK3BrBLho2NsFbTO5RQZid/wtYhdkypYru6Ic8aO
5RJE9cnGIpV/6812sBA8ifkGzpQwVJgxjuky557vcEcPZRTGGaXjWSKqENzt/4YHs/zk+WBEqfCq
fRRXmyTGpu+bXwX6+78+cMBeKFTj7VzGrxoUSewg77gaH9veCt8jjpbQSapeq3Pudr1oMYb8Vw5G
Z1g69yE75eVQAXROnlG5J0a6YEGiLMLf4aipjfwfD1rgqIUgqdxtwdUvdDv7I0VSzzI9tQ6hbf1i
+VAUHUb6CaPEA2/x/okcV3QzHQQHtw7tIHVYAz4TrkFUkXwYck+Rt4Frn+5vi/JBcon3JmMJpjzj
jzY/pqABo6AyQD6XGe/M2aoaYSRRzkMChxyznFXzkZkjGz0/tqIE+Va5IW97gmsx0SZX7+TlE1zq
Krm2vKsoHV27eMspcVfw4ac0pm0IPDjxY+1v/AtcaNofDYtVKwUpPD9DJkDzrXmLTMvpUxTJOxKF
+c4tQVbU39MY61XjTSklvrHLRojtfy2qWiDqkk+mrC8kgkjhSVovO/eIEemmAI+TN0t2xyyfFr1N
u38SvomfMg4FfTrpyiaDKYwMZparOdYxyz2qRNJb17VTcTaKh2zHUF+71tSt28e+45OxLGLLhTbk
JVQkGMMUgZHivFfxhEGZONt6d62bifu4ozSX9987PQ+3P5y18x1aOmvYbSLXuDODnUDqUtCnankK
6o/eeQZfTzBL70Zg39PUm+aV5oE9Gkb8wRneTe5SK8RsvSjvzjosXGzvPdkXCukDRE5rt1Lb+NVs
+OfYWBOpMj9/Y+UYKwh/B/CiOKow3UjPMMIR6jQqWAQbobHJ3bPsSUZAkH+SIVe5f0hXitm2/79c
Exi/P/XF52HZ0JpQO6hZ/ffYW2FqFop1hd+Hr/pWrx8bfP2Mw1l2CaMOFSa1UvGaT3gxOzAkk9kM
wj9uzj7liV/qfOwQ/9AKPMr5sjQVnKBTbBF5oYJ0S2M79wPupY0vq9KEhOzZ5n9mYh53A4SDgZhu
/9ZwEXJ62Z8ErCb8r+6clEZQlf5fljoIUfL4pqwD6+u/Mqs01iTmHRkdHhPA3io/9l0b2hJfIMBB
1HNcqo052L6daJ+ZpgTmviBNiFikT7ayANd05gDHN5eHFdPx3QGb+g+IRHk9cbqpyreW7PnB2Hot
sk3RW5GBvP/I+vw942SxIfDrSrC21LknAFCTn3bMu1wPjygPepm/TQE8gcPcLYhoXMyGiwM48kt8
Dt2L2sLC6bv6O1Bg3vjgRQ5zIUWWPTRL+BF6RR4k0mneSB2g86jiLJNg3fkFW1M+YYP3jr5MpG5L
JsvIVtJqptakngxXdSGHEoKVe4sMUvqVq0zNZK9kHI0XfZRLc8ROxAwap5bQkVP7/nYmgAys9To5
JRvv2NJNLEJLQ2tOjaJ0hh8MaIzHzlZ9lftcif5xmD6YamVa9S/8s/DKBRxAJgZOiKHDnLcWe5BV
YRC908cAaFmot4ubJX4+UBfWvo2UIDrpxpMNlVk0fqDsYHpLsS7aP+R5Se2rPTtoEPUKkef51vAE
xx06PCjcNUVDaPEViBQq5/OLjQy5Lowt3Wu06cbZ1Ux3YC9hjZHGGfcKkUhtYEkqJxLZT85t1nI4
u5lmH5Yf+gR/iGr8/sS/6y0V1AVE9RWgfl6QTCLZLBZpQ4UoRXE54GVu5sRVRCA0E1tTq3pRqe0q
o4cQ/wIyyxtQGZ/aT0NIalLEXywLKOjQy4twzEhgLmtI+Kp6WT0WzsTiM8OwuALXC0xnmDsxS64u
qfknqDV+ucnm/F2P+ENSySlTt7SwWrsU1FKjglNJuygo0uLaBb6ko98LQ+51hLfvPd6AUQLnKLgt
IJvlhl/hofePivODaWac/aC27IpNiDXa8299PmSDgOtMuvzSocnjxACPTiZ4EGsp+CbUK6UNavXS
1Ut3FX/K4nqBtefXqxerGlLsSUIjHb+PbqFl2D+bSc/szl5CIcNKOf3gdLTk9LGQVXIMFzn8wcVQ
w6epFYqqyUf2vXF69etu2hPYtZTApKSl6JwmRSIAjY2E36oQxCh4DQLtnib9etu1empDd/EHDleN
JvF1+UWUteA14lDrIylHc0RL3vHEJfN2kGBaMx7QZWy8Tx8EdVz1CJib6RvhiIclb+XTEwwHftyM
e80h8410007mDZgw74rQSjkbi16MsOEXcG6EvLGL/rDDXGY7hFSGQTxHYpGoEFYIoksxNumicLFm
PXEkzNX5FgAEZ949oGzH/vinDDgblpX6WWYRDUFBAbm1DMeiIotfQRd5/ZGDfNJa8BdiPjQGg0Eo
Dkcfw3EGwBR3NyoucoxmQAtmGg6vaecfpQ9YjqheNHA4qV3N8kUGTsvtmzLJTtWNR+KFa8GPmQJ0
O1QpUm4KVp1ABbLijLFaIBS8178seXkBUgtml6GWE864ZD6jCVLC9BJ/9861+knCIfUD2NVJukzD
A6SFkuAZbipg7qBi2MsWmwMHLRT4w3QVPiAfqReBkejyvWq1cqlC9GykclN9zBqHqkZNAmDdvOo8
xlohIwJ0U4MEffGTw6fJ+W0CkamPAiScCdzT4apCgQkhOKp2xwl0v9OXjbJ014KOOQfOtOy8gtlq
dM1ReKLWLTIuHFbAZehRZy6oH0xLMatyIIpD5Iyl8wKIvE83t9PXgyTkkMnKHP5LpYrCPD10mrny
UxDNz/PAo/EuSfYjSFwLumyEzjeU+2KPRSaOy4T0gjgZAkyjdrS39r1LIxj3pzbkBnm4m3Qlw3Tn
ULEt+Aen77sHjBHbxulUS/a6lF974pyPIOW7nruAM0S5r3stXZTr6j6vS3iPP7D9n5VRgeQ3jtxC
XLvVsK6S0MYjLn9iJQbBqB8PhpX5hAwLYi1rECrwlCSnZfjahycI/gGCfslXlLFANI+3jUuQBSSk
q2CKlqgjOgbejQWANDBtpEOAM2wSn5ldxz6NDNs1OMafADhY6Rwd2TAUc/N6SUL+Go4qiV6BIuJb
5eIQzTkcAMGH3qr/WZIotnZUQHZRt/OP4MWFR3DF1YODcuk9voGm+K6PugWkRWfWhg2ZbBFRItCB
6eMjSalA0Zo7JhzN3/bMv0dQOP+EfwCWJEEcobo8e2//C/w4atPuEz2lA35YE73EB9ErUfF37oXj
QaNb3dK+jh2DsXM4G4sHohBgnxLEWgH7LF3ikGKEgf95AtXcBGhGgXfilQ9lNZXnfkFBiGGOEuQ1
hckTzyNqar2nxFjfQKqU5SN2xWPFNDsBn58IBEsCIpqn8AKcqjTECyURcYrhROvh9Z9G/tV+QbV4
7ZFsZWsJVxtT1+2i8U+d4Ci7ezrkWB+O9G9XDxi0t5jXb1tREB5pO3zdlW+b0HAgYRRvxHC7Ye5V
5aVfNVoJAF5DT99zkkQCjdnF2kfyNvuOWDmh084GEYy2zDgcdmZeZOyUi8HSNXXaj0AmJXnLQakG
I5M9AaNEctGIVi4k3GcHegt40gPvo2FZMLYcjtSoB0J5ZAvbxQ/GU26czDK4CQkUV2O3WpQsXo86
mFu2JJ7lojekr4lX9HXY5cL22T3Ya8Yz61I5hLc+Sl3+TZtu0X0bYb/wX3tTlPnugFvvc/WNY20k
LGAqEX6htqikLIZj9mE9Droa+HXmhxDOe7xMNik/hngfI/XH1bcoHvvgYZSjwYK6PX/lpa2Ias7s
tmY1XC18sl37gorIGPzW+zJZhoej9i4WHVdDIfT/omCU5b9PbCzCYAasvoFKuGNoAE0X1aMVCjHz
enJLM10RAh4JPpPL0lcCyMQpGm+ocJIm5K/YaHZ9nveCgBcI7wUj16vwF+99oef+imziub5jVmOR
FbxVsV9N3/AFPG7S+8LlUI+OeH+6kqh69OwPkNyuA7Bc3X65AvjDg2pnVdfXq5SEb6naJnilt/kl
9oY8suGOQuck0jWaKfddrZieBssIjhqyoZ60F5N85MFxyBjscMPWcopSzK2PU7WlMLC9WKbKJisY
RJo2Gs1qKcWQNAgO5RH71/Z1K8avlu4jWZxUn0FyviFDIK5eZdakjiePFUceoGtElgvm5w5V/CB1
rZGvW9RiQpQCNzBHMjCedMgPv86O+UehWcLb9cifqULzf+QoXovP6Y37LPBpQkgMK8hPJwl7fwTG
pvr61f09aWUoKyDvaeETN6U8fjD2e5OwdKjEsC4iSxITGDgybiSSnRi64ca4ftrgoVFn5JrJV8nB
JuPy8tGCNk7ZlPACGU13X8FpGAflYIB1NQWdcEnFJpnu2uZg532H/EdoGwIIMFozEZH4KM41oIb+
sH80TYV5ZShoJiY558jgbV/3ueIS2MCIFRJy/nXJwQjZis8PCbl3nN5VyFyxFvULcWja6sxSoTpb
W3ZqnZUH0lQ7uMp5+C3Wji/RgopG16ytWnJmo4LhccADb9zgJvUvY9QC/OxSaVDOY+T35HFcowkU
7TVer2eug12wjoc/lm2PXFVyEvfee2rb//qZjfLn1MOD4ZdDgXf5GGiNexHVfAlOTiphu2eN7JuW
k/blxjYPOg1gU2/vdF12bLgQkEaJcH2aECRX99QrSy6DNTN8UvrDgNJ1872uPMOdaHo/ewV2xzsO
s5IIzZNB0zWFRCqHVWb+lHhd2y+Nq54kUHqnASQEOZc0WlPd6uoA0bkaiwxKe6RuWaoJcaHgqlFI
xfAuU1TknwxAUDsDpYb1lP5a915YxaUAaM0ovE9NLF9WznrQDCnp+WBW2zQzsCgZi9C8e8Co1Eaf
347Qt7hbuB75P4NGNV5t7Z2yllKvBu8w//6ddHHsoNXu3hgFupQKjUOUyk4DzjcjeZNO7G42BmdP
ZsaQgoWjokAyz2cbqMbLeo12sSkdJ1TdzmUXoy03ROzwNXCriAsfZt0XQ8lHZGYx2jnZZGe4hpNW
rK70kKtEFxzeb/8YJQreCnVRgrP69GfcCWp1fAWcjbkpolXKrR/sjg2N3IRxVkPikzS8T/voSd9e
zBVeqrKNvfuVoVtknPwf5Yvg+vw5TFqASMJup2nrqICePWIxwNqiEDXGdYteSbzToMn6By8mBL5b
awSRlg9zzrzzfSKrL2SqXZbyVcpCxmHfZScwkRp/HybjuB+3dNwILBaTO0uQeNfpOiCZaWUGyMXM
kj8fT/ctGEoF4rLjUI3ChErdRh3UCJeRKhC5ujOkgo+LS3vKjoq3ihQPc9/2hIM4eAhkmDw97fIK
LmVpSgJyGskOTUW9vbOv0HbSjM+Xfcw/XNVK1dFen/06unTzKBdwPyDoZlNafIB9UKSbk7CSs9He
F7u3xTsp6pFBjRmuepVDavnQ+OPJRQrIt+vuLwGjPWzvSQ8R1jVemJeMnqM5SqbTTPPOKanNEUMu
Hdo4juxGBnt/DUtcP66j65hRwjMsOR8Iid+VrIomCj+rF+O1PkRCyt0bs6+mtEEE6jV+PR5P3X5p
I+d+YWqaHt/C7ge/wkq7C4cEihNqWR+PNaCjkWLM+iAj2tTVUNqtnlp8OG0gAZEZicCz+pRrSq6/
pR79fUbW5iKNQJ1pCSKUBBXSNVWniOVm39uDkpnar8Ao0MSqKF65hQBff6BN46/YyE9QKjY99+em
vW1Lzcg0wfCc5Uv41HPSCDTFOL4z7Ts8DE5gdrm5qyeO/5vIg9TsHnWRNs+VuaWwSGLIIQ6bI/kF
OJwWIaZTfwr6KWNJh/7ydzcvKQNUDQwbX07eBae43rIfbIML5QPWEwKzKfI+ymxhoZS4RmryROB1
Q3EFm1JX6SFm4la2yQEE4Wyge8DGvGskJnbPQa0otf+OM1+nNgvTf8XIS27stVwwixfH0JNkiGXC
yhyUKPwO4KhPlut8+zVaia2pdNxrkhvwRakrtNjNEcPQxdm0UyfQ9Bzq8OpALkYafSQR4QED5rWg
KEiTQ3Zfa1B2agXuQETjtzRdlAd1FcX3vs8Z/DNW2pEJdzV+vBdI/0OEEfWaHFe85IxeneJYmiUg
qjBKIXvYzCvaPSHC9InYJk27nJ+YHumeMucNIpb18FSd+w7VmPDG0bMMQlF5iDic9iLClim6bwHt
lCdhRZzgT75a9j4mFYQ6S5ExTJUAKDhBW9hWL1sYB3wOuz290PrykaV/xIGFwsd401GdW16/S68S
DvkzH8LHoG0+MmxxRq1b4Ebl8ejd9rU+pIlPBSXvXxj6czjGiKEDog28QYotz0kWaC3ZPI7MSUWe
4d2/kocyLXc6OssVwW2FJWQBwGe7cL7xcNVGhQ6yiiOJVFfF5TWaZSDImLqNL0jQtg3dv0fwKuWD
1m6zBREfZBxg1hpB7qn61mtSN53LDlu3801ex5o/5PXHiTHnUxMIbBY2UQFNf51/c2hH+jFreVkz
OdxJGE9z1LmuPKYKswoWheIk72K1NJG31QgKPgD5WEUI5jhnRP1rEnKJ3nUH3jmS/ZdT24fOvKJM
xHzdP1C4eY8U/CfnmffvviLuEo/pEXXRB+Ok+DHLg08dWHvTlE2nTwdhz40cYYbW5IuCfASbYWaR
dZ/XoS40SA7G3C4b08ba8D6xUT4ouxHGxBTGri+92zyiKa8TpGODFgDzCxyqgo6iMW1FAX9oox9d
t8IYM9mUfuQmgZLig1lIOIhWVz0FIF+XB9gYOisSs+RRMXaIe/vcXUwf82KoEZOLPEq76gp31yAG
+iCc/S95sLtE0h66eRE0FjTlhU3vO+S+Z29HySDK4yY/UGjig4+uYg+Vw3FW/4YzUX19sYZ0sspm
pTz8G9VQgxJ2sY4gqk7DtKtSqF4Ckk8sVrvZbvCT71RMXo/JVov1L7A7/LAFhXCsqPXcWx4i0K95
k9aH9ueCckIjOo6K83zwNkZjjoFAT0Y3p8ihzUyFUr/Aa4r/fXe4mTXMVkYGaZDDpO0+fSvcMpFL
nTRHcQE2arkqoPJWuDVB5+c5YmXkIN6TZbWPaTlGCeEDP24XLGSHGiXWckHHE3pJqsAGtm1WUe+A
oqTdPi16JgjoJEpHmXXnoggg6NEdbh0myI6j8NVLQVbxcdGM29GwqhW7ynFLHUeOPax3OfTnxOAZ
41okc021gvkStv39Voq/XLiWnxPncFXrg3rnrviSj5TkmqAzkFX2wZyNC9icCt8qVqzWCoXyqrw9
jeAvjJF9SXycxL2GF3ke6a5NRcsjTxMkYt3dUZrwATLugxDw7WoOAwHoDd1B3sEw2Al0xeHNPJQ2
TdO9mZ9daBzW+bCUGIQni7yUeJ13dNo7J8Na2COhHF7dZm4GzD1ntOegOt9r/2EHoJ2aPB7qYgDa
QkPDGGNKziiQnnYQiQGdoMd/8HDwYquDCB+Fo4+LWPOnwdtdAB2clYoXV2sxJ9zjUB1jxV8/Jc4E
srylhBSwXDwKtVU3R3/JdoMFa3XFXtIMhuY+zuYFmumk2e8tYX2To8kxPfbBtyDFvSdhlPuqWqDP
NxkijhJnwJVwkjjV1buoHGPcqG07gOxQdg2+FMCG9O0BaWx9LRl3H8+VWDSyuQa4iyoQdM56nnjV
rXypQuo6p1wVq3fLqRuWC+Gi2199zwU99zPTX1ZuANpuDzLww2N/psRqxqXahTEd1MILG8ub2VaM
/cNr1Fg0uUb2ypUE+ErxLE9oMHlunWvsMWWNk/y66JiZDeqBB0kH3yzzLPm9pMMz4lZJTgYjycni
/agELuWw/4RJRmC0ktI8DmBKzbZK3oyKSuQ81HGkXInGBXRqwbIhwhVQyodr2NxoqDsvLQUXc2NE
3TrZrv19FohclPeerIEkzmnW+l7Ox3nH1mzzy45R9pJ3u8U3oU5m8gTkVd69r5RFpjvX2jNkVHAJ
1dAMq/a9DD4xd1UoZKGgmZfM45Ogsl2LC4A8pkPBhqbA6eWTdfQkzjZcazf2ITNPQd9GwuJLhoIS
jXHk7DEM6PyQqTfqMm6cRrZWklTQOXKtN+LKz+9ry7MXMRIs6AjyFK7p1n6AAU6EsLYiLQCz5Wv6
qeAyRY+WTaaXNaJHEhMMuw7GCmcbPX9q0xtz4nJzQs8+acypokfBKlqQ4WjyG3v9nqd0DMt9chve
z5hL5asUKVYxD0raWbaebP2toEHtsESlLgbh7LhpFefJtxsx0wu2bBpGPE9SYKqzpPbmQJV6MSTv
6iQBz0fRc9Wo/lkeDOB51LIEhPaYm0NELn2zTRRaFAzgVE9cM54DaEukZC5vwiBvjWS4LQ+U0/dn
2T6KC5TR3QfcX7xCAZ4x8VadwT51nLUYLrEfKKXRssiquPgjaA9Cw06Xc8UI+xrkxsVnBRID/JHj
5gjN0YU/vKzYlzDrdCWMf1MPlAH8+QQ1FSO674fyYmiRFcOu37QTb1PF7ZmpxXJZpo3vglOg0ge2
V2PffTeq0nh3VkQ3Kk0DIDoPp6JMB7e7N8Xx0Np6ajG9X7DBiIe5V1f3/7Jb1bcpVQLOhMx8Hu8C
XvAtz+22/U64vNiu3/x0e1Xx+dSK3OgsYsA2BsgRqSy2FiAbOkBzRUq/+L2T3umY7t7U6f8i5y/l
5OL0rElj06dC5I1eUwgHnQkozva2RyNNobu5w9cyW4CF+Mv925I4WzDtEiRuuMeld/cjqRJpFzoz
5sSbrtxZecybScz85fBeLWH6CKuwPi9zSBkWPErPfQZfJL/CaFUkE9uC6Xgh5vge7Kbqdt/reYIq
2TVqaprxv6ZO2zbirWws2Aah1hemoF3N+uSxNnIjnMJB7vg73rzPChj7lQw9cSO7D0dlJsjantN4
UwdKbWrTaV0V6uyYahNLPdrEZRbqB0cXrwxqgCo7PYiQpukYOTIs4bqT+f/t+K3E+vtyy+L0Y1eG
f0oyufLtQ4BoNhjx6pbam094wqzJCVJBsqTtuJs5SVvsPoFYOpUkyJv20ouWsDDqjoMCmQjzqr5P
FzaHTV1Ag3cRVX+JMZFtlLGzXCDRae1gMRGQTS9fXhqZCtHdo7+oyjUGEfH/ze2hKffp6SyA6Bwt
DFe8FGI0CCL87GyiFZ011phW2G0m56O1BzBwp2KFIVRLEr9FphRRMzeU6md8eYvMV3djo1C5dpJq
SsmC4iHbL2fmCAcfByEWBSQXy8AiFvncRwNzyP9LfSw7mP7nsR6GjLssQRmtaemMaw4WCeBaBuK/
IbiJcCzOVFrG3xGTq0BGiXE1rrLhcyE4Qkcnao5poNBKw3THWg8V4Qx50PE2L1LD8HY7oExAYwMT
3sDVTk8luM23o3SbmLT+EFzrKSIvTHr+jInHqRRLe3Up3Q32KYTHM7s8TFLkVQZhqDBqZuAe5Ghz
KEdU7N3q8qx6jooQGrD8INwOkNL+OUh8u8Wt+PKv3YI52gIGIDnIQB0DAjXa0zHO994BueA5agXo
lvPLnqi9bSYM03PqU3htmQvY51JLSTN8Eye+F+y1BFe7HPbTT6pMEAfC+XuS4l9HUO2cF/cDnrem
Sy4gZg44ozlZ3OvtRYBdHM27P7FR4jYnO2SHTVvPrk25h6XopnD81smrkRmhD218Xdvv4NPKDStO
azZ7OEJGOV76bwnh6XorsUTav8HxmA4iMB8IYZiOfLWdf8bCNfgriguRCnLxbxR3Ur9yBZ/I8kLc
+PDsghpTLmdQiG59P4dL2GVZX8pWmRDOdIXN1RmFla2Q1yG26EzAeMjvbGEBOZ9PRaxDPx5v2wIl
2J4OK0GJhEh82tbawqrKLRmzAbhay7twjOinfnSVb8T6CnvQ9jEV/lWD4ezl44VnJw2CeBqP3tfF
Nw1Uc23f6eBUHOvv/hAXCfGvKlXfLph5945I9PGyq5uG4ifrpZo1OAwkZVIDqohBZeobTCn5EM6Z
TPGrraZF5FW7ougV/fbpeZ06Ic96rKUeZMENcLkFPcEHkVIrhLmxeALwGeAWbcYCws+PUpiW5eAJ
gKYC70P+OEq7bsDuCl7dEuaffIDcnDlcvmMDxv8jTUKtSOsGEG/We1ZfM+a9l1hSzBul9p5EOpHK
3GmdEloLQPCnYo+4ZhNxTTxwciiWYkA4K3yeanoYJHm4HyKki9EyiRYu/pyfjQQWi6JMNV7laGSk
fuO1v6Sz18bI1O3LgmB5KSg0ul8yY5eCpOV4Du9lZftl7/fesNUh3JKbppI3i6Vc2lnepa5BYy3g
1JNI3ZFwAxXLC3W+MNTYerk7EYkwoR2q0h6DOq2lVScrg7B0HliccQuLbvLDEBG4XspiYjoIj70o
up7ZCubCGDwmp6vQBHttTvCAbV0dkrbBPWk9rrepbSW/MrF2naAtJw+SOrOpb1ZmymqtQhVe8ubW
ZBSbTZwPSz6UQc6TXjwoBndNN4804VUI89PZXBp0RjU0XDywrbAFcukY1b2sKYSHVvEKxs08OJL6
K66o7MDIxIOaYTjtHeBTZvELQrQZxWHWbFe2SMIOBzthJYeC9A0HekqnnII0P0boVfQ8sLRFsx9/
DpNZf/bjXKsoDmKT44lZAHg0NgmZcCez9XCdKomn82lPjLB3MVTWfnMNOi8uo2Rz6Web5UP0FqSN
zGDlsa+BECTi5VuTVWfNY0XchsLxFGF8J3qXRiJcp9i+Pup9HISz9xmE/8n+puBcRkrfL4UbyY3p
bymAsQclPQr6ID7u/hfBE5QQ7QUQRJ7sqkwG5VMEI+Ewi7JuOmc0OQhjpCeJf1SWWimc40gQu+X4
euzy8cpKXowQP0AMiOnqSpdUb57Farv9man1RJvYZrYozUloT+ldxrBCqp0vkNWkkRK+AvnxlPee
J0jj9XrwNgYO1paRjA+nkfUGEbUGWlsX5kp+loihGWtbKtfr74VQ3oQHS6vlkI18Hvd7e6wKT3Wr
yQXM7hDCYHnO46Gka4IBNeftpQFN5pUuQKAb2cKbROElNSr48f+VjJXp+wet+my+IeZtyNh3OWN1
iwSj3PW5il4Moe76+wRpfpkiPA2X7k7sedg+DkmojnWdOu7Pay9aINQfRTHkCX6/fWUmsTi3rAoh
YprodQo0uYcKumnbNmPp80X+TiaiMkHwfygbyrEJ8Aezk1IVL3Zb0UUx/jPT7UKxSkEU+P3gfhON
hTmEQg6mM9woydfWA6HYQ/jwUEa81JjekgRfKl22A46EFKDkdvuSV+sSYobGAgBU2FTV0lT5bTlh
NOAdphpfdaN2snnvCfVn+FLg+Txv8Lp9bbPjZ4xZW4fq7yxXrMZ2Ggq3B2FAD2l4KdJIQyw5VzkZ
tEc3mIVoJWyxrXyDi3419s2Gceq49OM6YVFH19wNpCig91g0Ns0EIsgYKI26MxjBXy5WMt0q+o1z
uDvGAjJR/Xa3f4LW0CchI5Xgeh77ES+FWuuEyvxQ7gcPrS8Y1az5Fta5uKsHEwH/kDNIEq/OsNIr
AKua+CapEaDYhqD7XQDGlSL5ZdTaWlXGGG4JCghU301mzmekseKLQC+S6NCFitpln0La3RUP2jnH
DTbWCDyZLSlHVZGq6h6LF1Dulj+G7HzifwZ1wutEf42bFvHYysoq+YPUOG5f6epnYzLBSV89HRtL
a5bclYggIbG0MoprRjf3UI752EqLhGfKdPeMMwwLcoI/A7EaOpTfZKJbtKfK47VF381wsCBeMMa0
UnnS09pLeowfxqRf50vpeaK67oo0moiAgD0u/5kxTVKfyGQjjc4X1ad6jlA+g38gSDGGN7eq7MlM
hG14Hp4jLdhKv2Fq8dhU0ciBmNHVIKhvN8TXaEznqYuakAXP25oDw8xRwzh3mDCt0KuJIL+hX+B7
0h9Nj/D7eIj/TRBXnuQWad29QXXrO6lg3bChXaVbAEis86Lw4d0uKiTxJv6HZLwgt6L5yR6w/xXe
K1a5gC322re/A7MBEcSdfObOvw2rWmhkQ+4Q7JepYJgcrPTNmf4EE344pRwfYeMDfTzk5rX/aUrO
uSH2GcuxLBwyfJTe67woUp6akrhjjWjQGQ9Y8Z5fl2Ak6uoO6qmox19ow0vN4FBtsYFE+d2RQj8l
NgCoK7EqeC6BZndA17NpdCYL5KuwNvxsIBpOduSSB1Kxh6CaGKnBPNFx3xr+xS55NadJhQfCFKx7
OveGL4D9wqRzaJR78TsvgUE0SuwCunm4dftblwwx/T9EPLt2+elg06DTKaVE8E+vBlpCcUw/0PGb
QMVprgbeBTEdVMfnVY3S+QPOVOoqDxrCoHMrk7lLU2tjLF7CTPf8MqsKmmWGuEpXdNBNQFGCzlXm
xJ14XpTGRmfH3//HU+vtM2A7DZFS4CZhR4prs/oH4shd5GrOnNikO5ZEDUjUKcruwEkmJx3OdkRX
Dlh6o3epSE9ygMk1S4QITHKqxhwUUvO9yWYEEhYXkbNzC08caleoK4CL7D5C/2/Y6GRpmK1FADdK
Tjm9LyqCcmOVacl4kc050EjZTXeZ5ISohF5a2HXCBgyaFM50SSe3sO5UYd+Tp00qsf1rqCqJ6uYn
9TdiIig/oDWRmHZgRjrZ99A7V7KEWkfoiOQAEAZeHgHCdxEEpqrnMGuDBuSmFgKD23GU9VxkPKTI
DG8P9BDF8nBwVwf7zqRp15RVhwb0SWyon7wXOAc0oRmsnIEeO7wopWZ6xSVuykuLOZfiBnvGJz93
E6rvxu+/JH8Bz3ZjD00/vIzl6G2xgMXsNS9UmJ6MUNQntksEg6rTVIkrc3pyjTftXzW9rON74hqP
l25VKAe5qoy8ijNi86D7JTSqY9sYlV2nLl+aogKqyWmB9n0MJosd22Ecj5HSN120g+5CM35/lV0F
xCxExp4pS9lgi+1TfNqYSHesmavDuWPMYo+5G3nPk/xU0Xt1nWUm5N+Uvi4g2pLgNdyAGib/eo2D
wIrJxx72I4UkohhjKpWlDhq7wm6pm08jZVX9eDmUMP3mqpdhyOjOC4zMPF4VLdL2Gvrkm/De83rz
D1hS+A45rFH9xM0hD7UUodNY6AAmdFPoJg5JKj45Lv/R5rsxSjeP0J8yXVqHuf3nwv44Uh34Ih7j
d9sZwBvNmSi2YWVskYvZhJXpXSCsei+vw0VkFNwLQyd0KXXV4aOiH3kGdafvmDf9Ws4DdA7boD3L
9dfZIcmOUxmfdVfJdE4EY5+ARuDhenEo5vzmx+c6pArKK1F6TaOsX3pg8z2IsSrHaokpbomDMrdW
qIHobTdTLukYIws3W/Mav1f9yvFT8zi9BMrjPxcgZsWQ1kQRMueDxRgQ/kQ3XrJBBSQ8McKNUpQa
jFqSQJ0EQz0H6tq0VH8ZBiOlLTEJpypR7fKFjgHCeRFZR4oG5T7t/9aSMhINZp6gNjxob7BN9J00
u3tJZ7cW3qeQwZg1qpfB/0fGgVP3UqDxCPxoQoXUIYiIwrWznC6EpHU7UlnB9oMNzx806+lAGyTJ
cDy+GcD2Lc4X1rWMaRXBXMXj2CqdUjAR340LgyjJ/Fc6LYsGGcEbJgJAeqmKT9nl4F141r6NwnAF
4mPTYEGi4WqYUBuHUvTvf1ks+biTsNOFitLdJ8lDYOAe2XdaEYXK6uh8HkMjluO0lHog7rCOxp4J
n84g+Iz4huqSnwEPhLcZTGCiqgDuB5bYWbvr9ypf0BPsszmN5SLB0qwVeb3nVLNFEVH02OTzIufP
GGROdv0n6coszt0aTbnGpjldQC7w7iBzSD5Q0uji/ANd/GiIuix9MSmoYVWMreOhcBJXB2w7MreP
T4IBs9B1XFA8vH1XdGMuCVWGEZo6ucNLnb6qOQToM7A7+VH98ORjyKawDIaJUKBFoshGhGyfNN5i
7ZR7pocVDquSIyi0PqBFLkWOU3CVts4GC6rV54GJoCn6ooIXx9rCwNpjgJMgn/MErkXrbVNgK6ZL
Gqy82Df8Vt8Eanz1qHopevgtFkwdUV6MQ3Mqq4e4tDmLUBZtw0iOA7XBwR7c0SuTSI93ITxiydQv
wIpuP1J0GP22QRtCSfnLoIUuomWzhbgEUymZ00SuE2YqlzmAjShQf1I5ONR8g840A56ZcZxlZX9r
+85Lvdwkj72rxtheO08f8BsfdWuO9xWgZjoSlZJll7Ur8QCmUz2VRXUcHC4jdpOmP4w8rZ4VYvux
EYHyc9lXXCbBrmLs7AeI3tg9ntHhk6bgC1EDdC/AN5iyfeIKSNaUMituvYdQ5DycZUsScBfjsYGf
eq4d4mq6XbBVAEf0CVlK4mgFizGQD9oSbKnYOn1DKRvOnDtfic1g7tnGvjDbudm+xmuddcmFK2Hx
7CNTJT7u014YyRoVRymhl6U+j42tqSOyxd4MqYDKcMHk2B08/pCG82dI1JxpdBADcouSlKfTMILI
QYngwJSwy70gDWaa9zxVX64ElCw20T6awmtKsTyY8lNDvKPUneYvBlvoP76KIZGU30Ld6hofQLyo
MJ/aZud4Aqa2FTigBCaP5UDtB5vkeDjgmrsz+UJEXdGKAbB3EhCz0oXjDp/9etmG38lP37fdBqRn
QK0ujO1VjxUA0tFdu05bdPPTd8K7wiqi1kwxHnUic4A2yXxW9Gwi8g2Z0/ZVHCFhuBP9S1xt04Jd
Csb7a2id6nAWQ0HrCyHOWIFY0V6ubvLLt/zge1cDjm7DOxsMq9aHHKayeSlHnfKo571iTrXtrlDv
k+7fPgFhNrPcy5wLDQ5cw1K7BsJPE3SDF0WFBDRku4hf599cEE1DlxCqHpbV5yhHGfLV2xZ3/T6a
YgvX60cOCpitH/hD0rS/TqQRy5reSgvsSgjj5mXYCFt4xkGQ60Jvp9Hz3Yc4DullmIZxnKuUbgpM
VXbNfsql61493CRUd/uYyq5cJkLBK+zNGpsJWdzkRzfrjI/EPekTU2LjVqkOdnrKBTNvmGXJpgfl
Ynl8xU40JKjQ5tjf5g5tKnlsgiAvSIQqcMK+OeHnr0HBjO143JKlUQM7SJRV8v+glr2xqG48Tqve
Rn5l4WfZiY0sC6v1xBRTMxmDF5vzYNquR2fYSxIVqHFTyXK4BeIobz70Bju3j4GpbzojiOsUQ++Q
b6tX69GuUE4t0rQZVXVkaD9va5egUZp6sbMo5UJlEI3VmiO2poo397/IBdf1926p0YTOvKIi09yi
092NMjCjUe+ZGKl+YMP5NEAI7yrZNLMYX5pzRW60dFmiZRNWNymWKAd2m1evJ3NZ28jzZX6J1JOn
8L0TMvX3S6wBVTb7wCJ/jINkCfrFb0YWP3o5/RM6F1+7KQcLzrPViOa92paDq5la4z57Lo0YFk6g
wLhvuuvwWq1aXP6khvUO4q0Aj8slv04IDMzfilExocMU/EWRczAeNW4KkWo0/GcNfsMdvaKTU9oR
lQAC6PBkpHna0bjLXB+Hu2kns05k2a1bmEXbo81c7PIKhFd5CzUAi07knRfdnVgzW0P0HNbCIRmv
o6J4Nd4/61Lh70x+Uo/4QYqVZnxg6iGRI8jdBZvr3csszzI4mZV5SCn/L305n9uwscWGIq5Q3O9a
1BvwDTDK/tcvJ3xMg+nPSGgl4flWvdSbb9nLE8UwGZJq0uTmhgYp4fvsAP0V9w/2+hCh10tCMttR
JkLTFQpHU9moSsWdPg/aRy27itqRVdgDYgUWChofotKnVrKOUmbK1z+9GVT8ZY5eEnwzhZc32E0B
ggEoDfIuDPt24TC9WvL/TRiQQ0oPFRXHVG1IMejfatxmj8vBBUHCVMdDpx/B+LcOMvAu88o+jsQQ
4+m5L8mNUbh0Ao1OuzsdrkpDHLG8/nxVkvaRSEYcA0OLEvHRifdYmNEsKZvh04ynEsX2sLJLv3oL
GCFDKh9j7ounX4rBvZqYjnJXCDNquMy0UDZD+t0sRkURPGHZGjXkahLsNuxxB+mDahaOwcyPmjBt
Rnw9FmYeTWuLV+tH6XCFZiK/rJD1p9KSPDtAa2OrTuISgCvOzgxVaS/HULwmKBRxKzpoZDKnMNa0
FPdniQjQ8nrsXMC/rA7CDSI4yTq10p8IbRIMVAyIcPbDTXkX+5/4h+T27pZiGL0O2/ysE3eol40a
Y0waDavI5+ccziP4KD0FkxRz/DSwlAbYhGqwqYMuePVv3nUaJtSdGQzTc21f6HrGzURU4E8y7Szo
Or4LZ4+uJ56rtIWoGKeWPo1oK+P/+rK2wPataeMaGh0H/QZpAZncTOkCl+qoy2+yaap5LUqA6Hfx
c6WqBYUEY0CLbY9AUFkqBGPJ4kGhz7YV/7Pra/cfndJYjaYBpctw/6VOh7Af+ju8bu3mQ2fi+aHL
Clrhty3iLHgtTONrg4NiLkEwbsHIXzNlPyIJZ/u65h7SYZaeUKTmj+SwYjPMZZ7SEmb2REEBEckL
orYabnCH+gkBwwPavzXYNzfCDm3qwsA/cdnwTUcJol7iLj8LZokMyQc0dFuigbV+jUd9qDh4BrZP
qrRsuQYUS0ajFqV5gVwLDRsUwoFVXFrGnirdYjTgTTuNXfqZ4aq2pVZLKh87TTd6EVDHShEf5Lyt
1O5xchadojVREFMWzLqgf89Mvo+3GvuRBpLB9oZsYrUkUcia9lowYmp/5mFQXroa1FJ+DAXT3rDB
NKuKoYtegNDOVW6VVx7O9x/91TFlrrGU83GSxtAc9uqwfuObLh+V0/A/J9HZrKTlYXwECfInki6y
wKFWnWHjHvf3+At31bur+8ovpUZc9DRIj7oH7SxG5obBGnqnlBzegvyngzmk0skCEsCiUt9o76NJ
xCMaLSzIDFx14jTfNtBdI3ZibyYdiQ+t4dacKfVM/hIUUqus+nh2T2N1DKA5dzz2ajQTSu6jS0ov
im+F9BOjUl15NnIOH6rqR4SCbgOz1DgxHt7f2PzA2mc71Z+M3XFRHrpmF49rvx3xuyMmV0tNIhpx
NAQnXNva1XR8L8xxu43h1R9YVNRJAJjohy1qHMw2SM79+J70wJXxU+mRL7c/gVKzdFpjMniKpLnL
leO3ISBKk1b4lHUKOgQXQHTu9dEwZVuZkZkNpBuKpVimvcWlIDFqydUPgthWB3aPfhLNMbn7dBv6
pHLJexiRtouWeavQviaF9ibfUfKpNiT9EIop0LNY7LIYd6JDPas6LuwM7h6F2c22tNSwXNZZH6A2
zJcKP18kurTiZsWazOKRlbqdS2eRu1kuMLJFy4YwD99aNbMq8aCMMMpe5lEL/G1CNgWhX6UFIvKG
+Ehk9qxPXvMydBWb+5T0LG0PPtbpQvvL+3fvb81whWcT3CcLLHcckq7kF04tXO0XYCWYCe9Z+KDd
eR200bG5FnzCjHQ66BGdQtho3NtgbJadi8QsiMnwG6BLIm8WCeSZaDiRTEvnXoDyE73WAZY4SKAw
bV2f0FFXOX2iHT7jQV70OoFDNtYyYY2u35oxeSctGVd7/mTykktaspeN51AzNh0e0LgMKR3Bpp46
6cZqxsDIiJoO7qRZReHpQ19Y8ggSEY7yhAjEQihLCp7wtpPkIF0wEH9ibfKs3RTjP6AMgxd0LsH+
BXfCxmwDl5XOAFJaEtZ6T46OJJViug5oJjfJSxHeAVySFgEkjOyWVSvHpj1TNh2xGBgXn9wLrKaP
Jq3LUzteCwsOCvuINpdVNLkNqEZYBJExkj1fHATykPSrsDc31WG68Gk4eiytZ4yBJGC9CdmWuJJK
s2MTzt/OgD/UNdc1xYvIHDH1hQk9GHFw7jl05ywU58rQnLWiH1sXIzaj2H3IS5E3jjcozeJlUItz
vwXefiQLx16m+ErpHWhymVQlJ9L4s9veqEQnOrzH9KPeX6XOH+D3LMydpLeDei8UPLvVKpwKCUKz
StXbeyIGvqO86ovCZpTUKKelBa7XZHRNdRNtVFF3MHMh9NQ5ezpZw1iy3RbxbXM57Kx9cbu2eAm/
sJpRWqW6ijHgKMy8QU7G3efhOwFrNsNLrJWVXawqJMyzglX/N3I0wjNG0pQi/bKw/W1YfJTof/mK
fKUCj5btOINL7fKk2zS8M0OYwTIRsiaaRHrV7rp7trdvv0qPvPysyZanBBn/2ZyMOClrPLUeJNBR
11tBcBn16Ojg7vbKhTC1+L6N+19ozX2RdMRfhn1xNgNJ2qQH5UFDSgRnqYlTevOl/uFikOoWI6+3
J1geY3dycoNoE6dBEY4dcX7fN2nTp1Fhbb09tbsDF3ds71twFE1gBAxCqwcCwNYYb+VkTOPpgHuW
SCDzIemwIksZPSwJ4877xjD1DVTTLKU6MHXiZHOHF17dFQJ0Qwo87Kp2irhNw1LNobmnjcroEsNC
9VQsMr5MGSV1ZR2j7v3DIQoJeOh9YupSGny14lslmbLOMP9vbabhxwbgE4X/G2kaPwpvW///bMHF
hpheWP00D+ZI52vM1H3JabZhS6Sr+OWjn6LEcYe6WQtrUDqkS9fpwaAx1CiR+hJYlXfWMtPq+Dq5
TT9UIZnsneEUPiChUVeOR+v99PYcvjWN6jh8d09Mn7DtfSaiM4fbAjfzP4I/V+Xu/jpDDShdvr6S
V96GMBXEoHKhFmDu3H7RiGQLVkfvssv32pBfDtmdLvJhIHyl+2CDSRTCkjfPrbo8zIO9GGbRW+Z5
j5onKJUlJ9iV3kTc7K4D3rFh3Hpvg4i7JzcaFD2egFYSvVoNsc+JMnVrXzvgqPANM9O3GCWnUU0C
W2ug4SMgRyioQW+osfKabpwJldOotO1URkjoaXSWhjZNCy45yMEaGvCvBZdbuLWdQRNMjOxs0i/W
mQf8Nye54v4fzdUAsWZb0wLmUzjOG6EFgQR7nvZvLvSIkgmPd1rmzNyCn4yeNY1qp+eBtD0rMHaE
1W+PVHb6KndjuR0CMNZ4PyF+JJdkkTwMQ55VIommz4/L+PqSW3wsR/zGghMU91avXJr8KIFKmP3i
J/BtkMGLgWa7nITUEjMjYNw1lzu2Q3pjVeh6N9ju/rkGq5FROliOvMbUl6GxUIM2TmXJc29gYpQF
BO+GmCGmAO1+jMKgkQPCsBaNvveH2FPeuMdtSOnJG/8OXOOgsUCGA4a93MSBlls9i3PQWONuDXAL
eShywSe3KUslnUyo/CrQYns7JI93ujlsL/a4lQ9nHtF3Hp0IRt2t7D53U1jTh7sRt1QvSHRyj7P3
YfG+subOCMVfJoPzgrVS03WGq3WGnTEvJVXiSI0we5SLMFwdDoFNpS2HjA6UguMQtDTIdKemAqs9
LOLq6TckcQgYyxGSyAaKG3i32q1EgciclTOyM53yNk2OeEYEkp9FYdXSDevam6vy0OrtBD7pUYk4
Jfi29cFausn0rxMwu3IeDV8c6wqUEipO9aKqgaxZvH9+MjATMuuDE30RDCEyFJ1bmktGaOhUHNN4
7p273XS7E2xzEs459zEwOwVCPOyXdZccyE/k2MqhZW1zb2yL10elw+DPovLiaXy6zjwx4GPqeiI4
OVeZaY8204p279oWxhvgr1F6vb3mDDOlDX9jVOqWTBkq3iXXvbibCrmn4eGNhR/9py8YG2URrauQ
Mz5D0RaS/Su4g/eyzxED5Z+AqydXsPxBGTQ/Mc7pRo7tEV5kTa4v1+bJa4rUqjoDO8vvUcUcw2aX
fN8WIoi65Zs7N0K5+ncTK5VSZzCAcCzwa52gBBEHvfktuc5M2+6MgiK58MvdZgXn+TvFYlbPq4CI
x3iDhqQbl+YLvyyz1n+CXO2JVzlFZyR0J+8WWWO9uFj7CqfImSRBOIBSj0uENmXzvBhfbsY8ggq7
lKar3DDbwHuk40YORiWczJpHPBBz5PhN1Sc8ZLdFvD0qbjr4//CfJD0KeqCIccQtzjI/PfglYWEu
TjSFmR+bzHanpSxj9yESpQPZOurmdRMxt0EDP73SNEUTxoCXdrH3PfIqjgJMKWpwuKa+lwcSkrrZ
fPuWg9lFnOx5lRT1RgJMfnY67rv+WouYEAcsFueKyLsS4LjVhIU8STATuDVz5ZuN368cL85Yz0Dg
kMlEGI3bK7D6nrdKve/Z54yHWRj6T4xxSmLULgrcXSKTehcnlQVQfhdLV+8FjKRSkhMRdqOZ7u88
cXEokIGypw5z1NEoZK/Rj9J+RlwyXBT6v0iU4WK2+1lccsO1mPlhxaxTOHnqa1DEbyL2pm4zRlWJ
HoqjUo5pEBY+x6mHjMxnRFAn+eB1cSldRS2sRZ0H5QiufXOZC0JcCKiv+pWwpMMyjQbQr0Kc89ez
vSD7qBucIxwZJCdHqqCRaGZdIf9tWceF2VoJJRYVCbpEW9s/mtiHzBmjHJ1tUDuZczpgxkOUKs42
K4PFTPpqyB77vphtYHjM8Ek4BVVV9I/XA9sAGWP4O2qfJtHTHP0G7xfOd6sTx2x2cBdEfuBfuw1u
s0Q5UPpPGVDbhlWOyUfPkhMDtLVk2/N1zIM/1Y14RhP/NhlrH6WXSrnX9bSyeNxxKvTdg/qnhWTz
QNt6yi1ZDmo9fy81pB0C7Zf5ya36hO1Cb6jGiWP3bOB9WCMUAMbZ3Pp8xja2CB4VYA4HedpXvc4D
c1pmodLSYkZYri7Mdtc+8p0c7tBHx6gJaHWAo/2KqfmuqCFnsZazrF+vB4GdKQx4HLxX4HgWC7/v
SbpV0LBrCY4Mf5EKl1bK02kH/7FNni77VvRjiTnE4NlMbQcHUnsxpsJrpwsw4be7WsljMyDxO+5l
Sv/lPLSN9IuZRhXzlTibNpUc9JRch1nByr72USFW2l1SzKL0+Uqa98DT3pMN5MtkNcLA/XjdxVcC
ikhWuBHo6j+inuzCFqt8pRMbd+tLYwmlToSxPVmvUYzhS5YjJmOJvfvyvlFMnI8lhwyYdHUY7qX3
WR8Xh9qQSOmcVHVCesdMgeRKppU0jbOfPdQh5mj6bhVMUIqbKvQUzdsKJzdzl3/bnDwnPK5VO5mg
BV/2gK946rPLbvywX4zWiLxUpxVq6izntVi9B5t9ZkPtsWoYhTSRL9b6K4hyycxRZuftb8Ba2UKX
FR4Yxz7+F+vG9W4wyIgnHN06R16CIWOf+G+sBrf/SgtE9tzDiloXpmfJQnCOWsBe7wl2YKL3fg5M
z2hsP20IsW6Q4jzPCNyTs0H1dxu1Dj/Ge7naoO7AP50+hDRPQYq6vAKjtFKWUzjku9hYOiMWAF1/
xfmlXmpAXAxIaOzSvsuLh7HU40OiSF/LxLv7lSbgTEt+Nk9vttiv56kvnCmm2aSYjo74e/2d9d+t
4qtETzqnBPk5WH5ZdeKv76dRNFBMPoFykLPq0+DlxYvpuah1R6JndM7GoPrXw6QQm/L2IQN9uyPB
3txcQvbB6gav8/ovP2TjvK/JxEDbDiKRyeXsw3UPKTsxeK0Wj5JWfhGwGf0dcn/hEMdETjjvx87H
bmJNq9BWMpmSoWsUZFT3Gt3XuFUT3QbI1VX4P3/zPY1/kCY4ydQxLgPtu1wWfeKlT2wEnhhC8VsC
OennzpHrSg9BHue4vp7jQ3HPZVVoquZVpym1ZS9Lp4jS96Mql8jjpGeSWKmkv8Zypj99Q8tNeI7e
RRMVPovMTR2ff53Wd0+/pEHxEEEhsFrnvdw4xw7o80Qe5Pv61GxeTNC4DHUBcvJj1D4cB5Wa6qTh
6T29r9pbdf586ZAzCWY4X0ANMtgFrJYdG2y8SXtmRaFCmbRuN4Fe0Vd+WUXPKyYyLl1EOX+dmj4u
44vBlkJ3EXKtPQERIlGB+l6hhzOa5x9W/0GETvb1QxZ9iVVgSbzFKWJdBwISDG4OfuZKLT/9THDc
KXyhEBeBICDKgTdGB4hZrGJK7s9awADVNlltzlhm3cqMMh2Tl3/eJyi51yvg1M6btG0ojhzsP2cd
/VuTDfrnwnMNk2qdJq9vb88N7tI/yS2gbO576RPqmS5TNlc4Z3rIDXlkIa0D0tPvlp1cXDgG0XYW
ija6d2ZHzR360F7IHuVderXLtyMVU0VE7aPcmAbZU0QbJGFDrD6dV1qctFV1LtPqdTXXg0hyRcGz
tQTiScRjCxDOd8IIOX60hjh9j1oJohAmk6NTBKk6CKeNwrM9XVO3WJMUq5gBJG7a5gIubAf5MXdG
bbMpltV9P/Dp3TM1yzb/wW8znHVfSK19kqgJ696Wuqm5nAbdyOG4dm0TFm4/5Hq+BZJZ0Xhfe/99
reN+buMfYmQJSQ1lgkEN3hurxc05++IUsACXuvNWt5yKO9ffy1xIB0Xgos500IKbQr9HvGbyL/2M
iPpcNJ86eZKsiHFh3BkF0tS2tMOxFFsR9S16rXJmt78gZyK4sO3qlL+MLfyxqYvDq5hhKL8aKzuZ
sYtdMEUiPjrbFUxEya+46/k1mF9w7V8LOav3dSpVruLWBvRm0kVwYdN22f1mFlKnDLoMOqazhWrk
MirucAWnqOzdD4/7uQQ4/fk8S9fTkJvV3tbihxulaySQCi3YCQZofJlUxlybiF5E3otQq3YcfK5j
hFy67gZEwcAEO39G2bm+jtcj5u8sITiwyORvk8TzyP6N6HpMyNDhgjj6Hkx0ysivvqfTIDrCxBgC
48pqH0mZbBvdn1mTda5YHOCG2qM64YGGHaQEdU4nMUSTfhQqlYyDK/YoaqPkGARtY/tZEtAynlJb
Zgp5Cgso9B3FEgkJ0FbIXXtgr/vzA/raQ9QJppo4wx+a63DOQsZNIHwGssHMhNYn6mjR4fK0zo4z
dDZU87ldi6GLNYILok+GoI3wan6P1yUHADDh7fj3TBITc1G4QFhPWtN03F+T7ZJ/Sc5QakvtDsLm
1HFz1iv7LZwQV+l5B+yghCH1G9B2sOSLuosL6kJr3gR7s/FOwCBbMcLbQYMPlUuUhjhuCShE8D3W
8/bYI8OSjQzVYECXYMqdFh06Cyj4UIgAlMkfxbRG28rWxP7r4irU8J7/LvmZiUesatN/+GvP9Zkf
imYcyJ2H+E2gWHsH6or222N1PY5v7I0GSc3Wk/hai2QYNoSYnPa0h1Sm0XsPClTiz8NQYrknjeGI
dWwMpxS5EWccRXLbAX57qALcdpYLudH4eBi4DnpVpa9BeWfrYz/uAlHGPp2+Xk1gIIkB5wSiG0WC
B2mVXlq8msVTKBBJy5nEIeWEbft4uGw5BGyK07EXaTpq7eQM0LqQTF2xFJf2SQSP0jqppMgK7izH
RDhK7gTLwT8krpxHmMmW+CIV9q5EZUr/qugZvyWz2DS6citqVRtmizQfXopF+VR4MLY1Ux2TASln
ggmxgwiK8XG1FUO/oHW0I5N/hvAQfND05bcYMjCewwROiGcXbfoUXIQ88X0PsnAy1FAlPU7ytUWq
1KhTlwRV+s2uICBrixrwIVEsl/2+Xl0zw29A9ddF8Eg6xCFwXdDI//zPHaOLa7QcPY7AYtSStyFI
/uw/ABhY0ABF0kiRdgkK2nw0mrDsmoxR5Npj6SOzV29bQok6JstgHBYpbCEB5zrWEaTXi8HikVzu
YrXGyYAIuMtQoC7BUF91/ACHKjolftpPR07YP/dtZHBH/nGW3/3MpuDc9iVLEDYueIKl6SiD8ged
q05GMWDvPjt8tJy6ck75ECaLf06+DqSdxOHyMy8H1JRybi81rrW/7GsOUA7o8YlxlyQ7ml0uYt5p
ouLGQ5AEElCXkJtkDzBjajJHjvHUBA5QzSrp1gDHH/ot/3T15AS0l0/q3hAy0UvyxT8eocXWEF7v
os73RQAjy5FoQfFMKqlzCn2q7cJu6qwYiSEFi4KNpudcGX0J7Q+nNIMVxLJaTR8BM+HctQ1Yu3Kd
lbI2D33UA5Xj++5begakzsDs4crR31kSMXJ3Kl+ZwtB8llB58rQTNBjDrsKh2L05/O9qbnDF80Wu
IdxsiinNEpHB8DM7WI1+I+Xnxwlx+Fk2nuMhYsAojuZgMHmGtJaKz49iIOCQ4pqW5jey0EzwkjL6
8gHI79y3fQufgF0DNyrwBub2S/x5RZSkeMIyli1ofVGwgaO3WH6dL4O/ujVFknMD2t4bH85rY1jz
zQ287+oFyuepLK+fOSZyX+RMc+UMlJbjcsPVKTqisdce6Cf3NtwGcyM9+pX0TMPGTXTHNe+OR3VS
8uQQEym92AYttL9MLEIMvmRE1zuDCfj07EevIsQii57CTViXygHykcxwCJIqcDCtfjYJ8tW6ef5r
J+DdFI1UsOVVDtpAKGCoDEaYFIiCIkmrsxrvG2nB+Yig4nKZ6CnTszr3kACFyPpmVzd1WADsTI++
ISbptlzvO9OHwkFxIBlIKIE0UYddHWtNSNSz3CP64E4qlrapdJJ3gkaBNE3vBENZdbgwMSmLtovL
jCZZPe57LCuw26k40g5JOD7u3xJOCbv354bU1zEozg61edYiYzQorXtrQsax7ZsJJRGRt/mCQ+qf
7w2AgXgEkMgagv9NE5ZZWpIfVltPViLB3cuheaOE1f1Hz+8F7wj00OhwF9fBhzZlX+KU7D0Ytv8k
hHg6c98r5YfFl3CmRkABN5Avh5ZKBzW2MUWFcZgQJwLYwh097JiNKan15IZP7ysPRfGdJnHhdxF+
ef8EUYAhldDd+jHFCEpVaRuuGTE6EqaY7uc2Cj6fOzN1Z/HM/coEQslUkjd46+y4gimndyiqctRD
P83KWMUoQHaDp0AiaMBihjtisEXaxCToTNJSFj5Kgexu7v6Os5oXT5N6RGpfesOVVEsckHw6IVWd
Zl2PillaDMnafpEnsEtLJfH+sZMD9cbkCSAbcj1DbuSn/pDHaOgiikhIskfYhvrZd90O9UOn8CnX
o7b6dcZ2fkpoiU/OyS4zhzwKqTHpoULYv55e1/Q72vIZT4MZ9OTcdNDDT7KW9SzA9rmGlVJS0/2Y
BpjCb3LzVttfiGMlUUNz8FH/5qtY532akI02jDpQ364xXMVkuVNGMHuNBauQPNZbOCPPPB51aQ1K
CJ4R3b9TUZusY2htkNTJVlnIucob1BbCjV99RwuLKnu6Ci3Q8UvtMP1E187pemWiRCYaLhr6ssae
g9IE111Dtgzbm1zZQor+qWnILAb+61Z/MBt/Q84rydn6B2tlccvtMOZlwa0cB4LshVLNobXeC0P5
vATa6rrt7e8wlDX2dg4/AknXlsYQS0QxsXbv38tK2W1bhzGgvuwJuKQF3c9I8yoUOe4XxSFCSVJo
pp+dDxBN21EAmsMsSTMdsfqKHlwkuiSbPgG5ZTOTCuvHKG87IMvQIr1ZTDL9KiGF7Xp1vD2YZagX
TnR7ZMyWg0UO1UDTgB4wzuKLDzUt3ViV7RhPgBzFkgYKlBH9lh8Z/4Q1aWw8NtV/68dSlV0HJa6Y
PhI7etKOfhf462+BWsxlob/R28LfnLv/QntYY8xMEnOpAHHKsv0lfwP3QodwEm+Ck86AY2XZaw21
jNAARdoy7Z5js9DaVg2dTsmDzeRHFHUNGNdWdedS49vN5cTEUpFSf0e/TRmNAkEBMo8hE5xa1cQB
fX0uR4O60o5xv2zU74AuIkX1rCJV3EQQdYJy0CLNAt/3xP5n/cT7OriwpuaVlPiUxLdPcqHLDR1R
hAfj6sw2NH55YX1tidwmTCQM5Jega+NHSZR7NmeZL3MkVR8vxF6u+BAjwkflIf2k49d8zVMvC/LV
qjh7AuGFTK9bovE5txLnGAKC6NjJsw9ldg9sD+7rGRijKJW7e0wv1O28Z7vlHD6i2EJDA8eE9C1W
EUZr1sq5dDZw0lnOVL7AbsBGqvsrfpSEqEwzZrrAv7Q/fOKn+XhYsYL2RAYyQiKdO8VTPcbkooZM
dNk/I8hTTi9DvFaB8O6U6KfY9XeE/HA2ECSIpbtJXNIp8K1J98+OsTvap/Pmm/fEx+56mv8JBQpo
NyT5ZBEx/lEvFckkXsgFnfRlSZB6K6Z2XTE5mI7IP896hvkuF8JXTZ0/Fov3o/9AGO8YKcXsHYB2
R1Nn/1EqAnYC+4evakW0HiXTnISQuqkVJyIIQHJ1ho93d7osXB63mmGuwtM1GGPIYDoo25ZJ3kRZ
qq44MiUSKyb3yFzV59d0WTnp0Gb/3Wb3yIj03hOR506g9epMem0XZHj1HvZqb5+1r1qsn21Kdi7h
5gOB8xSoGlZptX9NWAji4Xc8lZbRanob/2vjQmFd6Nz0+L/BO5LEDXbDTCJUX7LBgC+KgCVXiDIH
2gRdUdcAz6bcMgUOCMKNF+Kl7MPc0096qPFsHZgchmTBHsh0g0jCjkcc4t2W8IqdhVLwiATSkcAx
rx20NXtqYAoGFCevlEyyQgi7lle0QhnYo7NlfW63uGrmXb7dPgFe2ueQnEvFlsS2qsMPe7R64GFz
gc1EFSeHmyikXhHFVCjt0NVStRpHwuKAk15QKvhZ/srjKfhe6IuQQBwVza5IwLMx43Z9VdP5Inbs
1CUmdCf6iRydhN3VccNcUpl+gEJXgXdBQ8vCsNN32ri4ISvI8J0W2fAJoH6Li3x1IqHOCjJISdAK
1tlP+mASCXMhHgKJozCc16SBgY8KxcYMuiJKRhZrCNlufatvWh44OdJnFCBYSp7LiKgixFCxfjyA
uMPWrkwW37vKWxQsSDijLqqgUll0gc64pyG0p3jJDxqpte60EzQZSz+2Vc3KDMPMD+lXf1aBEKAO
6br6N7pyXhosIJNO+e/F3CGPIBuHSB6n6DuPFQatuQD1LvgAOt4V7gsjLjE3/r+CfwIqssAcfv+I
CtVjyMzqYHCbFjEdvT69IdHYGLRvkAoZOz8oZ60egWaNIYRCb/H0KmqO3rNZd8O5V0qAO7ULjoIV
F4Sq+LUXIRx8IUGDZfxEO9IPnh9IZ7MzrQf9hwc1z6KgnUUjimbJGdtJoABfgsGOKmta1PEUhQyk
tIfcRzxhxYBVZhvbkRqu1WHd0QdTL8cwCx8jLLSq8UKuqxxS3tP0im+/RM6S7r+i2Fx5wRd/6INQ
zFL/CrSCjDFm8/CAOw3o4eRg82dzpitJIyBo+OcuRSeeCn2Oj5r2PXFJCwDulYHB7EW92hyDHLcJ
7HzUcHyQAgLzzFh1C78TslUFCEnROPhFqu3Q1zeCVgdkKv/k3NNd7XVoMTuEsziP9wFua/6HmbJZ
YjJnImYlcAIv5xbeyuyv0tIskwkoxInM3KFaX+E2Zan2E/mebLyAdCcs85rNOYxgbILduPY9XGxt
kpBHVFl6LkaakO8ueri8iwDx8yBNfs912WDv1srrjWb7J3lwBcxB4tzG1G2bSTexjuA3Bx0gQRY8
R8JzCVBg2B+n4Hu8RSlp+4u4f8zM7ml0pXCPN8K4GrAcI95q2pmYA2ZaZCl1KQ0VGrjgVLDAbREB
FKmKTmqurYX1aSn2ZGwPm9uZb5KfFIwRA4+S+TLEDJSqpMismSPoiHvY+4nXxGy4S21u+exENKNM
0l0+6YenQ8GE+xPnZC3abERkVaC8P5We90smsAgvZGBbmyrOXY4oXMf8WiFNi3NwsvVQcvyj/1t1
tcw0aWh1s0L2PwEUQtstcd7DfS56auQhZ+AbefYKiYajhDJmZglt6QzNzKSlmF68QYiTKuBZlU6K
ggRC29W1qzNe1GFzKkFXCpqC6fI8JhOeHfozFv+DeH0/35GdKiqB/f8eqo/ciQ02lWxnrdZtewjP
KoWqNySXQXfhHWE7g4Saprq+RunxaRic2J/pC6nrEV+6aM0Yn4oQK8OstyhVDG9r6sR0dFfXBK9L
DRfUfGmhniua2JAp0m5+yvQubOROfM7v9oyg3kGGbjXzSD3AbzHLPB+aOab/18H7PhXyz48wajD0
qGN/6P4sndTuXZX/Xmzh4hS61q/vQTCeZF8MzVEQXuZ5VHq6SqF/dPgpDiyL4uk5cbk64dM3MQpr
nI1XN/kq+VDcLRtKFG0+2oC9bLhCDjUMYDT7UhcWUpFR4nyDOUhrIsnPYFR/MQ6oIYDc+nfjV4yn
TXkc0zDDDBZKMHss6UpfzFF/MV00cn0vVvYY/w7f8zXI6AbbZj9MmTVTG+xTWe8l7FZibuPcGbjl
29oSxfWJeCl0fHvK61ZYpIuk+Lw5dIDAhHTSVNaSu9vJ1zaEU2gAyGm1A9Ibl4iElp8f2We5PNSl
Rl6jcjbKyxF6Y9qNHWCfj8etq3X4dczRymr87k0kGNIGNXXkkEoX01jW0XH/Jrb6jxKLAVpzZqgI
lImmo8aQrZLHylXew+qN0hy86FbQVpZlDH4Q4ttAPCNMVShFRoTEeec55AAi54PiqFsfs04P9YEF
z8Y+4PNp3wZ5IOnwY0UeFxwMXzOeXbowx0AEhXxVbE/2R4K1hXg7UvaAQlrUaHdBBJ2OHOv146eV
nhBdfTQOK3UuvozkSd6PWLE8lFxJWGT5EjkoJRq9P3Y6WYYwa+yfkMpoAvWGvAINupY8BcIUEA1D
AQNnwP36X7mfksA7QiJ1dH0XmJxrE7svwZqix8HaNaC5ddRZKYSiICHpni2h0eg1GZP4rBFdkizW
S77KGIhh3/wuQz7pC3skPxe2TY66RMzBtc8VEzpkXJ8JF5Gpb24LUQ6JGxe/ZyJsAld13xzKmoPK
aj//9X5duWQBsLdvcxhgLcMbEvtKyt/4jDfXCvz7DbcDbmDG3PMw+bKhCLhV202J6LmPracdap/P
lexx46+vr/Hbn875lme0wvHLt5OcuwhejZV4gsG2z7thQxSZqD0CSkpsS4SIlVZGpqdKWCGadUsB
w25puCtEMvib0cS16tn8TqzBzDpVEg4kvVoInTaaVDGkHRHgVLXmIu+9mtTGsXFGZziCQVkvWM0e
97uKhB9Ba4QWXMxt1Olhrosw7iYB9hFmb7XRPdRflHLB7N8M7y7hfLO1quEAw9VFLcfq+f5hvKDW
kVLP3392SLcx0Yw+zLFlZc03I5JOyXWzlJ6Ez+sHp3rf+YFkzoXlCrNcqIToqPQEb35WlPNqwPgg
/8bmEEkFoShqOBQqiqWCUHUWeT4x4mFn/y+xuV3udJ7OWJ9WP9SE7NbVJDw27ZyCOi17f5OX7gAx
mxxVAkvSPP+iMQ20W/jZxTCXqUBo+7K8IhXKmMEn6rsmD4r/C+T8bXmkWMY9CQsCdhmd0QBpB0pX
8rld/Q72nNArbEuUNUibDxDAyh6wwvsryH0hp7QrY2zfDBF2PxU5iSBW1fETgPAwlK8ryE7xJ8Kk
DEazo2+MYeBMaPEihlVOcFWlJokxJZpBodPapfqNO2wkP0y6k0QUs8XtfKDPxEV3hclEyg6Imixl
FPfngQjbffnX9rWh6DOvOahN+PXS8/KcBh6kQ6dEeIDI87z4lWVPe4sv38vRYrcpgBxGlCChajQk
lEFy7BIhzEy49yx/eLD0blHuzoV2tD2t0iCQAq2doj0x6oSg7lQ694ZQcDZvcY/V6Nt27BwhAFc0
f7scbVVrG3rX976TeEaQnBJIQteiVR+URfIhZXnIpI6kyRruq8sYDLUT2e7j4I+HXe6LChzEPAQg
4ELbiwKNoxiIRztWBxqqMHgxmBg0Wj67n+rkbzNGYpTtuXVADr8k2wIWmhwkrX8bLDX64bmMF4wC
ostQfwyg+6VMQMruuvzI7J1U1+ApnDJaglNWEn20tBTRjX+TxXyuT1oOsTvGGO/g/Odcnh5Oz/xx
agMANCLPRWvzuwclmx0sidM8mKNeUa3uBPekqXA4eeQUY58ESNnyCM7MkaOkZ1l7V4XY0nMT+9//
RCXBAEY4X7rU6TdxdLLLwim61ZvYiHIFzkVBSnc0CSqwg5PqpAlDaK9o64+Dp2oZYVm7MGBNKiYF
E7e5YNeAUQG5/vgR8ipWZseu4Wg63Ss+rIwftTVJd/xg1emu61J1W/wY7y1QIYJiDn61CGoO50RH
DbKGTdPSJj6rUT7TVpsuyecgT9l32CB5d3+4l/CPWj388tAUMVvZB1E1QivfIf5Fwo51I4VL4DIQ
y1NAninlkNnp7er03fJMGps29a38g+U4JR4GSQftGcRurSta+yYhOJmNFVrdkXqZO1euSdJYrWvx
CrvM3eLPeAoAf5WWjQpDHzl3xHDNtuDSPidxNduFU7ard86jkx6GTsEqed3i+V6IypeGJWx09Grz
Qo0R0Pl+QQjrVSwQ01cRoH3ekw9ed2hVblT4RZAYj4FOhDc9bXiNYylDBSKAQgRM2dkrdkvYc643
599MV2WlEZHUAoXqGMqqd2XVTZYsAgPnq4OLdGCS8CXnvwVvtpLJ3qMmdCcFRrG09/YlEclreAiq
Bi63JDSEMAcIRetsaaXVb4I0Lg4AWqbfpHDytzBXIXxfuVizp29FaQ6TOnwfJRcMK7Ef536hV5AT
fLrkDuIrrsgsHVj3UccdjH6cASZHbqK/hHKuBu7v82oU27d+44AKSqMT5f/3F2HfIr1t0fkTqF8Z
4/Lsc/+zIiiWrCIw2X56I51XirGWO2y2Y08OVa2MriP5KC2i36lv6I7rVct9HlTk7yGlSNWhhP7F
0DAR/FcrQDUUrXfDuKyd8iMNIMPMNQGUvAi6TuK8hElOlOgluMhLvF/a6xuZCKQXWQWhDHNm3GUW
4bCTCSbMD6lyP1ZkAnWs2TDpc1AU5jzGi/mgS37HPj5bQj4jaPhFIrjOBz5yWqm0xGO6aVq5nWgO
w+sM7W69W+fyw+8uIDptT9WcVfr/c9Ar622pw5CdWZa2vB0FxSzddUFElvrJjcwGE0gXm3hyfDAV
QVYFtDtm0Njd0k92ecQ6QuOoj4RdZJ7Jf2Yw3nCL3bVTS0vXr/DgL9BQ9WL88XXVb2zmORjx30VL
zlcVU5cHtJ2/8yB9Q3/py4494DBdUaZ0e1ah9XETs9G7AkB9ErAtwfPyLX7m6tSipWDa98W+u9Hj
ZofhnoMCX6bz8UvpBhJSNfTKcizSJ1dapvZEDcxkM10FmCK78sEASzkWtpSshrZXt4iVYw+4GLf/
T2BJzqDP4vh/DjsQ4quFxlodvpOn5fY9jNyd+Hbu+g4t7UoMiVAwAixzsVVywtCYY5EvxZbzIMLL
DgEuLuUrADxsshMJSHe/ddjnBETqQKlXmNP2wlLQRuXwnpQ7fcrbDc7ocbnjCsRCFrkLUxRc9YjX
IZRzQUN/AkhWVzkK0l7sh/Bi4qWi7G2D4hAh572phQO+J9xJFtyiG99SvxsJnfNiWYhiPibHWHFj
RSRq1L57ilFkjSr+8PaVdWbGyCL9015dQLD33pyJndEe9HYkKJ/BCmxolUvnqF6iEGWSxPJacsMD
fcKoBvFpQdKp3JMb+zgmBfl6R6opD2iq2vGMS0e67XdKnOG/feIkcZKVhJTx4KWJqem+wBTj1RNE
HaLEf1QPu34qLxJe0SzuFidEDxniJ6eEEVU//K6Ux0hDgmxLFed5YXYADGsvDV0PYpZzuE3SdL0/
ozjUwlINN7W2yG87L+av5OCL4ngF+q+qdmeQoIsDqe4De+R+tC68hhRvT6ED6oEKO5ru6X9bbT/l
gl+07nU0/eb2FVPCoKtPwVLgoP52Ug0ASXCt9NNjvVhoDTiowq8nUTkqOK0jZVvIVFLgsqUCK17Z
ggF8D0ZnlK3wE70zETU7XvisMi1iz5ZGYUFKx7VNNbhwO4a2X9gh2wU7l1U+p0cBf88zd3McG/Qe
RKmKYFJ0mvymcuzrX9Ps6JnLbpp2aTQf9mdj+GF+L3iX+9wKD9h0fem2qzIjowlEedFliGCDRyW6
bVj+nsy995wL0W/5zs1Ske7u8Uq2SbhvrCAqMEGoJQJycmPVQX6T1oqtmo6SPHt4FrcH73wxeSho
16uvPYz1tQQvIBuifQftU9LsnK0GWi4aAV9DC//ZVlwC2GYLCiHEfsWsWYOx3svL3dycJa1qAYKu
cReF3v5AEqU09MNNcPy8OwOhMSXd9vI4quImd9sf8Vx7wSERF//6pRBm3VW5cPFQ78+XnPOOwVvR
1KCjlwLobFKfpJD+5Hu2BGpP+9A0CPkdH+ckhx1ABL4nuMIkQ84se2slUwFruklPtjPsjzYlXBJR
fqcqGEUSOFVigMHfgIBrvvVJ0DcQl2lnF6V15jCjExGIKduhXa2xLtlS4JajXlyV3WX2i0jMnpQF
QVnl4RANKNX7Ec/QYQYwlYcEJeAg7g9INFoztfgF+ehvgpbF+GE3AJs7oYFof5K2Qft0Jzl8oG3d
U1K5ypaPNzLgFbpV0OCjeXwhCDQSQAWm+o3vqobWKEGSeYCLuFBe16+wAN/bV6GQJ71cbxg0MGk7
bKj5fn9IeG57fB6+szVS+JTj/e9DijM6p6fTYx/6OVhkJMc5ruYfXq3Pnl8SWO4k5Z8FIzWQOaUN
glTgfFGXAXrIfFOevvHSCROYZuztRBOyvhERO81S12mgyYrULgwgIVBBNWcwD1uqoSKZnEQViPvW
iA2Z9CM33HPJEELFkrvCs3HuKwWMBJ+H9A5Qq05etIaObBDx5NJ1jm4aHuMLR1TbzlMyVg66bSND
Gis0mFyYytE979stWj6PJ18bC1lY8GBcyV9Q/VJz02LrouTHDsILD7S824Acg7cTMGpUzKLZI03S
pUM69s3UxHaJikBcd5WkQH8Z3aqRJ7eDmkJ7ES9aBy4dMxNvfVrMP6OCRJPNb31gJKwc1UZ2GeMr
0c+SWPBOcXQwshQPWhxo51i96ajXo7MsZFdv+9tDxKLKqdRRljQ/XZsAu3VQZ5gVP55K/cL/wxfI
RcVgukg3bm3RcJ8P3pEcXpYw3CFYAY0KLC0ZNPcyao06nXu+YcDg8DjDsRNziRJtxOBaYy2JB8rO
3jFW1hoEKz0VLAh0X4eAiJlkAuk9tvbOQZlCrRKAg5OmHiX5BtSh+juwfmvKUDAvxs8SVDpjZl9H
NNUChesAPHGhKU5BCVrHK1+uSEXOWPo1oDj81xgqWk6jeOTis8ipx1JYR9ytna4Zvx1iLK5lMPL/
XyyEA8iNVQK7WfqO/yZ55nEb2Vh7nbFAtco3JtAzegqNdDXrYjpkAiJXW/kqi50YQwshPaann9fX
OETME22sVJrUVCJjJep0MrVRQvRVRQY2VXiNE2Uvtfl9tmgIDVivpmbJBHmsjZRWlRYkiLs9fBLp
TDksZupT4H5pr8caP1d86rR+zeybQqnZjW//Gmn3xpNjmeqg7MTjal9holTzj6C7kioHrzDuVU86
l9z5Fknr1d79nDQoEpDNEzD+J3zj0ytzWK7neMK6toJDqDAhI72Ko06kQY8IWqNvC+INmTL1pvC1
wOmoJvO01bkjKVxbyNQUQhEZ0/AsITdfmcZLonR7XX2O73QLleVBE07kwBq2ETx2lk5D9R23JufO
WPDKVw7M1W/dmTRNlDPKO0souNNCUdUZE84H2XAp6ZGAue1lTIfzEC+fSNmYbSN7Fvu+DTVMnYnl
4iClJAjnwHk3h0KXj5zlBGcqxtjG6q5KmpgkbSpe11AATteZcf1KLywe2WX526gokuYug1FqIQo2
cHIknCa81DknyzcZcnjWY0tN8xHEhD8xeQsM3vMkpqhCa0mAmvrpIDsQ5MqqyRPJvKdKAMt+n7Mj
pTarLcxLalrzeXX6w+dmLBwLcBo2Q5ExwP+cCxFNppTyw8KY0XGw8F7sv+W3ZdEdsmZbeE+DvlCb
F/HKONcCXFucLWUVcyHvMNM+lBj2oYTgoJX/+YmVYlTHqJi5XlJ9yquVSpQ6XhmoVbVQl54EmlDZ
ohNWPA/6ha45vDvK/MSIlj7t7Ar7rFVxHbDSgvOYNoq/j1DboyYBEgKry0fb+v89EgN/D4HJERNT
aLIeEN5ZS9qMr2AfK8My0L/pOm5+flQA7BuhWf0Ep0YrdCCfwcXK7EGP/6ZbBjEISxwGHnuQTVnt
NouX22jZ/m9iTCYw8LzwUZd3yNhgMgUG8quX10OjwZh295GWpM7AvRgnqZQCZ2CwusLKydCT0E1G
NorpPwgHfleRnI42sHtGqFwFsIneOp9+AFHYhFocmtr4/SY7doyWMa/HyWgw6kbqqdEixwWmkAUz
QeJOzfVNlJ2QP/VDdVr1Dt9tjPzgyunHxQ71xv32Whnq+HjXlu7KPVoPWDpsnx9sRSj6SsByQ3ls
XP3QOcbHiuLiuIJx6RgKNqxU7ci8BO+Caiw/fNS/lxzJFTVhc2zkiOTmg2LgveUo/XxiWie40UCf
X4A6i36i/fQRePOLIH/ked1EIRC2OiagV/lkVMqn0QOq3WywgfrkHhaeUuI7LyqOHWzkWekD9Enx
EIQXS775FPSPFeRB9JTxwbb43QqcqMoGhLCJM8hePdRJtnZdyctw51lwMERwvdJxb42WcpqO+s/f
VcMtVCZaTICg8DmExI4wmtNLCC/VkBPbi6SInD+XEUH2AZEUMFACp7Hi2+p1fSA//PSXv1NGckG2
1SntuKw6FHQ61VJnRKPBgEgynbsPw5pVKFujYokRWrsKtFXBWrMJmuvZ/vKNp12bYqYglEXmwuUJ
bOYryNwDHIHjfO+qSeEwzE8F28EHqBme2iEti1cW69AgLOFqnT2y/Emejf/OlqYmzc5EQLquz/JF
xeNIcRPzDab0Ia9NX8lh83jR4YO12omLBQrnZE6ZHKmBxqJo1Rp2eURJMKVe/iCnAxvRKmzkCCHE
DABOgmhRJEREYkpuNbaR+pRH7OB5zVP/rpykppg3Bm6+GUE8VQI1/46/3ygCeWQXaGVfyaMCpdig
v2oN5sSfrNuXdi2sHsHpNSv4DR0JWZHhQ8vZg72Qo6LulcjxvsXb6TiNm6HNN/OPLnoP/CPy0Elz
S6PobAZSi2bn+Uxq5IRjAQD6NBkPaOEJjvfXs1DY4cchwOmFaRE7rHo0Wo8sHG+BY2sHAS7spOzH
8xMXpvUzuPJ//b33nzGkVA7jFa4C6mK58inV/D7tMCk6fu7SSpa9KNRNvWTgxRKPXpF/LxxKmfcg
fFRei31130H62VAmFTPvvBe4TPgJxW/5Pz/IImwPVWe8q7EeyxtETEddagDV6DapUw7JBMp6EqNd
amZsU8whbf5QU3B+PadWvbXEvN2z4JkJ8L869FyZOebyQXJh1yuWLMl5C5IQk24ievMeMaKiv85k
GNaCS0GNRk3yvjRTDXfrPg1RqVkqONCjowQZL9vTJemWdfBzECUEpi/7qtLJ2WOXBDKnYCPd3b+P
kKkXx7CtJAuDbN4gtKGgF/mBrOIz0D/AhuLr9qd0iMxoxDx0Dms+GH3sYddFagDZtGRs9YcdokyU
LOHBW2JwceT8oWYnlRcyb7C9oqOSaiH6mtuM5+Npyvn653qWtutRSB0so5OReO8d7o1DtWRJVt36
AgeRGj58n8xw4IxCqSR8paTgW7IRyRv/flJqzFxfly2OJkNOOoHaUKWoMJD8axyxrdRFwlL9TMt9
Gff9rbn8hfA1v3+ak17DRAkIZ1lnx4P8n7LQ24q1fabK42Jyr2cllSycrj+HKkLaUVXPB8tIYOrC
iHxJkNqkjCTE0SmAXw09TWgveKhCKOmpr9F3t8cd3JswWElkpVTCWCpAOJijr3/oBHFPElDAEtLo
Vghy0XEXtsVPafNkoswHxUkprmlse5Ygo5Ge+PWaqFkVATs/JLka8YjoD9rO/W5T/90A1gDIzoWg
9ayU8F41cL5tUIxdlppZDJwdppDpXOphF8AhAjpACScwoNhQloNSSiju+8Ujma1gCZzFibS4XujI
o+gkc+1bx014NxbUNYtE+nKSok8V0oFcc8U/HzdpT5zX5+JZmbv8EVPmgZkeYfTb40uwXK1JMWSb
32hqZa0DTciAnJiUTrRMbRwEp9Iw5KmFGIEr2WHqyEiPTFlPFi3QekvII7w/FEGiQRnsb603vqgC
5iMWTq5tMv6DWvuo1vJGIB8EffjQXYeV8jdw0AiyFZSw1TfPj2UtEY6bgJTZWMRbNZOpqdHiVjnj
o0hlL2Lo1AukEvOBf4hyBw6o0mZHNwrhw7uqLL59Ns+kiCkrGu6zmY14qyoZ6B4U/yR4pJXY9SqM
ScyxDXL+F0exxn6Ku9ZuhrAQmwV6rkFugtPda/IXyBsJv5f7bsp2omO4czhskkI2z+rte9uzrcWb
obpIYWHWhsLfDPauEnuPCBbiMSsa46+aNZQhV60rIf7tFV2zIevyymyZVIEvNrHZtRDAZXii+//E
3KdLyUieGLh/SksADQ8yRraXPMQbcBCYc1zaIFGLfSs6SvWLrG8uwv16NDLATcjdWet0hJvBrccJ
f2X7upqQ08wGa052U3mbdzldLJSgVzkfSrgDC5INNHJW8r12jimRWFcebdLgmf0/WKc+wRlmffrU
wNRoQ+A43pTCb+01vjT7bH+xEEhpz5w+/yO/XQgkPfxqUq+/+iDpszyG0DyeUXq0yzM/BbOT4xRP
z07iUIfC/JEo8sUydiwXacYONRUp7Zi8SL2amveuIdeEFK/0qEofwDKHQPbe2zKJMkFyx10eqxeu
N9U7FSWIdb3+1VU+5mKed/37YOZ01c3TGzbxUgfLBP/3RsSJbR5z9UikQITfa0TtvZ2+7paIStpx
/xDALjw/oOkAayECADxjV/uOHxKBoO9jBPqgcAC2VTy6YJklJiUK2pyAGu1aqMQ9eH7PJx+24ha4
+Il2oCPTEuXo5obp28adQuM6gKcbW0edo2hIxAbGV5utKyVniJibd9PMuFGI+gFjQLYK5YGJovjq
w4kggY622uAOW4UX8EBX2QQHN2fYZAYtCjH7/YTSH5JMfoA63Zi6263On8PA1qHLlYG5D2wKhMh8
N9/IdorM9mR/sQJVpiQMYU/kXFqn7JNyCjSoEkaGiE20Qij4ZCHoJFAjsPt1vkXN3HMvyXP7vEGr
3T2zOlZ99rHPxkC1Xj3LMaUFWSfwTxpt7mMb2XNLnB38lqPpf2x+0ck/B11N6wZZMZl1XWEXju71
80DVc7DDK/fyeWEFzhBDHDs+6fUEvnGENs7kVumFenUJ17hNk0yERzs7kP7sHQPuud4BI6QM8ayD
6lsoLqY++JdCh4bpmc6G4HH3WXY5ekkdibVI7Ia9foeAbMh42SzHIHcCXGC8I8cG+zla+nFiSPj0
MgYKN+Qmq59uxXDl9ClqTc94Exc2LKZ3Z6+x9YCBN7x6jq17hLY6eLQ4GQb8KRJx+pDAwzvX1gB7
bB0tJYuaWEuwZg+TANUuldVCLZH+6jmLQ59pYPX33mqms0kBMTki7F41pHto/SaeOPwzfC+fWkoU
cZkDr4+FcBPcQgrCgrfddIlj1cDwKKbygKSk5Xnvt2mXkbCXI+hebhP/9LbmEe4j9y0ocfrANwX5
Ai6mGzk0k9T7wzKQwv5tSGquJSyWM/xE91Ya+LGbLJ2nLLcyjoMq9c6/7qAVnXObwHLEoR7pAPry
scjYTzSjFbcD8JDJsbQ5rDmT7E+SrSTda2egFNsKXgZXFQGOqoln/YXDCifvB62pCoHFWSUbbroL
G49jzNLjB9Ix+xq2bimpfEfPdrSK0M5zp9y3HjwLN9cFG8VPrew20bHScP/qjBERvdAN0aOuAtv6
S+XJDwtAwpGIuzzWKFvKKxZ+yvnBu9RBiVbWF75DdEAVV+o2wAYHkHlU2wrd0/P0uhYiGpjPsBnx
XaDkjPyHwGB6JT7xJb0Ww0hhUYpJtckaxMUbiskEZ0sP+yekP+m51fCLMHnT8MlIvDEkaH7FAe7r
p7imIuPPUWNe1T72wg66OlPEoyjEZ90YTfpp6wPKGZ6+IamnAtcXnqTGtItg8JYBLZwxNma2kV4p
9KJ1gYLJvz6T0+II36c6GrpNkK+jAW7b7B7YwU55NeyXcMmjMHs2X0orVoe6KZQr4gPBUAMYR969
FbhW3pAqVVY3bxG+1e/rD58M7ldfTOtJeZ/id5lNF/JAe9Ul62nwIzFu+G8LUwpC2mLJkhPq82cY
BViC3RwYWifw9HLKhHV5MB6dTWgNzQtZTG3FQ4IDw9C00DUXWKUuMdKxw/YDmi+ldUQHM4TGl10X
/Wn/fKwg8NtV/kejx5x5rlOzQY/IFYoCo9zfaKaRRkWHo2hKGejkGdz8bhjS6D3MAtv91+HKYBtk
gVaNTSM3v0rgvBUcuyFz991DYMdTPLi6qB2X0u8bk88FSJHFZe/13s1Tcf//Ybl0CVHAfJ/SPAyG
q8y8YA6nUJm5yKbW5FheEBeAXubC9csyIJEjwZDAMZNGHpp3m+qwFKLQvr1J+nx7p8yxMdiJD0TV
wcZ/c8ict+Ey5rD7GfJ8CcOBOVpf8N0Z9NFjGO5Jb/hMxWgR9t+0J/M24I88X2k2A+UMw7Sl1YdZ
XH6cVrrJM7mB+nOfLr/HaUdZyoF6kLGU+ImWq2ZwDZoZZseLk2O//nuNpc5IHI5SYyyWcxxqVGp1
dOODQphQUuKNUdf5gRaqEkH74IEWOUC0S3Kbky8F3rmOZDRNLWREu8LjzFCN9voftkFMiy3FP0OO
1ocJDL0cQ+8I1wYMKC0xTX7GayfYJWlUW8Xa1Fx1liLNmCpRVw30+sWYDQnPxrLO10bNt2A2dSby
aaegaBhFDs9wOIc0TodZl1m7V8Ox9Lfp3zfSGO8CzY14TXgNdmBwfC8fEopydNujNL7y6IBZfueb
ZJPu+XUuGSZ0Pa+BJ/ZIHIUPdVDT9DA4zpiFnY+K6RGemDIr2Ccx9WzPUhZ4gxBNjYTy3Mfioki3
/Xr24omLxS09qIJs8kyeiWrLbxG3RNdL1eguzPFb+084QZ+sYEd3J3qUM+o0s8eJb23pUp14d3Uz
J5h51Y7bx8NCaNApqASov3VG3hlRMdjP1N7LljIP2CkP/DAAz4R4QDHOl3tS1Bke2mex/R8ydWB2
NZhVOl4vgv8iXf4fMjnj16eheapU3j6vp/PZ7Flje1F6sx1wLdPWMS10QmTijcmErs7DHZo9DmB6
P+VPU8xnQ4R/zJjzv7sYfOQeCgauLotEsPhx6+fpJub5u8YH7XiCWqxGPwMTPp2Czoxh/zhoEm64
uET2Q4SS6OsV3FxS21VZVGY6ChwKisvlAW7wUBWQQ/Um5kf9vCJtNfu1+VsBxWaK3nfcFzARKfEg
JcFosGRLVUBOd8hMsKiuaL07HMGQ4oUKWupEpjuvPzO4kNM1la1WpI9qTwRnSmm3cUkPQUrvN5lt
WwnoQPAx0RiRyIICl+Ungx6f1EMg0VXThWgciA2RQt5rzR3xgNZwlMHJ9ecnjMHV+2UuswhXXdZR
un7VhwaCJk3AYggWuWOe7/7fzuuV1ucT6d7pYb6SyGG2IBf4MDgMaa3x9zbIiVALsGuD57jsSTO5
4TYnI1HIEfV4Q4C+EnBGgR6+JM6VSbNBuo6cO0vDDZCws7ViKSPew3CWVII6NdsCLnUlOHSeAlGN
Z2i3cy10TLtd6DcztZvWUXboPwO0kvpMMu4wsHWxExWCJm6ry/cSMfW0/YOSf8uDpl20iwx24FyN
BJg19xYDgvCbKOKA5o/ti4g8xHlCohrWm4nF/K7CGjKBtFgBmVF4duvULobdofFkHVSi1C1L8ClC
+/Q24VARotc9PY/tJrVLqamwRUFHFDDTa2ti7U3GVtrs4FHYBlpmNjOfOygLxKKjFdWnlC/Jj1nR
b+WccR5ETatHgjnJke6UnpCU7oJADdDLZcDFFyEqzHt9eXO0LlhPyLg6U/Fd9imty99p+2z8dMRu
5AzqWJIaCbdokT1Qo4z7jmBaiDBlrJ5pEaCWXIOM0vBWb3opt+P0sX4L/oR/Hyp9b09lDZxQ22+I
hqQAQZmtT8vGKmNMhmyR+W2HndwvXcQY4wEoRqWC2voR67GSPveofxtWfJhRykjlEgl6uF/ecCMl
UK6YlHDXSyFeaglyPsOdoDFcvEflCtfsPZ9Tv94RKqTKQg9mICUFKWM75Qq3ulZ6C60Jz4XSzqkh
mwl6JtXzOR/vW3Tbyx8LLu760sGSgGchpKJaY/6EUOKPXRjlFzWuUkC4UIidsr+tzfeOvSaBu+Bf
0Xhi/fGPNyzZQWwERmlulsjx0w14BFeklwu0GfJtH3dFxIhOSbRGrIZbzkjB4pAvYxsZuyljf3JG
L9zZBvGusy3d+i/R81H03EGF7nj3fKKXItqZ8C9LVam4i4NYm41+2re+FJTsakLOhl6pg2Pajnyp
Q9oe7BqVQvu5ufOz01jDnvEIlrSnAhB2qbRsBIE0A4W5uXbRuG5/uCe4eQqxXDpDqmgs5V5zb08C
76EPOK7LFSDl/sE/Y3/Q2N+abJJpngTpimYq2F5odRoObbc/gsDU8XN7xgcaqbPnhXRtsPWImZMO
YbAcFUmTxLZHE95oBJ/NTw4jcSdFqC5DIoeLEZqw3OVFL7IM0vCrb8bvQU1JtMKHfz4CNyXeefLq
gYiyKt6CTeM6Z3CpAaqjCioxjUxlJ39SydEDxoMGXqnepcwvat6D7+DmXxDsC60Rcb9196OTg8Jc
cJCaK7YBzXGcJvIgcX1I3mHcmLkB0NjxiSi5+49hO/z3T/gN706WHo4ZjKPUxOKWYFznUSy0Qpc0
HP41bhmEC2B2poDyVCQCw9sSAQ8YemV/nSDxqWmLuFPi3y4YTi4cX33GdvwQZ9hIFhcCjPrQ/36n
MG9jsRIBSQVbcCnonXko5xEoisSQ0atbSP7SAA4O8jNK1LVRCP/NmstW1FFhPZb4E6hnlr37aq4Y
c4s7IyHIau3HVIIhTe+I73uPO3K9PkudkwKE1GdgHm54OW0P0zfW+xUTHCkq62of8Rt2jGCyFodV
jccwNK8+YYXw/hlnd0Ux31ROJPd8HJbtw5W7dCqLwyQw/CSMwupIxerIhBhXVQitAfePj64yG5/w
5xJ/xkfjhPTyHyVjKtGiYmRIEpssNoWjGiD+OVptslUnINb/82n9GWCM2E82yEDZRCOXvTmLLbX8
Qi3S1ejumc5+BywEhxa4utTrpYpQfbbnHN/TshHn2UKLvDu/7rV8BjHjibdDjifjL8b2gbqg3W0N
wZ0TU3FNYAw/qq0ihULGnVPOlmnWJB6nJMmsOTOBQeqWu9ka3sDeKrfmDd+QzLmO3niZbB/v/2xt
Mu9PKs52ylBt+f98O97cWtmNsnTuVbayXEuUKH+2GKUMrKLcYQe6ovN0A7fT6/ZdfZ73+tTW5TX5
LEomzBk/I3em8pvkoEUzTL+rDJK/a1aUDUDTYnyg0ChRzD1+RAF4WSwxcfevPUn9omq4gUT25MtZ
pvdXBFrSWHTEMnVmjCnSqwZ9xLFaYxzBp0UqtdyLvbrdlHdp4j3j9QSOPQ01zcHXa8ZJ03tlOGEd
bizcXwQNo2F79ZTrnKijrO+NUn928CE5JNodoXi+BIvYnATD/w/DvCBmqTSovRAXbIO/jkrNyUfa
bgWU/FWp05AIld7KTHrsAduC8fBYHkmpCy8TSsj60i+IvUtzss0JjllLhOU2I/xkLLQvxHDl2l8F
WDSiRJ1V6QdJ0ZJCYhPjgdIFGAlN4LBtR2gDIPlB57QgTXS8TQt4LUrqVvYI7hBuflKtvXeDtHHo
4vBek8R810FUVa0obpgOuMZ9hnwWVUtIfdALRaOAfOHcTnvN3yU4OHdG7D7q2U3ooT0kaet05zNH
s34S0XkWlj0tWdmvMnFYDT0ynVHmieoN5vIid9+rnJCDPJWwP8g8ulumpTMHbF6T17EP6qKq29TT
Do5EM8Tc9M1RaKnqJ46z2DTECvpUP+UbAwqU2KY5Eg8pt/YexJeT7tl2KHmScrU+4cHSoOUh/oDb
pfX2UvGXd7fCfAJRMO1DXYkMsq/b8cHO7v49msj9mqv3rtObLB+1yxPqds+Q+Wndr/ywTH/HvO+4
boXCFBklTxoLap9x76VKXzgnsLUAQe/oO6ddErf1eoBpx9xdqn5zg5NRmDqDEsh65/9iRwrLvJM1
5lu2I/sCZZipbRNTHezb8KUx+ljXUYibxMFywIqAHqK861rxaU0KzyhIQXg4xqekp1yXOsCBYVN5
WtQnUZrct0QIWUGPrpc9G1m9qVN9skaevtcsEdSH4KUtjKV81rYh3pxrdD0qMr+oCyaEJN7Vl1D3
MjJULgnqC4vO9GeucwEP/hDvxjqEUM5dCZvmeYamNYvznH0sxjTOVJ9Yi7d1QdCXaGdVHTy4KkJm
2Ym821RvXI1cNljCAIHmh2r0GYC9o73/S7JMD4chR68uRTaNqrqwhlxOIF4CA4zOtdFTejzJ9dZE
auE8Uu0J6lWGz8q3kJQe+L3mN1gRsz0XsPYhlmQrQpSspCRjgouBemxQmzXx+GBg4SHFC5BPOQwI
RuUretq0KH1R1dAD498HIT9K3tmtneR8LUWxc6paH8WgCUW3o6Mrpp8lZAcqi+ngxN60kS1SyzrL
xOl7nYs3rE67ZJbCv6E23/NkFLa9MR7HTuNFqCTuZyBbTSyrVPpfoWXtiVXCmNFYR95GscVpU01m
199RQlW4RNCNX2iCezz/D3xy9joEZBD2w6YNRyck8JF7E+inQZlMOejdJjAj2/lk8P3H16AzeyqN
zC1QfxQcl04+7UBBHhH5EBRGlPMHBvmJS00BQvWfQeQjSmwKy62hnH9C7AmaVlP5ZQW/jnjT4P8/
8pZLtXdsUQWjaHWQ8ksjDIhhsqcm2xER1BpkFB5B6hV5e9vK3F3MhzFezYEkia17KXs0lggZ08Uz
8j2sPzDQgbFkxVl5Nzo6l1O1qK9chPyqwssBxfvguhP19pAthJ+buhJR1MTDP5lDlzzxThpCmz6k
tbwcBPgMZ5l8IqJiuXL/1ESKc8zaX1gPX1ISuI23VU4+Hmxo0iYeqyUgH303H2UhT4FHqzA1VUvS
oDE7ZCy4o0PSe05i3U5xGOrDhDNiaF14p0MzD07IQUIEiyJrC61+iASaS/gAbOocE0b3MY7Zh1a1
V6VNZNhsOMPy2qP0F+ISMBgrnGE43nvse84dHKj4KGPYUeGvFkwH5SOqduCOmkLQCm8PGklc3N5i
wNhmcK00TZmfA5ZP2ak1wWSqDbx1/oqZMqd2E1eX7rG0GHjs+vegnr/vR5D/xFeYoQaEslgDQG7a
j1mA1R949ucPixJt6SVqXgueAhfIgToHwOcLqmi8oDz3VKU0uVOorVGdWH/z9Atqiii4aZK3DzQ6
0SYJni4Koh9t90NtKFoI0zzBsd1gxdCq6oR7tkeQFQrahd+jWgexa00UxMpANUjmc1t7487zw+AO
HL24JGPb9stiD3CTlx2pqROshMylKcRiWJgt10vjaeH181PPJyAAAmqT5fe1D715YiGZxdT6ou4y
R3ekiTDQsQo+vFznQfq2KTg/Z5i5M4wq9N2wHXK7crYTPtD6vKo+5KUE9MaRbz/9qBBbqpthvWXN
qQYCNG3/UXsg2sOR4VvFOVHeFizghOJE8rbmronWAr4rh0DrNBCMELFPJ0LXn8fkfDTBY1P4+mYN
iW2+12o+BWhKAlF7OcSVJfHZ0xJZZfgq64NUeXf4FiG6AblQlJz749JWqZGgvRO0xL+c/TEr71f6
aAzk8eDgqbOz8nKnOdTrkpXQnhSIVhLJABXrFSbSdAkFQ2E6TC0Gq3B24oP8ec2MUHhMfvBONH3x
FJcvCuK0qJQcemXVY7toCWzBwXbaK9eLOPAWT41yhq/fkX5YGZJ0Tptq6SQnbFcYyxE03wCiJWe7
IgCG62oDxfu5pRvH2GBcZcZtmqp0sgx0NAnx4LRfILthFKzFbbyB1rfd3Ni58gbMK4oXt7dpFfGp
dtUhUUDRvVLTSbzDTBPbdpUVU1e9NSv70a0d7BUgzXB5Ac4mk7OZZbf4hkbaZqWmAOE1zk9KNc9h
mJlPr5xIs1zh2JHX4REGoReAN4cgA6UzYWqMcmfSi9m7jTE2s8Cw+TA8YSw9VJPApLA+Z2vD1Hwa
ht1zrj07Vu8lso+2QiSlL0Yz2nivpkfbylD9as4CnPMQvLSBcUfFE80emZjTLKtn4X1PF3c/LSLY
S949UiA+3WZ+9Pd7Xg11TwS7+X+C4zYgMjeu2MqS3oN6ZqyPYOBNAoa5TnQIvT8wIw9Z1qcJ79Bv
nxxWhKIu5nAej5eGsZdRTqcVNef5a1EfdNFeoR9YUO4BLtHlFICqVCg2EQgQwM3sTFV7lR/TrAWL
sT7H6d5GzLH8308Pxv6MsxjBdC/+rEG0rMfQ4GwT7BWJkY9Tve6FaNwcpcWOo9KcU2QmFxDQXx+p
ba+0nGP2q0qhQYMcGpCxA7pym3Nq5WqAKyaPljUkom+WxMJvMIInET1sIzAWZoOkLeWIIm4cBv5o
YehwDFRpx4eTKpWYmLYkxSD0enhqPO2W2Ns19dMzm7jkMMjL0RR0zFq/CxuwwI3KKROZPmZcLE74
lC8gi2BFk2CVkKcse7njbeSTbwltKkgNSzwCzlh+XglT5kwBDJG75SEVEKbdnMI5cxe9NiaM1byd
vQC0rb+MDCvIG09v00BN9pFUTiEfX3JXU6dUZ6C9cxv752l/frmj+Y1tiGKGCwhjuBkZT9kxOX4m
FrCDRHsK6goyW8upT2jhP4utgP2D6BqdZRXbLZH1E1BkffT8nrC9hdM02/y+ivXrExSLdMi6HEzC
bhmg1W3d2WY2LcM8wI1zuiki2WpsHVxl6v2WTcZ70QCDImMCgknstklMonmhjjRDqK/uBGRuNaa8
hYmYKm0z4rff9dSTxv+jOO3tBFA0IgOzQXheZSFRtbUAWaCDtK9FYtErQe2Dr/ke+ykmpHj+G2bf
SM4/NEvWzRKIWMCxtemdcQRe76/fhhzH4qvoTAZIqyOOq9+Xr0DEi4YoAmXgoh0caMt4XOF/Z1av
cqHoL7kXhqwfqeqdcd5RGKdZpfNQQ5HaqW5MqqNBUtZRqOEQWXIzoe7Vg49G/ceywNM/mTSyC9gQ
iJvcfpTuspXhRjBVMplJQZ3NR/2yO41cP+nSQc6dfOFfo4iamTd+/99SUXcOGeO5UOpFPEVEXe7r
tKbzGjMhNiSERLIxutu4i+V3BN93dpjjFw3+G1nUzoUI7o3jBflyP5LIwGcQRLJkRj/W7KJTyo6B
u/xbusUzrbc+39qgBKdHhIDAZM2/uzs8gdmZxrPxp3w07a9A5pYCDE+5LO1T3tscPZMRTU0JqjsN
VEfJjiYokgZGzAJNnLzXnnu82Ldj7mkQjo8biMZkDkb7dmbdGWYHbzDVHywvdfR3YOsi4yiBMUQ4
knaSvFAnzgcYUkC4+w8Rgy0RKaHIpj0igpoylWQmWRvdxbTgy06py10S+m9yvGo2YUR7mwXWMd2B
tilp0jJ63CfmGLztDDjYL6TJ95sM7q3nU+1/fAtl2EtpY2wio7VjX3aDT/nspwrG2Pf/PAzQKxWn
KEg4W8JMRDHBZETI0OXdy+lq+qcyHfXCtzHoEbxy+4Bl2VvSLDMQRnA6i+jDsN+8T29Tsd827blh
sVckokgDVaiqrpzQoAFEcf1AHIHPRuSgh3hReKvm8dcKjNTtFYoVDtrcqkI7fYMEVCgkkiRY9yoX
r1z6k3pTq/kOwMy6AZXfCw7+Icq8nhH4AMy6ywiulLyQVxoqo9ej1yfLXsUiH3ouQVqY7iBKVd/v
JmabAB7n465Xj7+3lXbNSTNja9m131izAcB8vLHIwulQIZo2dR/PY3fZAQWPDoOFFRe1w+SQqR8C
KsypdqOuvfiyu7FktpBDQmt+n/atBW634Grzg7a9mOCu46/hQg3BA56lrWJe4VOvqBp4BE/cUwBG
6+1Mx46iAIdtDWd9YMrTHM5xWCDmlDq4mf3bR6ZFCVpjJJodkxV87gXPl3VVXrKOJd2dTk4dDU+r
XgwzM6azwtMjLRlKgBLGWI5y28WQqkqpWawaFVn4IPVaNUmSlC3av/3lFIBXgOnSLs2CTw2PmF1k
lRRpmSsGswMWCd/eEbZ5D11rw5/CIE8/8w0wjDxZfga1qiBpgYZKUKskicjhWe5pmIn/KY3gTred
9q8PuO17hvg4BrFhyrRd3Lu9GFI/QvmuffcjU0LVjdFF/PQ0ZnSn+qKM5OE1sb2DxNfYxTBt5LPa
Wbz3Kb7zBjGbmJrqm6u5vxOWf7OSIzN2G1JOPI8qazLRnsRLsarPUcdjgsXQKbyJmwGKT3TH/KsQ
OcRqHbkpRnptQN/M/V6GUx6RlRCrqR7UV7NeN+jxNVET4an90xbrHQgRa0K7huDNdoKb+zOnIEAW
7J6c20ZjgEXgJusSm5UmxzIBfEwmgLKWSfpeMYmP0coiw6yIWmOl8+l8HOZGtY/UyL4p7q8ae8X6
gmTVGXsdITGKmF/Eapc73wUVnmUUR1UX5yU6mF8kznADkfpm8VzU4dQ1+k3OzbDbIkR+PDZLWuZj
dmcpNUfy07PQcpXo637bc/K9jmMyptXX+9yWRY4PSFSgfKJItf0jeaUWxtz0Cff6wqUICkVmwbnw
fPPxn6jtYfI0v6Z3+df9NyDoq3il5+hQL37qCzW2Gk3iSSHBQeyv1iO3Q/zaAghWtouPbdvZe94y
3m6Ak8bW6NSuIuaZDi7d+dqaBXkPoBGHdBHFYAjGj+k1rNhBLn3C1DzRur3nnapVkxBO2FjSe0L1
ikXTtIbxolujBSk+Yb2Gbw6qqarN82jtFcFCTic1kSoyVICOcTdeiwSfalnOLqTssms1OVBDp4Ae
rr1QyhXiVgn4R6wtO57ai0T72rz2XhyRdLdWHAP21mxj63/NWB0mA+5wsK+raG4fTzUXCnQsrb5O
0EyL5blDnckRgYzv7gOxNtztOeow4W/qYev1WTme6Pl4IyAgcEFMYAXF2BANRJMRQ0PtP56F+CDj
4POrZoc2PrGWraqKYcJIUuGmuowCTBd1DXev/epBrqeLqOdlLDJRUvrPGO/lc16h4RcTuMwHaR9k
FJ1cEcS7hsRNvLIGNFgOOot11CZQeu18P9c6OTHEnWoVZ56DskD6Cr4Jiplc3Yat5XVk6Lw202Z2
JnGLGfiUgVCg63wF2CU7+Kt8GCEse/S9rEvlp4jaDDCQW02HZjiIEExg2x0J4G9TqGTR2zGC1Uw7
FDH7biCjJXNA9YwdRW6+dNBPpXiAJvsuA+FpGSOALxOUwMor8Ny84Gg5tIojhfMXWk3JCpQqiOtr
oqpxUYBO1IfjibjDMy4WpOHRP8de17fkQMfP9/yII8bnOyGPZUgHKaLKuHCj6vhwtJVvtzzZYe/Y
5u4pUEPZn1cXBM0uFeZtmWNuCQheLWcV9FbUL4ptTGZdAy7WTseTlCIHNfzbHCxQe8B3HbkTSJFo
fQZmbn6L9EF5uwgqej7JQ2zRoi4l43NmawGWf3gDEGD1rfHI5XsR4MA/mHk64t+68QS8C0LSYqFe
r5L/x5Hs60IXOiUt591kJm5lXWS44Gr7PdF2pCco7c5975LNuWoRl8i01kR9UDipHkvZjbqiy5YN
KX44AV/hCOay12e46OW+n0eNXAwvZBbm2UzI3pgDyxRqW3mz7r/jXM4luRBntrVBoqlBdEDMjapb
BTzOf9IQ95iG3A1zszBE0rBSdlP14gpKWbXxbev4f+kGHD00VeTk8GX7fKoRqBNF9jWHfcUYjCYc
A19dsMV+CuEO5edCMz5pU/8d2XmKL+IiWEXjngjUdSK/xPYGpCD6m52vOnjHhRd2f9aYIF2Pq0EB
+odhaF1Ev/z3Cb75P6Rc1Qd3PYJgDDTwyV1PbCeEY71o5pCJUDI6dBr0P0q2txi28wxrH3Nr2C1n
9hUusc6zb9XH9R8ZvbIloiMpoJVhyvA0UUBNnP/niRAlPfP0CpEAXqKAFti2Zz7Ya1qCvHKdUygR
Hcl3jFgAVq+kwBxGUWfEpRQJFh5vgXHGnSDkAYrKBGO6Ba1tZQe/IktjW341WVI6Kg3qvvUSp8a9
70hgds7T7vGEfucJNx3Pq7U7w6MuAEUC3shAgCprfOoDtTbeF4nnf6AsjH4cYsCXvHdgQIO4gDeR
g+YUIFNLSXL8g623oQwAeAEy3EhjGicWba04Ru0Wnem1xmWkVRVXo1C6zSJ/AeB9pCM0Bf5ZK/Va
NdAn+6qxD8STkvB8P6jpiICg2UivpH7JP/WhZEuKtSOnzH7wA8QN4NYxRBeisVpZVIbGmwhQsGen
p07Qj86/OduMOOoDohLgOELWsGm+YbxhInZY7rDDvPea/AW4ID925sl95TaYR++Y9i2aDjCXIESc
kIJGfbdcqRYwZdbegqLqYN0HvDS2H1Sl5dSIBAYy/y2vdN3qEYQajihZPlud9Iuezoc5KNemYI8g
f+Cc9/de7trYaXExmm72vvkEYeqIyd/io46E9Alb1IzTFcYLeix4jd2eLF6Q6wLguOXszuyxv5v6
X0dQkw+ErWovEeBEXjuz0YCKGiPqVY9+xwPGFuOFImLQhFnwk5tEjmT2c1QpDgFLGoa5LNFoBEDX
YYReTFcgd6wgshalNff6thJlhRuf3QWTEG5ZN+f5gB75n7V7AeuCXb5XqsYgzJ4ErlN9l6Lcol64
PyW7AHXyFbwiMf7QVl2FOVsprnimy/uRh1ea68CkVlC5jJKPPA5RAwGEeb/dECgv3NpwuSKamo2e
lL25Byp8xv7Od4jnkZgCXYMAHGvgpLSjvAcum+G+bLKFwdAo/V4GmuKl6tN1okJ40v9arqy+4qZ2
nFBcKhNnkZLK5dbqzfmrfzhJVVMXaG5P032LszjBHusUtaZXQXNoqMlsa7b6y59pXSKZ9evfsA4Y
KAaY1PPKj1M0ZiDekTVCbZfPUf3oFfKe8JBRLfK+yy+iPIVKlpYtGN19sVUks+l8lC9tqM5uXjYd
gc+cE5wQ02K+nQf81sCXhj1V63KqiXwlq3dIETA2DaK6rr5q2XjG5looWFkv7T9V9UUxMt2cT1uT
oBb3/KU/Dh6q/TpI9xWgoQBGpcoWwvIdM2dBc95GwQMcvjkcC8hR4CidvQTdot4LfhwyEOVXC0LM
4LwfDyX/WH/y60UlugcU7Zohtjkywz00/v79W+FCg3brMKgDcXtkN//OyUbCtLri5x8iripEeSft
0Mb7/q5gYuBVL5EOW02TWJPeJVk6xHrlY3Ut8hwFdMjATCPPorhxwpHpWkYtNhBrpoUh5mDB62mJ
EXzDZYKKe5c4YlKyPptnA+sOViU4LO5YYisZELKoTM8ipC/aGE4XoFSWhvynWD+FwZBwp7cunmH9
v7f2zZb3qu1n4JurIXLYjhwEy11WoPppIr7M5/R9QtlDIW5tcRo6PRSgTHBG1pi9JOTgq1Anrmk4
KISbb1L5f7oRbkCsjEtaogYXt/AuFc7Ii0D2G/TXOQkcqs5SIxEdZOC5aeae6dv7zejpRWg3tp61
gQK2luaWz2FZgaZWGcu481WC0zF/75XH9yhsdvwEsbnGfYJntKuZPFt77xNnDb5FKDxFpqZqQ/5s
epUuoUY3ohOdNjSLN0nnuI+XQCxA5rbe53djIdOfr3BvSiJgktJnz4p8+UVDksBvC7SFGitAU6TQ
sZSpcpseiYGMJnTxF93/0Rxb6TQUs93D7ZdNDjGEKUMYYCnT40JQ0K3q3RAxSRntxTA71dXFt+yb
sMuvPXNb7Upk0BEM0mtXbnY9cb3yFd78Rsmj1nTP4ggpPbLlfaGEKhMSZzC9knTJ7WgDE1o4qoou
qGqr4TAZ2lltslCNY0OxKzK7VimfcyZk0VrxfVyCVmKVsfuuqTsdTALj1802b+PNd+q3VjJ4hi4F
t3d17sS5uA9gXzEQlOyXUMjpzKgoVGrkGGV4d3tKrqz2U70ECs0GE15V0FAGOkpR1JA/RkLaZUTr
6ls+GTwqD8dlRwuFnfOxZk8iU1b+K3rAqLNJTMbQgzSlxDhQz3Rtlo1oNzzyZOBJduvX6FkUk8ke
K42XbVMcIiucY4o0TChbz220mOml6zPYmbaTjw4cQKpSQP+aIB0uQSAn6HDLVTAT0hP2gdT3uX7K
TqvISfDpMeQdefnYB7Oh6qx+l479cMfjxl6HMWgNa4OGb0zaVxJda2ojdA/KC9IUZm9f0Fv/s38O
WTwZJsc7YoxnobNMH80AooouVQRUjRxjiG4alikiGPIa7/JlI0cpdNv9vlICZHVFEydE3agQXgJj
u6bSl26tJB2RkoT6sc+kNtG+aq3HGgYecNnGoiinaFo7+PX2cISCsOnNPnjmMquES7Ob/Bwpuz3V
ziXVZh8E3l/Ugmwg2AhT2gpr1ldVA8FaRUMsadNVvsUAcOxsMSGA0vPPByt8oascjgoFGpR6YDnd
1sHLrN7sh7vvm75d4DiA/xZSWy+rc5mTrJh4M23E0PiPpMpkKQVP6y1icCM/LBDiOcxsDciOsHHI
JrBp8+imm4YqBr/IVXV39vxSOKVVwDatwmCoZR1oVCz0lpHKKp6EciOaUd/FU1dHjDA2cqJpTRDb
FhVJxh0IRWHWx//lrXTmoXJE+3vv5TVWn83uD3RLb5m+wB3NxEodwCqzik6gHz+n1XryQFnFZ//D
SAh7xOTgxB9lt4wgSfGxAZfdp86mCfSmg23rVtsXkhlnvXjAjg6nQQB3guIWsmvVxQityCWA61hX
Fz4HzmH5J8Hn9cRFGT3VVCrmJmBZSYzwuUMsQbdEaYfT00zQYJgceXQILMbCg90W8ZtfT1Yi2Ode
tVwvbTXccHFUpdkCZPor66lfIFQJ8cP3fZCrryZi5nFPI2bTz45VvR65uXsorYmXGZED7bo8+Pkf
1M050fUqmEOjbMbgFw/QVk07E+LvOZ8e3QxhBRkK7XGutfE32XPt3HNoblZnbksxnW3D6bGnLFTb
0uplsU2oSgtJD0xw6v5QHRGB79EgTMODqho1kM7BnkGN6dG27bseyKrIKChuNUNEZX82kNNTjzsm
QpjbkoEF0bPVxsbggSHfvZGpx7Of6vItNye9WpVa8IYOTqJ/5Ygqh12qGJojg8nhFZKcaxI4f4XT
ZEH80JYUSUXe7d9m3xWH+BZ1sJKBYgweF21rIDRMOhuYVdUzTc8nQVTaGP7jksPgIRU80hn3CXkd
ACvDW2PsWOs9c5XUDCUmgbpqD3U3IoLUkhCiENMAkW64W+7w82WNgYQrve5xNcsbkRyXZsiP6Ugs
K2UMa8ZISjTQIuzgxMXUmkqdShh1JDvxAdUET35zxkja6paYW2zf9ZvSLK65GtTKNdVitqTHYdw+
QIy1vt2ZJRM07tx5X6tRlLFTxzkDsX39ce++WXN9eyIKHTnIc5hQUY/TZeqtAcwoeMlFnSem3tXM
Bm1W8A2ojget/IK/Z6Gl8lWjU74Yk3V+BpmvJtH5mH581nLeX9JINeTdbFHQuiRh+jC52fHmTQ8Q
IwVLX+hClEp9DrfLzdUDC9WWjDaEqOXkUWnGELuLMDdhqiPmtjLpEVvFd+Ux+mxBtfw8yAXAEKdO
resJiYogcAo5ANwunVes4EbayXiyjl67AcUvH84Elwh5WDNiIln3zdfdmpTx5IF7Yus+rtokMwCF
iQsBRg31hRx+YB5w0O9oRCACiY5UxBQi+Z1wY0lRNJgegjX2ban+EczejcvDdnFes8vGDd7iEZF7
hy6Q7eUFIEPG+D6AunK2LRU4kX04QXrIFwNhaWo1XduR+sI0gKL5zxZupbfQaJunaxiU93sdBchh
WxTsGSHOHitIdHNN88ZxLu6VnyEb5CEmO4jvVZX0TLBZ46W3fKAdvW8lrnPie86Id3c5imVOYyvO
GS3yAwFf1pLVEvFH1NEQPfiTqoIeLJaTBG5hEiewdMdhQ/Pz9tSsVpI/v7hchIdaDC7UMOPmg5WT
ZXeOdi2Jq8L9QzmK+dR/stDtrgfowzZ9WoI3WAIxLsP1xAvmNktvjuWxGcAl31VXC95xZ/PfuIrj
UV2TcLp8O/xeDHxiB2dt1C0ogD710FBrREolj47X+kvmCZAhXYkeOBmQT0QKvX+JC+ffHUhTL4P7
QZTWYxkwXZZ+yfSEJPnKgWTessbo5Eu6naHLndEVXgOkr9+r3a6DaLT1Pq14lp7YDHXj32AP86fX
k4jSnZJ5UqZDg7y+G2PLtIS2giP7Lip31Omrf0UmANDxWSmtq3aPZwNXtzZIV/F3WICfXRzBzbPC
bHqBYZ93oBDvmy2jjT1LoQjZ0M4miwDlhwx7w1vHJsoeUsSsryfkbYtHNzJzo20UjQEj+ufvYY00
7EqUW1rbbM283G7WJyPm9+sdNP0jyhalKUugDW0gSQ4XIo8XZDkBd2uQEkHVvUV4ze7J6ZICa6w0
QaahO3ew5wytLuzKbc8V49p5OObf9Hc6BDk3gkNRHjFfwjOO46swDnvWD5IQ7kccqOgBmnWNeDVH
/NFxOYWSKjMKXo750g2+VpbmvKFMzlITR9HXhnhkr+fS1IqXrrLEQZkRp+UUQio/OFuyCaPymFhk
+g/8VbNi0ltds9IIj72wjA+Igc8zpjjQDyl7wAeYn06J0cUSA5yzzsSeTIjhuY9S1qWbNTelVXNj
hbs4YGEA+AuzSuamriH8G/3uy2hDm4bPtLcprJkUUiuZIqcakAJZSIMD8wXFPpKmyvr4UEvOibq5
jIOqLPHDw3ZnHiY83k7nsg7Ci2Kb1pBl7FZ22uB9uJkK6bIg4kqSFaO4Woq9mKr3GA5nXquN9Re3
OFlSGks4iLac3hdf9LzaNLw6VYdsNtFyBT6hi9gLUpfHI61U1kmb/Zoin0CPRvAVl5TUpWgrzIqo
fJ7w0/31ku5m22OJFo/JUQQCM5zuLbcnDr2JuUxUvfP2vf7aJz/GcF8LBP8qtqpMzz6UAHOqg2Rr
KxtpLwuecv0TqZ3Wc8dl3uw/ZLCWal9vJrp9fwWWrg7lw5OGQzlCT8VHCbajCF4nHdFrDzj2fcFu
wza/xDDa2OLViIBEEKxNrNy+kIGrAkKXyzqq8yI6wqLPYiMh0ZGA0MYuhtMwRoWIomsppbd5Okzb
lpyI/GmyG7KCm2/x4yH0RS4KKcBg9AL1OCYvAWCW+93ZowNCECbwjrTJMxVgXqOA2qOIbuYpCBFJ
slzX6V6olEp5eHABJtV5VHrHh0p89co4L1Y8gN2BL6a6em7iIOHo2NxXHfGjrrVzP+1E7SpTqcsU
/l5kIa8kr/Eui7C2YS78q2UQ3dB9VTN19IScEkXsk+JQqvSj1JGSfOv0tKdR3Vw12VD5yjd0MTsh
qJMnRn+6t6bgQJ8rKHNu6RCanaKysIiMO3o4TFaIApaWhEzL763ad+a8BZHim+aAbkTCtjUlgYGA
zKrHo00XXiorxXTStJExBm4/J8gJZWfSBSw5dCzlF0jyB2GD6SQ0kx1PEsJJdlKsDbuNxE5PQngU
J2+I9QphcUq5pQVeTlmjxe/5KmIWC7/pu4mRw9zQidpalPsFlbQbUtF1TlqZx6tl8h0iP88Hjd7D
rnK97GnQpLgZTaNCLUv8yZqJgONUgo1EgQPm5ZIuaSRWTAfbXwHR2LbUgSDO1IQwNbUji7Iyapqh
SO6hIY+jP0S6QmipElOtmEOGMB3Rv1zTDjxv0PwTgLTCsdOtyEcZvC8ea1K4HvA1gjc+oajq95wt
x/wl7baNtLShAP6mqSK8fdXcIu4cZZvPydophGjKCbOmOKqw78XF9wBsFXhTpVGZvjEfbvN7HtKg
vXIIBJ6Ji+9EqSFh7mp2BoJmg3YZnVEACD9Il2Tu1j6JA63T0lquFHft+FkXIUStmfRDUZ3rytlz
m2H35iSXLYrcxuRXYPD+yrFkFOICxCYnk3I1aTtQtz9mRO7A/LBHwZ1reTR9zTAFuiUYvLLjV9di
mAcjkk7HSDLgprPzRrA8L+2rSIckPQ7143TKy1/NdDFA5+Uc/liiacI/jjXSjPW3Zsiy8D5M6Knp
sDr/IYTtTHJuUmfSR3lTi64ekeIyLjgQvMDV6gLMLFfWpu2rPI7Q4j5WHpMFeEjY8ULr3UEKUx0r
+qSLXn2R5geeg6jmbZAake6DlrKFlAj2MrjK7tO+oBv2TmcC48xIcxoo2MDMHLVF58KnbE8eiDRi
ICR4jvwbIxLGjNmhadxqrGAeqhkRGK4IFFMr/iei0onmqjl0uz1/g5svKtIZxoTXi8pF0jLuB6JJ
BkvhzJoV24rp5UNFtIkpHzFtalP5Zv+hZH7+al4d1jAfxD3sWjMW/rWCXatnldMMJosLKUZ8bBsP
j6ZCin2t59xqzUz6Po8O7G7WC+3gOLuOPlXL/YzOgep28aEmu0S7EeIK7khBBLHqdBpJ7QpvG9zh
fqzqXm2YDdjWR2+QAatG+1fuI6xcy5m56p+UKBukaAhVQ0FhiohPUbAA9eu2cgnlwYmHhze1qZdr
dzn82Tg4pnpedhuMVZBB9naDSYpPIcElHqJnG6OdVr6LcE653V5bYe9Q2ygXc4NYi6G614wq2Og8
O51XxLa/lMR27T6fNkG4f7kjPvEjf0+Jm2GIf4qjwj5QZF5oYoxOoreNr/yOFUS/i2Qih7lwlMQT
W1N5yQrphJXE0u//0OhBXVwkodhzwEAoUcl1VVVYlyd/flN6CKo+YSVmp/eereZMpPTSVQebSdN2
5nHKDw8DuP9tc4PoEqNz7UuolChjO6INcCfk2UDLmVn9MJvVAsMyy/VDaiTONm7RkOWEOcZvfx7I
7h2gHxsdlQ/1vGo0lzq7lNaw0reKdD/jMf+hpj/+f3oqtJ1Z0p8si+i04i1N4sP3yIHFoOiwJyrh
eADFS6hqjhgRSHi2oe0md5bUyQ4OhLF5WZWwVpXLocul5o8KSkCIBDew+YmMJGSWTx9ET/XY5z9j
1GwSd6EC3l7JoBuJngT0D5KF7L4o9V0I2lWwUp9i4SkmzXMK96D8aPy8EQAbliUyvW/tMcJgvB9E
X2JU56l20WPYi/BZ1ScGB6NZc2HLYH1ieegVEqshidGV0yQTKVSXcu0ypXNz0aTHHn4qvetjKfvu
VGksT3gw8KgESuOzOgmIqJBXjVrP5IfQ2EKGiE7EmOKehygkAJnwyvraOAJkfyQgtFgA07zm1ovL
/FZ1YbT/Zhe4730qLIXyJ3MLxmisJTnqtG5qovCUZtyMpG/nQKKggnP4J27URQwMKLNsQEiyT2yj
4Mfpyua5NR2kmMbTqpeauMfX4fpCu8cnK61dmPvDAUCMMLVPQQht72eeV92+o1Vz9qcdE80SxHst
u2UoTq4L+P6RNztWHmwzU39Pa3yTeRKAMhOdOn07/0kAPWfv7Ibqjw/o5ZuAwg4irvPnRpz0HY8V
vl729dcRKtQxmgCj29/74MjUu2nrnY/pvclKgwF2Y/bEGtrGsYudL5DGkFSJFSwGui9lqfb2ZJ+6
35rxk8Hi7RA5X5TAP/YhZ20N++bgDUAmoUHkaFdJv7xiEcrwa0vEM2qnoogR4lmm4cjlE/4449J0
9t1qO4bYHpbqU9vxQrKWFtWKo9ccgsZgQZyMkF7fi43NJNFWtCQY7G6uu9MGt7SzHTLws8Wcb0p9
WUXL8xAhGTlvrSQUAzJkquOhIn5dGHPAP6CsOGqsfyaysLIAPkKhUSsoiBmddQVR0nVDJynITBRK
JQD+fUYSrFLg2yqBBNyP8D+KcwuEkjAw4zkT6lDsAYxbim4ZXrsY8A/CtRjfSkjf5V1s+wkMAxn4
QDtfrKSs15DmLLiS5rx4uhLQy1/RVpsKY/q7FsGk1RUp0GZ67KGt3G6nqeXa7t/UoaBC1mqfIbmn
xGjhe0ECsqfUcioyOvJs7KcPy/RXHuzp4Xxi3pqxd2xR9BrFkQ4dLRo0tECr4Pgg2/l9FvTq72pH
BxamYxWB9MYoBa1s7AufeUOkyg2o8XSO+GR4CWZFlcsUVcVdIo4amCHcnObSyf3VYndPWNpHjBRa
wbS2EWBivdrE748LgpecbbiGiJQP00wXJfjePwIL2Z02KVMlj59LuDINm3k6j+O1vzTDi2KSl5Jf
1Bink2TfLy9bJsU/XxqrwU2Y3sKbXjJP2XrOGWgSw2cebHhKg3T1dkGPUz8HLhQzQlPfSccTwx5z
8jXgwfEt7rNQWS94gO+46p12jUYIc52lRKwlJaMLAS1rm+Ay/3ORnCoNYoB5nnYUq8lCqaofFjZ9
svfvBQRvfF73GXCSOdg3WVfEn+rmNBmuTf7HROL/mAQUufk2QaEragXBGZSHeGWzaYjOmC4OQuK4
uJI15imdllFDrOCvbAagd5g6+fcDcVfH5kEaUQKTY16J1lWBSFJXzfpOeYUZ6dyYABq/Vam1upWR
JU/J+SXFkwWtyYUgNueTjW0xq9CXpzHdZNfTM2KUt65Q+Yn3Sas6xhvHoktxZ2AF+W5wKMctjQWC
qmIaGJTKj/Tq8uSyjyN0HBat+UFH5z+18dMg/OEbZwOttEdUiZ/59H+g2r7pxpjR8kOVAsEO2Umg
qNa08So9l7V3F2FOC743JXFMuLpL5Xq8EzStXbOIr9mq/R9pz7f8NiLi41uk9lq6K5tbK03/PYrt
d9pkBawH3tW1WMex9+arB/Nt3yHcUB9h2KqHM+K51WbvUPv8Ym+WW2wEER8mbpV9ZxH8PimeDNZb
a2kh5M39QrVmJYATOVBK9iWVw6HOZvUlvQ1IzFnt6gOmSj74HGJhTTpunBeKbpcvUvucvVAopVwk
jGrfzoTv2eCTYNzxtMdVfrsXF4y7wY4C5EH7pFn87zChPGPNp3VkJtAB1UowUwaSPap2X/AmoFzb
oNfixwUpL+R20IZi+nJxagiMcSbOzblBYC7fpf5zXBtp6xwR9bZEL92YedYfeypq2I9tmjt0P48j
P4vVW42tfG3ziZXdPjSPtqApS6CovSHu8URxQTKj+onHww6BBQOBsVrw9P5ZTAMYmUfk68pIGwhT
0JX9hPiQQFkRaDS4Lh8+m3S15uC+CLk3Txe34cy5ZeKkZkyrmbDOHY9K44gEyj1GWWNw5CFO2W42
NmwBT/y25YftxmVRURifWiHPkSnkyFLRhV6Srz96jjSWWab4iHeNp44ah/nd0xaRVlwj98KWTz5q
7uMTLtBRb1UsbWEQjoAweDtGaU4qXMrK3vKwCiPz3DiHVr8GiX1IyC1eG+1iIceF2dUCXRj26wP2
nwulgEHhKxL0Q5/g0ryOdW6MNqsvFJOuVE0qOIT34XM7HYUsxNbt+tkOxpItVSgYkWhNHYbfzJsv
spx25xq5FXMI6I6UZHDfTFssALba00HvZ4GHH/FzkjlnxGYUBRxGPiLXgY2ZUbhDS/U2mgY5ahyN
JGCVEBk0WLCfqiGp8pB9edwga7hOBPjb3f2nIMnjYAnY0iHfGufMSYKEpnV0xOOyzfLMbCvOOaiS
vxOKq4hAsCtuRzc751N71RnlVnDNLde4JlldEHj2tFVL3J4mTU2fZz0/DKJ8eZnlFv5qSxgHphMM
9q4nAHcVd29nNt77CsmTNBJtDzUw6nJl5vQjofpYTZ7pPjmdQcYKpZ1fF9bsTfn/dfuXklWw/X3D
iUo3jK5il8dLzxIK1/GFxE7hRfER+vNkhd2ME5qrKUWulW371KyKJhXjTFlDkMs1l3hVBE/iUFLd
7SiCYo6BtPyx7nmzke+O7DckHkLD5zBjx0Yy6X2c4MlNSCTDFNt4/rzXtx2xWFR9tpqWECqjG4Ix
+q1A3uDfolpfuejFWLWMy5ZrAwbdy2x25H5sK/fQ2dc+uwlq5ep2iag4jZP/YAJ8+rs+UutVo6MM
b8AwIXWkvob67yx/0TFVQwZiUNqhI3H9SDwfyBYhzWjccCnArcUe/Go5uvfYFYQ2L2gkenouYJ8f
CWDDj7fxdIIJZ8qLxBGOWThnJ+HAnGalEdpv1VMIEgO0ATGpcZWQVHlrsQtOxp6aC4IKmLvg46BC
4CuvpIPdafQUJm0x+Z8gcA9lxRXDvCjBxvJjKiF7G8t4PPk4XtAyOJu2Jf0hmBh6+gARvsCC2xfa
ppb5k6V7JrjH2T1YhgOZjpC28yWbxlGY9rHFmoyXeYd53JKbnMDZ/CZYd8JTz2ylFy8pfth3Apui
s5Z57279TXR7L00zxtLoUZ/nID1WsFGhxi7V2ww7jTmBMQtpINr2RwEZfuk5/yrk+aKdcnVcUu7O
oFMffk/3065lmM9s7ahMfgHjsmemcUgu8mgQATBjooNrI3obYWbKhGDDvGVvp8SyyuHd4EVgB5Px
2+Xvh40O6uqC7fiwFsoDV00Mt/AoQfj0sJkg4CM4iDjHTY0gC2CLnYnSRIsY7uDOblGZ+9khm6II
D387cw+9EGGNQL1XvDaq5fygEM/yUsx8yGjf59jeP/AcVYlWiY6s3gKKhRrtCMVJC9P0T8DSYOHp
kiS31KtIJ02NKu9qP6oLQjGkpTgVgcApMg/qnhovMFaYgUshs6Pp+6nFfhLzdpBN+KnZ+XQxJzij
JYvTZBQgw5lIGQu6CngCzhVhZE2PE2V7PdX2ebwI2yAsZy2JCmkPmWjspEPmL14IEF2NCntkLMI2
6mB3VBAWhop/Lld/+rVXhHuHIJZfAUeCm4LD+xZymfp+JvDp2YPpe9+u91FnTJd5DpqMMAoDCLRB
HA9cGFODuGEiJLuGLwKtAVfx/w4i9lYLyPjANR0QgGEo5tRiwv4oE2i5G3dSyNbrozrNIfoKur58
7RCAo5fi6jCTLCC2m+yKYVyosGQKZSRZjCyo+Z4Baco+380Q6iZZIeUbeyc6czNqGoPRNCsFPrLR
E6xE9AccTFauFi8P2mrVF101CghipmsQeQ63+Yn+0OzLEKwOI1/UT/Do/2hUfke+zdA9DSnKaVtB
yhAvfqZru2O5X7fh8bAnTwuJZknHriXSRx8Ny9FChzQT2BUp9U0Rs4e7GrQWUhhINvCyFvq9bzlC
fSkGZraDXniy+VdrLC30HQnSiF1yXQO6xOC2GijhUD5xt11yhT6kxR1DxivaNGjrMltH2kTGLovN
d4bXWQPttaCK3PcX6UR4VFxNkl90Dz6q3lYlx/CqfzrEtMBl6j4KYUvpjS7hy2555VfBiUmyG+PJ
4UA9NckEi/vbkVpinhh1FYuj68puooYq9k4vB9wYrILeAPZiAnGI9ABXAJd8X/wGKQcUsy54gnKI
/z3ABQ6/L1utKUjsCCAY/RiTPNMyc9gxXqdBU++eSHsWn8CVK92IzKtO1K5L1ieEvscK4WEWLaK2
3wNAQ9gBlpv8W67y9yhvImTlx6FRyXroz/8MdGwaMipyjN3ht8zp7VF3gAOCfFneWRvDow+G3AmX
kqdSOGeOwJfAKtP+gpG3KJTAUJbgLa2HHHAMJ64fCgyzYwe+6C40u/79Mwkkrub/JRRdqatE+OFD
m66WmTVlJ3umVLBERyuqGAlkDfc4PqUBOS/fG0VimPaZSY5REs466GFV2gQq9/Jt2AvUIwa0f7Zu
L4le5mxYNzupKvGpLdbewXc0s/dW9Gv/JkzKdWMDupafT649lnnDUsMYVVUuxxdZLWXnpe3zlZob
L5/AqnJSwtsRAvz428/pNH93xy8ZphZTEIC1exebkBJYLUDvjo4MhlWpDSIlGrdN1KDwUKOPs1gB
PSvr5XqSKXSI3aiGT/MK0VjiI3dxCRycrdeyPyN619rWgO49xpn8WclZ+DcD0C8RjSF6zvMhZMc3
ZyWhbcYBpitbkTY7UiqnxkHJknhw9vNiNNHlLi1mGjW+cxn1IL6s8z1apJy2iJSMwQoVGCeML87R
rKbYPI+ZRPhZJwhM7mzgUGcPCal6bJuYS0sqzslXZNmbsTybgWGYpDrk+iZWVvdDcsAV6DHT8+QI
IVIy1MZqtzR2aOOdLv1dnXnj6ndZLoqdeR3Hgk/YtMspoGaRC4Z5wO3nbAdTKNHXEMGWJUA2lIsg
OjSRd0uFml+/YkgQcRD9kDiG8B6jTTC4dFoNIvW9FN3sRZmR4vPmncQ7Cx5H946qizXzwMzTEung
2X0FJZ+Cmd0YK6suQgpGOzhqLPDqSXUS9zJAfB80pEnLj8M8DHNUs7Yd4nILbrwTKa0NFbI1JGlm
mAi60KGu6tYM2cK1bqwi9uKGu45X02iHhY7MwdSciCNDbU9//9F/xBygy8kl7JVdjofI5VMFK8lp
WhUfALJL0J0MhR4R5cLR1kzh/GQeFXKqIfOGokHy9raQ5tDJC/nChNOnvcY5eo1EXA15G1NWKRAe
JOrnS5GIKsZE2L3ZJglKNko611HV3+htIJ2VEueYbh6xB4B/jL6HMii7BHpOCT31gFOSiLg+UEPX
sQkBKbdrIt1Qkpf25JLB6PrS3ap+JLWv2mDXJC8SYPqNfgKzgcZDIqFB5XCaKzPBtHWkfa4UxQxL
T9IrTSWAm2t1cY3qB0MX6v+ATedhUVc1Kf2y13XrVGjxgqT1QZeOqto3wV8ZfbLGqdzWwl2or3b2
t7PSXseCw3NXhg9QqyCuYqiedl+bcyCIS0wC3ZCgRmQ0zh+MySBh5sIEShp+J8HA0xdOfWWoMppu
CvAQwK4QzgFO1kuA+LniKkE255CdVTTlkgA3mbsw9A+MP0gjLXpKqmcOah96T52qB9UJ+cZ3F4P/
BNvJqNBlCQvdog5UTHGBfPX5+k2KKlKgviAwg9ckPbQOkl5y15JT/KN//JyhR8mLfWOwPt/JxaNZ
NBovX4S6len7p7CO43Jrao4jpoZvG4J7fr0GMvo/CyKgmzdZ1VlL74jyCZ785JgXqfPaNVpEo8x2
ULF9BPv7Gf1LBW9MK2+blNjcgOuApKerUVEO2f5SiS0rjPVPTCgeepzK2vTSZHNcdxDx9ckp/tz0
aATXYSxYGNmQJMxouIYKPgTNL2xdSc9Epy64EBVUmpP9ycvt6HOOQD0dhb8zcAcyTtc1T4fvMK/u
zWav3HTqyDqQoEzMjz/0iGdC4YhZEnwvi0AeAKEk7OhXP8KQfaL299+UU1yDRGfG+N3ESTHavQM5
9GgR27qdLI6g2k+2D4MoiPziYLcUam5hIq9iUgLCoZT0IQNsvo0KhrtFKnGFlbxU8msqb/dbWk/h
taX8lucM4df3XwSaMvUcY4xv6MTjo8YPWdRtQpdN4z5TYubkJN4nMS5A++vbDMIodku3TrpkpDbx
+8XefdtO2o6ljzKhyg4j7jaB+lAA5wDwi7BY/PLiF07hlFkVp6jnlLPvKkM6DS/Xwa4BfdUOXylh
VpDnBulXXBa63C/ZTYBiIccPkdr0KnYhPgyvl+inaiRPbaUie1e+oUlTMROAaHVwfdWCgAnlA1L+
1p6j1sLIvzdfw8Yx2UfVVEjLHzeK0h35viUCSY4cLvxmBxyJvoIcJbrYW7K9RM7UeTTLkto/oDha
gesmI0OhI05/mBaxyd/4M6nWMlCzaeXJhkh5gu66HJLh047TZnofTU5bdY4SOQw5pWKIAvQc+ImD
dDLbXyFk0PqdFk1JbUY8I+HjxwbRUZbNwDVgQdcg0U85Ggy2lCAtpMhrukdt08boxqkPo1lKZfod
Lj6OhSzFpsBoHsLm4J6EjP/+P/qEyWyTzTIHkin0Q6onMmzlju9DA1AeAeZ0wTIRYG+qNEX5zvW+
kXLZTZUjUaSr4UOTyZLH60Ei/BLI1AcYOCThJHEMSYLQrxkeHxxKYxs43TwYYyvJKBeFBVkTS1nG
E5cxHwkBRix+pJ66aepjvJbKYylk76BkBvmjZOf2XD6c0n+kItFlheVN7TB53jJRwRM7bsV5nrAJ
bUsgOkOr4FVSoOmHzWl8FO7N8mo/Y83NP7Kq2JVMrbhYrsiYVuBKkvh/q4bQueyKPzHUEK+6vGWQ
GbGwF8XxjgT7xbgU3A4jw3cSOmghbA9706jx16hKUOvAr0ugzl/9SUGyJRpTiKgZ7yuo4PSCWd5/
R+W5kLlyXpRhj5BPcZkLE4HYk1/b7I5YoTll4qBYcLqsNqiY99b+5e/5mVCLYkIDI77E61WhiEJX
yboQwGn3A6DSfbv/qUJr49EC/fZTMyR0CYlMfE/5Zlcl1ljSB2GFg9Q6KRhkNESf5Dq1bFbcblpJ
sLDXmy2KFannWr3zfIwrkqHJpHhq17MByfMIRCp3v+9vOhk0SirwuaKJNiLEJaV8ThEgqpPBRhKj
HIHLp9eMWg5fPGvQ+UOAqgDnFl2TGyMDLQ8b6y384i2nXgR05YxelO8ESQ/wC7Wa8aVS16S5aQJz
AbY+5zreElzhvn2S1jny+mmBxMnWDAcoWarMon3C9LwWuqkBnq4PPSdMYDaIlhtdofuLaz2c0JhW
pGDJLb4qF8Ajw0v6KVS+Y9ru/tHToNbFHg2L9MgKt9x+h87N/kDWgNkFRxfh8cs/mqMpvMSWroD3
pjbMsEpJQRAppT/3uT9nHYKpsoLDOeaB5zOGeljL/KpQtolHiv1XLAYNm9s1DxEY1We/9PbOQQV3
BlOWQTP4Axq/bgcZPl6S9iC/EP7X3l9ERzO9CN7YHD57uaS+Zz37YO3RC72QxunP902VlfvWzA2f
ncuPsANET1Mr8hALqINYpTE10BAQ0dS0CSetaXCJKy6cgbWfrhQ5xARBfZJmpKJcGzFNImtnEtz3
cT/RKZl3bhfFca6RBoUWee3AbIn/SgCqibevDeygEezA33XfScsn0fYnTSS/tpUOB9jQGligNcGl
E4IfxW0+5DQAQURQ22g+utow+RGE6f9MKrw+BxbeRF12gAGaS98lic89Gory1rUibb7X4trLrPYG
6pFZEZhsN/9I81DgNy31c7zCU9o9nHqAQSTlh17sq9E9uC6e1dRkcJTZbcJ2lWGQvWnoWbOz/Vd6
pjK4npwf6JkOG6/xu0889oQMnde7wSXdHgoRxaf295YMakGlejYz+/GFQcHx/TJZbWnJBVhWBEs3
vMKY7+yk01aV95Duw8L6KX8gB4B/ZEDypmfZXsXjrrs00kG5PTap8RyNS5mNVCKfIRtGRTlXPd1k
OqC7GnhNT7Eo0H9Jp7g7v1V5MYi0LkMBxSRKkx7ygXUmrvx7p7SMfVJhyg6Mfuff4vDyv9hnqEHj
yh/aIcETxgGdGxXe5Urp4CWwRZYTbrupGSyw0pE971mDHYhfG2NzbG5ZxTU/tUqWUST9HUwy+g54
Qe9e4Fn6Fx8SjJWCAJ/iBzveE5+/lXOtaqVLRC6tgZ4mwht3B2/hGJ1IGnTu8VHXJ4++qDzCYf4Z
qne4KBwZ/6jfeqZsEnVIJE13jXuzFjC1vRd8ujWmXVNlBfqNnKgEkt9YP6LsWYGYQBKFUhI8pKCE
PI4Ra4TX7T/uT3YMS7R999S3NPq9WwyckpGKemKAZxpgWT4N4pJpn5WCLZcdFJgTC3SXMmkPSOVJ
1zalRVSqTHz+hzZJSY+VdmkFbEeK0o259UF+0zUkgwCdiDOA+1RXWH3JE1WcuPHLs0YR32e5HZK/
PQMk1ciaHDl+Mq1u9XJU5QXzm4ZOb8HZGlYDpjDwlZ6TXhbPBz5toY/76BAeN71CE69lZFAKKKKw
gmVDRLoEqOKr5lhnuJBJTuqUzOOcks3O7ZxRyQsQLzw3UWS5/9jo4pMluH/aTrRD3yjLCApDdXkh
3YRTdt7uF9EZrocatEjpX1AprwI2F9FwCBpYNlRVvUeVUDkAJ9KvR/vztA3W6bgNdngmfDwf3miy
tqnN/MsDJ2TfyeZP6fYcyCoBWKTT+6bXpnQn2oizE3nNqJulEbNiHwiGFV5TIPLeQEAIfkOL4gzs
tooZRr9SD6Fm02zGOs8J1BOHW+Hf4c5YJoPDdHuk7WYZiPva/YbX5d85NDeLdN+BW2jysMhXOoFK
nGQa4G8EIYHBvwZ6gRa1szwxLwYhLwHcFTMWrdzUHJmDO9rcRgx9l/NNppKWGWlAPXlyYSxPhV0k
1jP9wd7QNUMQyr+hyUyE59Tf5yq4dmFQEXCUqepxOwQFD6jztfPkkUlyRumNoIsGrkKKLcWBO+R2
qYZ/GHxQ5YXdqr7aYXqfFu+fgJVslP9HqbChT4e401+1+qvh0XIfiossUaMGXCs7hppDK3qXYZa1
HXrlmD1rvT5BVaZHm4EUPVo9e1IcXSshzadT5GQRlr5zMbdP3mH2cBheM6O25/pQahnHGWirz81y
NXuPaDQuL0VGwEVAJmOyq3rjeNg0O5MRyjojG+HeoNkQyTRrcDuGZ8K+eo7dgb+Vl0FahCrcceKx
nWZg7zTu4Iw1g9RbLduReswV63p+Ysm/J5ZuxbiYqat8MF6xnl+J1XEdwuE9ZmEQvmJAg55+rt0E
sivnDbKp+bAck9jZunC7fH+K7Y/HKUp0ytjrU25Qs6KYvMEOczjQoZHMf95kc9/iC1BQ01n826GL
hCR/sc6Mti8ydJ5yiltX39/uAQDz+oXbywNFq7nKsJrmbyyXNqC7ldgrXdjIbClHNb7o7zfDE55+
QoG4Tv/uNTkOUzzHHOkzw3Bf84cdpadaFwhBQeREH1p3wM30QH0VwRq7qIIBet9EEcyTP8p3YF1b
iDQNH3mYcZ1r7GvOpIcvpkFErTxIqJY1h1NTsC6CSDkgOaF4LkkHVGnbTun3Z7shomvHNYvf08ke
fnogNyt+yBZ/AailNf24cxAKnZhihALhF85kz/ErWxqNpjihoby0Qr6kD9hCD+FvlVQK3E8NgfTA
6V/xD5LLs0PG1NEDN/43Jg6r5BP8JD45VBwIa3a0RhrA/GeSzmu4JTWKqgrWz0O04VhGmd17Ij2R
Nk5GAoJ1OqixWWRIWxmMkbOGkSOyEAZwk3ohoLFLRucAkueVQCCn7prWBiF85jC6mqGKA1jJazGc
1TQ2Wrivj7BKJnRDJ173djq0g4/gYeajEFAqrsoyefa8dqTMzckJ3Q5QFA6DpQjflv8ahwZn3BAT
p5+r88xxdmdoVpGljpMAXK1M8bKC+qstBZzgYUxP1KxSdjOT6gtkIk2Lf8ri9cgB+1yFFFLuvrDR
OdE0y99ADVGUbIvrRxWdvovzS8yk6pttbBX5/ticYRaNeXuxUlxbp3KLvDcwjMcc2Zcpecyb83bh
l/ccYw4nN4ZGUPaP7iUSomSesT9HSFJhAedMT8TyQ+UAKxPX87hap191fLnSp7KGe0dQLDM0AmSX
GcHSlFH5MR8OEiqEGbtHFMl+yALrO1mMrUlsDwwwQZkC4BLoNIYibAtUhdji7p6TedSj4CwJClYv
ozWwADKhNqVTTt6TM4Y6M55M/Fgf6i8TIIbGae/MTuGloUI/uPCV1IkNZcqcBcEF+C1xMlD6tosn
gjOyEG1uGlL+YPbuThAS5yZ/MINbLVquPCS9BBso3OK8Nfhvfe5kL80bOSWG7XnVQpW4pVIgOA2s
ZcQzMNECih9E1CT7m59dnWSEYjRI5z7Ss7quHEP1KjKo0MQK/5hVZVLshXVU7S3G7VRqcNpkOT1j
l5efQdX53KhSkBFoyaVaNhHhXXC76JKMkWArVXsZYVCO5tQPVz45f8vcY3UVKEYaNBo0pb+6GLqg
Lkzvt5oEH4+qEpUTLOoCzab7Wa4UIAIseN5PS22MIjFQK5eSp046nlq5HOmbxINVr+S88FFtnlNQ
0oeWhpQwLvIkHZJXWQlRkIXYBMw3tTFCF39hVv9JcmlDGrkX09j9ODmWeDxaqkPys7VVfMlbgT74
3WALbFl5o+UhW71BvOeQQfiOq8C8jfnP71ddbS95AkQwSRFOKND+QjWRCJPdnfW75ysammpu4dQa
SlmCgTdXk0OY8xpDlsT8BZ1U22Nsm8ivz7g0jPY1Hk2Cr8lTd4mGxyVLJHozEtX6mVslslH776kt
5Ylv9c57Vomqtp4N2bLMSXd/n8GlsFxM2Abegflt2ifJ90bbqmmXxCSFGeWzHU2N8cP0tBnIga/R
dYc17ZtK6yMoRkWTeXRO51v2cQMYvEqgr9iihC796Ylq939EFwPxVmMMbFJ4CvbGS0+Q7AypeiN9
DERUZ7rWyfMj90i69MbQoZJhiFxFaYkrfIWtsDiAxT4Nxarrh+wTGD2aSciKkuJcPLs3zz6cfmWZ
y3OeKlEAtJL5x3fc/PeIuXK4olh8M5uhLsRl3lV9h3BTQxIkRZEy5B7gWZZsnJaWVl46iPSXUKri
tDwb82Y0HVJOiDFT8bu5gNLL0YmpQAa30EVUqDLCmVE2dwDYtREyx0mdlurPLak3+O7QkkEqcCad
9qpa82UQ9+W7s3xI20S6QJrrDtbgL+4aGc5fVOb3p29JLHmm6sSH2FL0fVoyE9oyFAVZuAVzBkut
gYeDqzuMoir5C7sBXW5nxvVBC60cjnR+oclV2LAyk6thfx3IihtzHBQZEOyhXrluJ0ZkTJ2KaQ/R
7gLJ5W9XDL1doydWgM0t1KNDyzstc/6OEv3YYeDIBrXkdd7mS0Qxt1P6z6xi/UoGkR9C31bIllsw
B9rXaPL6Qqd9ngKbn9agThduu9+D0gbIlcCse9fkhXazfyEPImbVYe6vo283AZIU7tXWoUwYWWnc
v04tMjtZ8acGD+Kc/iHc3+s0TnPAe5Kkru3bVW85RuOE+4LivwxP+VePJz1pGKx5RR5D04w2QKXx
fwnuOHlHEKhZLfxDwOSUYdghonUjgs8h7lM11v82k2uyKN1HoKG/lbDAVQD1Z2IT1VOiUl72/NqF
tWLpxSTGJDa0uNdFkFpSHMRS/r7VgMMRdhQbIXsCgA153H6jRM5EqkVF5Q614CHq/OnNWwpnf+QY
4VXM++D6xjcNMgccuzNOB5864veO41ksfV+SrBvkyZf4Z4n/7gqGG3kyp2bzTGU5R+CobVv87eW5
LR/v+ugRRV2HjOOEK6Sy2yKDdcg71R8VbWbQ+MvR3MsFnQvukcGgV913PlVNMxfncQp0L6nVDta1
rq9Q4thlyiv1zHlJxgaISHgG1rVKBs485IpVOV+Sfo+5kMRlhD0JB+6ZxqXEPcyXdC+z1EvZc4dz
/+U2Udf8MzI+iop84I0Pvx9/XMis63ty82TPGJiNJv4NovBG3ole8R7Odfz0ZTydoS/esfW/vqIp
vFh4nuEDsAIH1CHENjWqEZZmgBoSQZn4hTyDzheaWI17tU826kZa/otpOFJxseEvdRI6eu2GW8eC
JqRJkPqjEbippZOX1Qxmhu0VOv9OQ0/LVv6KTl+SdjY1VqsIdCO2luIAcoyTnqneyg+jAG2pM3FF
i89yZ2oRvRX9yRJqorUoIa4QwsmLfbkEb3FLf01LkgDcH9OkRi4DJdUHcXOjYt87i7O1GMZSpnTg
25ClOKCF/fE8f15bLuXoCFq/widAAIf++yun8s5S702Y1Xb/Wo2KyeztZQ1NT/YRU7WpsHG3eegS
/oD93GkC96CnLr2hMzPnhWmYgFd0y35sM7e6E1GFs5qPcbAbS0qIF6ilc5sSdQeW7BMgW+d1gxVp
IC8QBAnzcO2Hf0tWzNepx3+7H8+zLcbpOUHlBgcUDTzSTKac+krJuWXrmtrRwYwGnZAtBYj1FMGi
b099jcBIdmfA1rpOrFbRvsI351lzfIdJoD06Q8dqAhJP8dxgvLDTOXOM+Xk1XdgeH2tp3qg5x0BU
rODmH4W1WEycTv/yKQBbv1amZyJ2S5dSserjmKuguZqP6qxcsKg6LXS+ByKS4Nd7B+hi+OPw9bMz
w2AIOF68A0zZxhn44UEIf7h56QSKZDkmd/o3CBl5CdeUdpaftihZ4prUYgfeBdhsd8Azs4ZpO+va
+RXZec4vhwBaSyta3h74+RaOIHBLojrP0x2jgudERJUC/7ur9xOlIBy862nFSFE1FrA79h0gy4R9
tG9fQHd1p7WOKsQJWHadzTfQ6cdL9JeyxCQREMODVecPQYBKrtLo0t7NRIHQAGdFaNi3oyIhqvo4
8GDAEsMhQy715iDvSP/50UYTKQVCaOfNEVe2FD4LWJgRaCzwIt7Da/uUstx4z+ptilBAfV2fwLgG
XyLIdZRlxGEDsnG1gdPn1I7yM5g9/25Tqq4m3O5TAYrdB9sTcoLxNeI+GqjRI/l8mpy0z+ob7wlx
+XqZT7K7GFmhcI3c4Ox9vZHwVWlVkCujjIbdMK81MNebEKdkZtCcY7tW2B7WQtl88R5UU1RgbMuc
luURYfQpzU7H0nW8SaK6CKFJysgOOrPsyWTCSdfM77F1w9Vh4KhGmvKPbsyvmJpQbIlVncX+Zc7G
+BW/6+k3G+3jz889niLIpnIFME+QP/vzxdmHXEceuMorD/1/roO0+BdK640xjZafypwrHi2uhS4i
d9/ZRBV+R1pGBPc2pUpkGwHz6KHFaRsUqLL7czkumVnzVqRvL06Riu9OWmh+eDBgWmv06RBDe/HM
fhKuUnAMP8VT1QiGImBdUZfv8PedYB7z7XZgd00UN6VZrTwP9AlAiVzC2J1MzKCAkhQbusE+AGyr
9gZuQ52gV/Pu855rI1A4GB/b6ik5PdLY4FgJWGB3Nl79J1BxEjvhhP6mKt6VS9HE+65435VyKz3D
copFt+aJ0POd/jB91DrGLJkw2e/jI8shiTRjWbfFMr7y1co28vu9GvX5qpYqg8XRjwlEmixs6oxR
C/Gfjpmc4JKl23jBo3moHvSEHNTe0ozpomN4nDKwRpmB7XWuPZFPY66YNXRzx8FBSwM9Faz2zDG7
igFuK2WSVViceAGLFWGlRhjcozyvpYxKZAw4K+9yFEoT0upEWQSSzXylfn52MvAJFSCCBx7U50Nx
ao/1i4pI2drt6UtA302eSX9jQGzhx/1qdVNxmF8rCDQiXPl+myIyNMKwYn/gIJdK2JOMVABoM2zl
4dggnlb3xErckqStU9C23vf9j1lcFuvaJ7qTWpSiDnvSVfgQtcwyTsp+ad+s+VjYPwqkk/2NA3ih
jNx6mUPFSu+l88Mobwddgj06D+HQ/epZo9RaUXiJScoYVB5nkM2Q+uiAjBZPmRzS2w74M1BLsXkm
GAoZyeI7vbskbprN8MhA+KTKUu1lISQ8rWmzqmIMm2cno/uNIIGeQeeWRSvCuVWOvSU0HcXGD+sR
ewFSC7Gu2tib65u4iF9KMFsjs0TcPGT9MeAAWsBEp9usuSXZlJ0OggX1rW7jVY+FEYys3M02aXjG
OcZYnx3oyCKZTae404pd1HkVtG0kiIaNQORjsVuvaFG0pB9s6iYjWADEH9xtGsNt6J+yDBeWtHdZ
ka5+0MAkspf2FlybWYPKXDo7zefwPQk15MNe6QZSYL5FTotVfk5fJ7FpVHoMIWNePXkIdrOF7mWT
C2tbT7qZSynXC0fyTillX4fX/ru2lVeMBDUN8eX04Yh5nqYjTA3K4JKi251RGbY9si9ZuNJHfDhJ
8V6WTPs7uvqzCLpNWaD+FBrZLzBmN4GwgVGhhAqgQhYrJCREwDqLIa5xvkZHYFiDYu7qAYI+Trm4
3sOoaPnS87eHQwkE6Zh78xBuaVAAmkrORhhO6Nsxdhmw9KKro3XGdFUivmOVvTyl8321RfD8kZMR
qTj3KcI9dpIR7+kpufYDoYqedbqmQ5nv8nXAPIX1aHf84d8rIn3Movv0Lo3gsMF+QdohTVdnnJ7L
jwpm/w6HY7lOZq9hW8n3MXysBe2sOjD+ZVLt7fzhrn1elaCkvsvvYgj7lTooN72EvkEpLup/mK75
el3DzGejcj2d9JEBR6+umDiuIIKJaCGtcKIprIIytWIlRqi9BA5W+hTNFQx0TUC0kXen8Vx3F8Wk
tiYwefiRJ8GmwKMZIW+0iG90+dRxOxkpbQjILhcZXBm3q9oObeYNOO3OiXYM9MYLV+m2a+685MIG
CMZC3Mq/DjWA79ih8uN8yvxjB2BA9AqXx3fBMDY7wwSVjK9RVc0Osnt8vasjgoC76mumwQ4fnXDZ
oVK3kpaA08uUqh4BFHy2l+w4BhEVay2nX3v3+qYCSfOHLUxdy9mwXvt53CW0Vrk7Q8dyrXmeTX5O
2d1BM/+GQp35/4PaqNeXeWNe7viQc+cHpAxjqsSQJX6n8TEqVchpQmB05qeBMtFqqoLFCEyQ0A+K
d9JEi88JH2qKSQyFbbe+ky0toQh1ZlHcm+ZJfm+F52zgoW6sBkFjKyggXXUhW6kT5wK7xKX2ChKw
GzbPSYqG8t8lsIwG9gC/Vo9aD5a12ew/5f0OmP2YO9LkYXUUg+f/+nmz9PINJqcNo9qGr62fuXix
vvSHK93Kz7YQs3gq8T21VtMtvmZfml0BErhMlQomXbeUX0kncdDpegPhD6gAIaTR9aB1yBPr0yc4
cSXYi+UHJV/cK1WofgCVrHPFbOJIerzrb1f6x5mqeZW5GShg6P88TCGmMHgZ/SGjlGaM+PvvnMT7
o/C5XsAcZZMVfuwFC8Fw5784a6wC+c4lkpylHi86hGAZZi8F09GZewR8XId5VcCy/dsvWQfPqK2V
ue0uSHFRMU5WHS4p3qJd2rwfmCSdAX0GZmnWASVHNNLj5uvJxPnAlINQWZ3XH+JuL6pQhPSJEm0n
8tMAiN8hL3+bzYdZR/bl+/dEQ0hNVoeFPlfEhHOTC5yjJB5JqwnyDnWEzQHlnbI/NcG7MsX+C+bs
xHCGwlHQQFlT0OrLSt92ZjkTTfHUymodVSo7X7I770uH2smOukBfQW5BzjD/o3SMrsJ6xo2ug4w3
nK5mYlLZThf/dLwmTUodCA1xYtcNPjqoONnPEEyPddYUEeRtumxCXPASDWi4MB1g+yY1VwP/Pv/w
13wtJeRNjERGNagnnjyKXdb1SmjG/TqI826g/VEFWeBMRVwoMsA+931wd2hL1T5HTgpF228IQFHe
ZbvOg6uAwETJ9gjnS01jDuYKPVnMzWs1dnZi8jNGuUKIPjpzPRl+N+Pr9Vo7OfoV7GApGYeNUxTB
/LrtLCjM8m293SMHBJ8f1/6n4/eK2OWRuO2sdqmqK3FO3z+BOQ0aLV5nwLfdtbnGG31cBZGuYEb5
/HvA4To/u+KDBFijL7owsQdQT6mrh47e+j7uFIgxFP/yXor0Qc92C2DC3p7cGjhgZjJg/ZR3+njy
zrpOXumr8eMswQF6ng/wXFHhEKFtwmy55sQS2PtoAnZ4GONQOJGehE1k3E2vC0K2a9Jtkh6KeSE/
GhOKrfNxrEGlhLiYEqNFNydxxtc4ony1RG7B6sU41R6muVT7Mc0rK4+7clBkdXBbUVoN8LDgvfYK
MvqgC0i87HczefuKBiEz4jLhKJM+7zwAiFptOAzaeirnkF/srwLDwTgOrVUxfD5IZ3pRm6U0BZmj
sYZDY7LV2j+mvA+cZUl4XKtqFAUi6iH+sdzj3jpliutx5kmqXo+b1OvwSDRx3m9pws5K+CnDrtHE
5a5HLLZsJB0/smB/llfFx6wvd8MGFCf9hkmpsAj8q/2nWuzT1J8MKNdpKWXk5Vh6zvOT8AeBcon+
NlKVDPc0iFpCvYtTmtawC7EtGTuIKXcH3R6PnQSKGG1ibgjl0VTgOM1LvPapcX+oolcFfi4R9Mf6
dWCh6zodRWLOVJtjAmkes7oFiG3BkH8Y8M1sGewISxT/c8++8lxA4mmUVqaE+V6ORTdQWwLQWnUw
IrQttuFUPCnbZfuFzzBGjhWH6TF6DegUq2FhOA53zqX/C3n3q/VyvEghMMwVwcf1vj7z4IFm73fC
r3ARgwCr6hYPqsh2KyG9Bw6yFsAjbQ7nU3FZ/bDMkpn1bN61SuiIv99zLBL1ReHrHmFc08QJmfCX
WCoYya5ITXYH/2iMtHZqUbnkYvnYKlUoyzj3phm9PEHeO7GgWyVMJuekzLN5MhcP8nubimPohR/h
GysP7Uz+V9KKmcIsgFjXKI/yvLLtqXAwUcpzBGHPFEpOfAbdUWpUUy0JzK88OoAA5celI+YAQR+U
EPuGXNR8Vjl1G1neIzBHvJ1YEfXdhISJf/xbip9NA2h/N+YmAL2c3n0VzqPyEPRpVgmxZgtwuX5G
Ns4SFOlIvIzoS5dWQ9TxLm8AZKtVnvaxsLTeR2Ba6bzdZpBzKWYRN7ljJOkt4Gk5CdkCVEQLBRQQ
PpC1D5r/rbhwEzGmMWXMzKwjC5WBdORb5mYHBdVhnpOVlD4IxellMDQNunIZh07f/ejva9qIxQ1+
1Wvx/wRL7xG7WJWXiRrGE9kxSOzXfVXtIECTbDk+XYYV1tNXkbmeieo6uOpdhFhftcbMXjLavqU1
4yyn0R2pz0V85yTvUPnaAPEN+A7l3MWHy9tf87Pf0zcoeAGLOlI/lOi4C+DwNAGuJlzgT46sNou/
HeQZsM+ceJr2JaXWKYYlmTD3twT/Pfn8Bi5Uwp4BqUSV0H9LUi3cUdt/RhNdjWlQO4zUtyQ8zekc
VMVNfm17KqvOVGDzja3dKfT+FDkGRY89O+yidk0Jc3cwpkpSkhZI4goYSd9S1JBB+ENhaQS+JwCI
a8UJVkN2qUqrUiGvzc6AVOaKTDT98otWCd0dg5QkBQeb92jHNCFEnSAh1wdbk26bnPZf3+/kp1yg
NRLFZBs6QMm5ROMs33pYyrI1d7/ZgcIbjn1fpujfzAEQKc/+OCSV2sdss4RmFORPumrwYI/Mep35
P5FK6Lyzn4woenrCnkviUTMFLMiN5KLfKKkyyHl/x5FE29ecABTLITfwsRykyf3CeGxEX5sMiOPt
1tacLiS4GN7YRdn6LpyhmXoughDIU4/r6Pp7EaMGiuPKbvfSjJmgjocES/LbIkEFJF8aTeL/ZaRe
dGSoCLh9oWV8o+eezyl40MLgh23yacFBYgQcbbIAQh5VHrSWsCvVxjSO24Q9YAip4b5I+43WxmvO
y/IIszbVn3nIX1CS36ZKXko1NtttNrlmV3KydpiyMT6vzvA4b80N/cFygtbDZ85KRCK98zmW6zID
a2lTKsxA7LbhqnxFNewVW84IOz2XehqGNN6BmMCVmvHx6yeu9YwAJspfj4tHaSLv6BC9ZxZxX5bh
ESYeSxfAWGnLmCG4kocp+wejP949N2M/mqfaLEUlIBKP6NCktyB5xYOPTAe/GiLMYtxbystcXC4g
GSiqtVKg1xErONdHAkNDv9yNdOKyQSB0mDFGoBbgNDNQyOekoql23lYzamA7RvwcV6fqMqXisEcq
BzlSD5PHvAwtqFRbSCIYc7p08LKCyYSHVUzS/MLKaVAR4lulL4Mk4HVIiymLr0rp/fGJfeDVCa/g
JUyAp4FdBrA7B3hrORNg4D6BlQR/kATrA4LosrfmXjOClQhT+l3d2M2rupy+wETqIaM9YIsmAOk3
Vl4VY+9l9fyFmKAI3Qorpb0L0Yj6i2USi141ILxTGDJJ/F+wfE/SAvlXBC2dSPtRH33ZjfAACSTO
KPpOjPU07o+msxY0PcF6NL6rR2s5vde9bZ7nO3ycqk4LtJkI+KcLublrUaajuk8CLrWS1D5T2z9e
3Pm+B5lTliVL8IoUDWYja8ftiScU1PJ00q1UlqdAfBFw3fftHU0nCJu8JWEMZPIK8LmB2RYTJUzO
hbLcR+zBvl1DuQPo5zczzdeUpDi5CoH2/tNyefBZzPeNjjN/rmZb4GFI4+3UsM+XvwPBppoWO6qx
7B+0OIZaK5dYiLKA1yBkIGLsNtsfgIt4A1uo/HPEkdIVWb/IxVg1HjdrDFiOVRlAMewEILmPwp4y
8FE7bkPnkD0dRn4WoRuy3vzfGn9CAHcDMqZSvDhmgf69zDxJyiaV5Nj1IVZKJ/Yw0uvSggXh9jw6
e9nlv/+MySh58iXnyUqHT2NCG+KbCVo65oNLD/bn5E5QPGeqOInC6mpCkagzZmlxJ8MjdjSQ8bS2
hil4/9Bu7RhLbyKfOWkxAetNyhqGerWBNwuxhXLjzsiVbXOx6ur6FXvciNmff6bKsJKZ0NYxPGj0
wohlUCufxJGTJ3GWZOeVoI3XpMSs8poyqHCHRezIcfPSa/Kjo9F52kF9Gf+N/nEezwNaPq0BAC5y
vPRKNGTHvWDTVs0cG9ChEBAjBP2YTRylKz0u1mupZp7aEkHGhuKFexmHO3FZXvoUY2WDJJijh9bt
sX/OYS8vS7uLrxW5aKgKMj6nQsCw2lv4pg0zvNKSlFKbI4//TsGGgC98eZawC4MCYlRSbuVB+Ueb
m5PF8KxUvYh6EhRB9iudCuzb4r8FOE/8QjoDizdk0gBabIYdHABgtSUlNCn0Nd7PgrHbUeTtTKD8
pCSmvAlsWWIX/ukHkPfteHQBc5FkNLu5txB1sO6MLoJ5J9ABlD2nz07GtzPalNG/LNPXtb/RYhwY
aMKdNfPqc60P4epwfOvs7Rab3EwRB7BUCo2ee9cj6rO3MRioYuwdm+ZzFHtr99GIyEGYWiEy6Gxe
f+q+iNjk0dNvtWuNwKel3t+17h93GXnGfTONohbhjS+rRJ5K9kvYBPj09yUrue+LcjB97ocYBJ2H
z6UPk5Sj1+yORm+8YYg1lgpr1V3U7g6VfjQBRnqeRJ90G5XHtdT546H99y/rar1Nxj7m1vj4PGGg
H82ywpQTbXV5gGDh99r6r+w1HM32WJse5YLAyFkoCcTPUkw1WTR9CEit7cfMqnTmAMhCcy/OHSzN
awy0J5XzmevXJHf6XSMfMdyLGnAJ0DjDck0IipNvTVjSyU2F00U9ejL4AV/MjtfFLGGekSOfWDS+
s2Pdm3jzqRlIZbPh/qDT0GCd/ao9K5VChSVj3o3kg2b93mraNe3GuTb68p+QUDlJ+NMJ1N1nhXKe
2QsNm5C12ReeuGh38AxRb1jtYSttpNExanUEhoW8S8A+PQSUvR9RnTdMXt5w8PMQkKnzJV+/2Nm3
dm8ECxQzGoyM7waEJuHRutw6gC+AKy4EzdigXdl3cbJ51fSj2w8RbY9KJJ4dzZJkbvielGsvuIkC
h+PLu+7NtwsQ/SrRfUujzUk04QpOSaSPNRLy/q4mV26pEhUaR6QtzTAxwqHaTpGOkkss+gPIc8hY
BdWtwDAKoBwbvoexzeX6gYcc/Bqyi7A0Uysjh6jkVPNAqFGEY/xQ+mwNC/JxVnb5THxst6XmIRTJ
kCjB4P9izhx1eo2xKohMmyTUaz7SVu0rveX9gG7SlFFm/bXyJfDzlNOTTLITDpjrnU7pwNfhN51d
v7VGd9lHGHdrc1mdicuzawTKGN6OAnJxznouD2iaxyErM3qVo+LMKplMGmxIKSFZNCXDjtWoxO40
Smkwweph9l7AcwLYFM5dqoEoIHVZc026ZCckTU0bniGGnmxfFv1qAcN0baCioFiR6prms/yFGNtl
jeODpwXBp1eif2pcty/6hO5eK/qUdAzjFXlmXWnUgnHPVwo/WRbPQFsocX3KD9sXSSnwhK+JxhBe
ZZCuPDytaQeThR50TSzTRC5PDxWWYvBkSlp9YHtJwFuQaEif34ulJNdjnYW+ZTUc4smU6rTRYEvu
xfYtztGhGPpysxGeImFmQ7RqM+o2JBVoe2XOKEqvaPpXux5wjf9S+kA5jWi+rizgThINT2AQzqJb
/1tKdb8gtUgMpNOWELMu3xgo/R7kz6k2fIjgGKfv88VyDoDBW8+v98LPr/DGnjx5nirPjbRWGKl5
11djgHXUnr7R8v9VzOIoOw1CYWOVf3tN60XhHGXM1I2e4Zk7nsljNmcdTklwukIzzxSFgBlUwMQT
f9lRtaZklkPU1T1Q5UQOEzQPbN+VIxO3hzB2CUfq1aJRypGGyk01ZyKM8AA/qA06ECi9XTtSO83+
ANMP5xrXnLiPwxIWGp1BUdRunF//QlGnAcpuFpohV4DGiXa5rIUZo1YPBEyQ0hio6/85nyczirIS
hiLyijzsu6/UO+m0xmnSGUB/Vbe6lojwuwkXq8gLwI2tZ51G0wCsPB8tPTsuhlBup/aighNGvwXR
rCJjJRXYL8kt07KFJ8Wi0f3YeB1JaXmEy6HigXyNVzPc1cSkMsoxlC/MxRgQaRVPDvINAG5DE7Wy
aXeK1nJJt3T6YOHn1f3q3WcgpYPgB55i5fQIMbc5dEGOUbRGwux72mYOYJKS2D/qdfCdI70sm6mT
Gztsbg4ed9bb+tFSPBNEqIa28O83Mcn8dBoHs9O1H3LQDu3K1AvDozuYYrnltUV9GDKRrx204fp+
qDY2bjMU25XjbEDDwZSX+q4jpNbUwy9OuaVBJ2hMzf9uBguawxcTFjbtu+15AKMPOFJzAUHE6jZO
hYtydwM0vWmqDPfg4nwFA1KBOJgmddJhdBimJscxdkNggXO0mZaxf5KWlgJMj0g2Z/q/DNIQPRo/
9Fcvg5Ouh7br673BxyHZxjb3+IVxKSseBlM2Ne/NSXjFO7oAufvmZHweNG6k2i4VYYLqFhLxt7Zt
X4Mu92LY1GuZu5rZxd72czqjEYan//I034WdMULnuTOr/i5toPy+3m0dW6TirkphV1L9IPy3MS8O
drodDBrxNXJ0mljoTD8TZb5Pi1NmS8GhyTRRjXNklveGD70CVQ01izVmrdfgrYzi8BMGBXoMygAy
qPx7+KrrNx+4326pQijeTDcPRilE4+EznvxMEZhKa+ToBXQAjuoaYUgWi5M8CMtNna9C3KLso1DL
hzQDS8FbHnucJkylGL8b7i4aKjMJQCpPtk0k+y7y0w0Hozb4QWPQ+HTe+78kc8jvIGCnmri7xzcg
JzBZHKqEnfTRZi1Utq6kt7dT7QiiQNS3xzAPcJsLtKXC89RSklQesmvmtjYjmmSJyTSxcEQXhbK9
nIrMgq9/CuivJL9x5ClYqHaz56DhvmHZhnZL0aPDmqtidSLF1P/5JtqWFgXipTCfKRXjHsYohVdo
yTY7e5rgZ2y5z8pn/I6BVtawpauga/OyhaTspEPqCdflHFpK1Xa7CS2/DKyLQFwX4IyXyreVq1sK
22DC1prEn/Dr/2+Vb5Ot7l51LH0+pyW7/FzCECd3JlCz9R4yrNvDeF9uUEGrKqbb7/MDUzVqtDff
F+ytwyn1V3AXRrn5mVesWRHS/uLLLGbOeCC2qnJ1rEmu7wm5K3suPgCr/VidsvENj6ECBDPVK1TL
hHqlUuy2hjPu+7DRu/dn9nhMXX+r4XfM/ROWpqybbYGm1bbl4RvXZVsbbR18lnsWt3MsMDMnSI4I
9ikQA5lSWxgG9oub+SS3nPcsrAAlsL1Dw8Ri0XVq+UOf7gfJFOqQBglDW+PDJ6xgiCifN9KzCub9
7cBJkbuLL7ekkqFcBC9MPiuoKOURiu77ZiQFpCrCPPv15nBbZ+d3Nmzyv3LpZgkel3ycNBTZ6lsD
bebKl7M1WjoL78hYrUyqvO0aUXe+q3UVUaGG7gF7mx+h3lSivjajlT/h5U0yHzW3cX07jIqPCg68
Zig/r7jWJxv5zWmV0sq8i5eSOKrrB+DL94goc0sGsnmg+0dPC/L3HHMvnJfpJX5yZacNB+0XfXqK
QfvP0SqyFS1h1Ep/mkVPUIRw4rd7yRW/oF1O98XoFmZOSZ5YpjQtLpJBF7MsnxueeB4JqoqFx4ij
Ey3WAyZ7X6SBw1y5mOH4wNbIpjkZB+9Z227Pad7czZouSGlMSufk88hKBNal+ax7LPG9KspvPU08
Rg9pWiO2/J7Hk6PfzoMCw64fYJH9gDt/umdKXHmfw5ldmdrYQWhn5eYiSZxp/FoXBCRmLszqWl5q
oNJmTdosnK7hdZKjUVu76WsIINuQP9mWZhQMMNEzuI18Yr33hePdQGRHlIoswllo0E+/J/kBE+cA
9ePWAd2q62vD+WALoDXa/jouYrQPPGBMrUyiXkNivrgvxHDrJeLDiyRshsULElWYRop4/+z5nBo9
RmGI2v4pdiU4EGdMJfncgKqd8hLA6kj2PWgmspzcNRr6xxeDm/rmJxU58CNCYNjtYtzzvNCa2GLV
S/s07LIjXAx7xjhZ6nSOXQQClX6TmDw6HI24OkDgzbvJC9FeNNuH4pXhQX5a+Y4RcZtSHP534Y1Q
9Q3ueiEKHFkKrQKg6G8yt+YlnC+UI0ezaxo8oAtvrlNj4ctGCfuxwK+kcuPyPhgykBJ/AXqlv811
mh9iBTOlyM0O1fRbFk9ZCnMi0i98SU1nK4f0bJ1PUA2Z91hNnUuInsTymH8rVgGT6aJhxYfnLATN
JUn+syn/JP9diN8lrdgJLLWLo/bnmpuSeYqkSAGehQszLsDYUwm1aIz2XyshqvbeBtenkdKgRlGw
JP4cw2h+TrqEWrBmhYEHKOMm51SFabIaIvxqgpRwc2Ymr1fmwlKWY7mzzkM9GUu6XSBQ/BmeKvuy
9qK2FDf2INjH+uDkGG1t35TvWxO13Ow5rHV0A0aFT+cSDiFnS4z9dm2Dg+VB4SmMZWHtSvw8RbLe
tVvrZDpurTDgH9TfsXbGf7GiZG8T0gBn92FXUrSqM+bKevGmLYXn3sJp7MIFVSwYyZQ/kkxR9Yzy
ROEx6zj0Vtvj4wILxCYQwdOsdDVudZ/oMFA6YR/SJ1cGzy5oweTx3F+Gdl9mqGCejdUORYayReOj
f1syD6s5iLFy2u38j0qHV7zavpoKLck2WnwgnrBDhlWE29vKnqOHtlJsJFSTyqt8pWJ8InXuwIPH
Ny9n6pyUTXQph4Z0tHBErLX7B+ydXQuolEcO0suJ91qP5jNtC8IGyn/ArYACN1OYFIB5JtuXfQz/
MZD+JsRpNa8qpOFkbdXyjGBVCw7A9o0Te7dIWKqlZlwloaaEhTNbgbcHFWNKStXJOLoHe5maXglp
I6r0jVIsB19Mv91XrUZCNlCspAjY4BCEA+XNnYsU6JvBMUvcK1E6RcXZgwj1UmK0hK56ipJuE9gH
QRmGPHR+B37G6CdOIRO0cLXDnkV9F0Y35GMQyPuD7p5zM9emLg1YbnufW/0Ico/S3VFp4F3Ca/7K
p+wP9+8Qh2yCixuF2c7cUkWH6TweF0W3M438Yw84isMx+miEGhNZ0qNPPeB3hfFAAMCY1gC05rH5
Gk83nxxYKDBWuCOyUeSRiaW1CMfTFuyxe8o+LIBQJ0d5DnRKYbf6nH9QxNI7ZlIHZVAqZN4O8HbT
uGTtnfZsP26Kui2P9TYL60TGvchoYr5LGr0445pjB7M6Cjig3CHBJp4lveyeWn4rP+aoNdHxNKuF
4xoCnno8zi4Z9V8Db7ZmwE8GVZCN9zfvizcVGS1B+NXkwljY2bTonIpGz/T8G/WtEmQMpkSpKpqN
PnItQGm9DMemPKdfNgQETEjaRHo9zA5BtcYbIMsoGE5roVrxHwnnW4lME8C0BmPpdyAaaayL1N5i
+WG0knHr4ktQ82/KaSY1d/scrmsE8nEcQ42uX9YfT0pWokZ/Y2l1L+jtayMThq8CW2mBY6SZXOsa
Wn1MquOA4Jog77iIYhd/a9PulzJ7AzOR7YLyKxb/UmauGPO0ZkbgPdtcuYHlbOSAepB2+6diAGwx
C9odnhhxkGd3La9dR3IkNHXtQocBfHvEbxEl99Ukn/PuQdD50fvkfevUepygjwqCLkJCrnGPXmDX
JCb1CPaP8CNTeybhomngJiv30+EYu3BeWfIXL57tEgyeZVBUYvo9L6gGSPqXHRUzihhizayJkPaV
eQ5WoRpeoeldphZ9IHx4NRIkWcPFmPwgbBAscpWhEBM4CnBZDJUANFWy4dN2UOKKN6hxXss85BTP
SV/Z+Yh2SpntjgY2l/DgJg5HwbqbpuDJvrLNflIJ33gyEDZJfSP393WTuURs211+Yo1Q1wo2vpqk
6Zd2SBZcjTpd0DH71blSP9q1ngqL8nUNVjGihs9s0kWmkJut7vtG333s6Ktu5vBQBxgSnPJbXp5O
OFYjfVRC04Y/3C8yYim36ia57Mz48U1m2clt3uILYSvKko5QVCNJwUD+hd9og24vLi0QU/uxZMru
MAfcjwdnnzm66Uufo68oASZo8k0LtBlr28inx6VUzc739fpWn/UMWR7K29AnErtO4I4Ar9Kvjppz
TDSxteqZ3xHD/JhNWNOBODNfgfg+nR4G/F1p0jX2BsKAk0KAwIz4GAbhFOLBIcJmQ1wI9aUWO8Cx
hqmp5bMQ7oSzdhQ0+s5KiCMBPOxhTTJm8+NYb6N7KlYvXItUczwhR+26B81IbkDNAU2wNcXAUu+d
jOJ7dejBvC60Z8vraX3QeR1dtc9ipC3YHGr5KUDTBNrXGzuLIVJhVm11qHnsguS08QW+GxXfhPZL
mq6qpzp/Y+INzrYKh3w3j7G77MIOPhx+48x0V/XLZC6zlZmqSq5IZkdAVMa3KjEP4ZqWvFk5SBgr
3EffTpYpAmsYxu8KUr8x+7+lieuF3MEQCpDYm3BevHZzWjBUbXaqiFmaCLEXsWX39bCv43Mqvp9n
k4karDS+4LMQN4pe257MzFleVLo73uykGp+PlUnlIYA2Dn4xyQP5eFJppHUo9na0aqXJyGs5Errm
XpNMWQDdcM0inBjuz+Nntal6LQqvt+G+Uk/LY9hNXfGBuoNTYdH4d/mBXhvo25MwhXS+GRFnTHZL
/Zw4f8OwiH1nO3FvVj031FK/Ox36tQdDNACQUx/UF+yQUab16XrDY0qmpJwKGboIEm3MUpd8ifFa
xmXGlBKzGkD2KvQ0e3Sj5cGlQprhWejtr2PA37Or1oC4OnsHU9pnAawYFmluQJ2xEqniKOlQXaSf
m1v22USRegNfu6EcpNk6xcmKC+UpwBEDOLV6elUnHKrIfpcfpOjsxDcAftNYKJKPccuXw3fq7+dR
3Nd6JO8abFfL/Lr7AaDkl+aEtnWWOYEsTnXJAECvGPGFQO5fcoI2kSOOsAVmNcSesWjR7wcEHvch
DibEXZa/2IKHAy396HJyivO4pHFq3MQf6toMnIJ0SBd6enqxTLJUVGQUV7gxnFMDv3IuqsKUOQsJ
xo+9U0lxB0TmsRX05tICMaZEDO2T0lg1c4aT+WaTNlwCTRZv4J1SFNgAwVmxVrzuudKn9hkKOJ+H
dw0FFe24T3Ds4qDXGgQ88SIG/UVImMbBYryqEJ9vBZb1RA7fYyKYYwYOl0+EC62F013FKz+B6VuS
TGmf+EMYK1kg9K+t03iK60klKExzpufa+D3Hh7TYQky9j7SH6KHhIzHUFyWY+Qx7mPwC5z3w6Krh
+qzsxMo0eySEaXiiyxAF6PZb378SE8lPNatyEKnj0Rj1Eh0oSdfWxt5bUMyl2vXgwrfKEEjMFknY
YsbjBGBa8TnvwT6k4sfdO+pZmDl9qti28Tj2RaYT1c4MAE6LrW5c7F9rXSxL7ujS3wxt4NZPxOnc
TJ5gzm1/JBn+46Zo++6BHBOiTLW6In0AiAY3jDy60arXhheQBz+l/Q8VJ5aRewZ8i4dzVkbCOnOf
oWUm5/MSGrrNUfoYH84eOYzs2bTHe+C8QYb3YQwh78M7iP1xKQx6pojIghMHlR7H05AJwflUN/Ac
WEw18HqfnEbxwSK8jnotdH+CH+aTuoS2jkvLqDu84xT27YXcLuAVrlrx2GRzRKRP6msY+xlIXTgb
0lI4qEWIjEEExSLwvglzeDF0GYo2jEdn1utdDMU+niJL/x0eG+yTBjJGnm7wW51tEWpmL6ZqXwQV
peIb1aGAVd90BYQej+x1z32kmM1ZvWhxIUEuBBjBa8tWjcXdlW0OGpoPq/VFAiwtobS5xQHfWkfG
LBnr3nROkdQZiZGCReXu78ILoCKM6QcjTlY6EZ0uCItsrjlYLo7Dd8c/JgIXgwtgqo2jK2YLtIZe
WvryUZq6QI0Yit80RuIZHdxvC7qH8Ntd5wdFazvR0Emsol/nP+DROa0UxTFX8kTRjsuundevhKRR
ELftS2OIpeWmr1A5oLrk7yYqSlgumuNpAYByhcvFVoV5S5njY1BK88ChBGeZPM0XDDndcDiSpnih
bOWH1qtV9xVPsBW+YCZDaqM35Bx970wAQYKIBpVVrdm/PgvESsmaa/vl5IMrCLqku6mLHXe2I5DB
mPx6YytGRrAebf6KoS1y5Vg3/abketGTg4ojdcZ8ytKzF5PxiXgzz1So448IA6iR5JdBIMiGaUEm
Gr0s4ecsXeCH33W+zJuc6OBEZqcrNFNKqZ1dVLzAt216IeS8F5S4s3SnCRX/SFLINHRmXtKZvjrI
3b/DX/ld1xsuMGHHB2/5W9Q2vdwCCoi0/xcbgYEj5OgdfszOIg8gIWhnrkd0v2b8KGaHie99fc06
dm1P4XpJEqVVj4+A2mVdcdgtF1Vk1g6eXyPeYxBEC6KkS18ILteBFdUUYwJxl3lnUB2K3rYsIDXC
hPYDrgMAvtX3FHzpBs+keKX5+sJRwSorJTeFblfw4VV/Ndnmt7+LKVICTT/4wHEBggC86HKzjfmp
ZJ691eqs0f7TwF1xFJxIWQY/IbbaApwDMPqFYyhwgOCjBvD5GCtkt+gDx49zJv4jxsjsMWN8xcIq
GRYJNLipm56QGR0a85ZoHQ02xo2Y9zgv/GkSzUvEzop6WNupFIbNeHMZKsXV5p2rgvsuA/0mm1lP
fKVXKqbW8P2CqZXhjIYFxWTis5EEbxm3DwainFvKoMydg725qs/Ut9WPf37gJIuW1CuzJjXzSUe9
8DCZRk2rxj8vPf0FH54BTcvPXCEwDwlnXkbVY1OIKEL1pTtqJtAISOeepvrrJhoTm3NkOHSDQ6S9
xgO7RA7+Jw52Q1kDCC2JMkQ+5mTrtWbGFOKriLV8qdHfPANRROABqeUUy0ilLEqKHnWFKDaruPF+
CYWLbgEc2XGZmOSK9Ngd8aUc5C5RkXt4Bpyt+BSFWhEnEQ1zUNl/61w2G0NOUKQlCfgXUZMaFTn0
I2nvB9Jr8l9+DITuE7iUDSuWSASmhg/KgHE7wM4i45cyaerYl6SJ/dhWqIDO0p7aRJ/O+tuOLQkI
FK032wZgX6BgbGP7tdKThKS4YHK7yV7tcXKrW3QqjHC4ItnekkhZH9fk1YfilKcKb1iTwyUsdLTu
d5FkMgmhs99DtyAQrafchQA4e80KDZp2HpHR+wBujV0wuEEweICT3ci+iiR5W8ndhIXwQCon8mQ+
MfCEvUahg3Lfrx0Rv3Ezs8pfKuHCqJua9xBmbXWaPQgNvMnwwiQo+3EDv3VPnRpmH9+bT/M3p6C3
bGvPPKuw9LMSQcODlUyoMNFF+ouBc2DcLyS1lziDgXetu9KqRNCUZntb6a5zKT0J/1SUFuwQK5yE
Zr9BdkH+ijVvSpVE2F82kBUglguhxEUjeTuIl79HNHyGZRUa9Fd4z03Oo9ylWdC3fCPmpJgnBhSu
o03NVXCZunai+znJ0DpEMWysXhMEj5/1BZtofsktb8MXU6KrGL0fk51kaL0BNXkByv+zSXgeABym
YOZTuHBKflTUJwEZnU7tem1lSyhj9+1oSb7S91QQ9JbNxhqW8TyXgOPT5SXGBxi59s8ht/V6zyZc
xuvtQGwkW+iCfpPeZJ7LZs2BxB/YKwKsnOpfsD1Z5Tz8aV83ryo4cBizW2BkpZxVxXmEfvj5oHus
hT2EwXuDSmoWNsWwSlNT2gh6TBmoUEnZw4dOaehgR+fw62VZEslviXu9FxTIzl1igVht0iHggJMr
uni/OfDr3DbNfDhdJoI67HTyv0LMGgOpgVpQ2E/WGr1JnoRl2Y1p8PJGnpbrPmAOB9bbyO9pi+Ef
thdvtyWaDHnB7hHuMu25fO+SIBnQjkI3hSStYV6733Hw9a3bgIAlg9svbSO22xrla0D1DI8Gcocw
/f/66szGSMj+jvniril9YXr0K7Fl9MX2aAEFEOP7doiV9hwEyQdpexwntkqoeTRyRJ7C+m7W08mC
o998xRX0pZ1ZffqVVTN0pN8VZ3GRp1ZI9/i9Ceb9kkP4Pfb0XobFKiucc0U5fnw+yQp5GIo/KIeK
EN/jkvhGMsli+oOgoqUPeVlxsDrUjmZd3eV9MXlJzeACzcXP1koWv0czhZc1ahFMy7bNh9cDSgAm
Dz0H7NXi4ICx9eFXX263/ZPiN7S5SpF9WbWs/gF0kkbLadMnpKode7pRxmi4R+1nFES47SP4NcIC
qmr8rQIQ5WlFwI6cJ0I342+xIcpHe1IWTrR/5Z3SNXdfqv86W9QJvZZvZBv+J7JR+QB7aHkK5U8y
vZ52If1ER+Um55C9r+9fMAkmeBX2l4H0mFYwCnKTRLy1UAMlyc9zqEXF0QP5TB12zmvWYrezfmhG
ZSbFbjkhbyQ2sDjguwUiRFuhn2/uSWF2D08qWSbYU05Bs/AhmQCN4N5gNioj1Op4KpQrX6fM2Z1y
ppgia5FDLi1u79igALDHS5QX7UqRuGI3N2Haefdt6j5yEN4WvGgwILATZwFWH9WyiE97Jn+FEnXO
NLgB48eQs5T8seFN0GvLmFHY7AAPJmOFOnuvclU+Jaxuh/sdMPuF6TiPV5Cscxdk3KsvJuCaosfY
NSp/5pwNany6RfHixP4kwMWIme6rJBUy3huP4A9w09UXAXGr111gnuGoIiTZmeiTIREjguUdSSpJ
kbm3/GO94aIuv/NrKR1PT9NfiNMHeiGOK7rxvliQ+ovX4T/4us1m/TrOB0qoKWwUKJLX8QVP+bgb
vht3YnU1nsgFupYuQO18GLF0cS7+tnyaYqECad23mKKPZ2K9oEI7GoRwn6gICxejhq0oV9nSJlx8
dSa08zB0Dtst6JxAiZ5UyQNgNJyxcDIkZ7Ry/uI+VGrUoAYQPWGG8PrpgI1XzPd/UMFIM2T64bew
a9M6n+87cCHTacVMoE20kz8Q0SlFSagYNsxU5ZMuZidt+STwlvcF9oIPIC1bW87FxCVjCMgiwsrJ
PylNlERrV+iiUSd09eoKZ6eZMoUETI3E7ntzMilDw1nIzH60a1D22u5Lm4YUOG9xriKOhYbVNFjX
GnkW0aG+5pT+2LVmz2X1cGnFIQINorYRhY3DpXexM5AMzYE+UfBo8qhJVchUDFG0ican9yK5F98J
LBUx7lNDdUyFwq0Qf4Bl5YOJrkaBqxiKS+sQZe7vDjPKJuTV8yN8p95fqhu6x7m8A8F+ef9huB6u
B7s+tKAAH1gKnMrrWk/3+H/pestHpe7DpkvxGGSPsZ5trAgyPA0uRvu03VhBd1ithWHeKbei6hzP
aOdz/wAE7hSgRKqVMIofAacrL/Zz9t8ukVzGdgxtWrDP3c7mGroUttH7TULR+oFdnd6sWbTllSMF
6j1IolCaX27eCD8guXa6CV874KGQpQU9r9uBDYm9HxvzfUStiHou1fuozRS/u0xsVBaCJSEw1TTG
dLtV0VT84oUql6qLGqJpj2UOFkVb+0tAPwO2SeINSX01qqI4ez//6o4hRn4h4R6xmKlEQdDZkQQx
LN5ls55RIalYaoqoVpUszm0meTGtSaT4iJayzv/+IKB+mxkk06NO/vXLmpbOvUMu1Mo3xvVX4jYF
0fyBGouKmROQA6fxOiKKlOR6Jx6OshKGElgmVlOYKNGiqZq02/UTHaX+acnGCbGMS0RSVDIzI3vI
Cyc30Rn1+twkjgrQLVUpN/bONagkAOYfKbKksl52ngdxZ1dorPVIbps9nvvPhTY7T5FOvHGmv0PR
/MS0Ei1tQukH96Io1raYD3iYJGoprOvA9Xh0V8XMasiqg33KxyDajcz8eX2eJyKbziQi9RdhrKA/
xb7L8VEjkzEO5U/ZHk54wSUdKTp60UZ07xxQ+ePvXwSoIR4a5D5CosRrrqPbVXNLoFU6WsBlLSl6
rXGfx3wsH7OCzlTP8wzU/p22M2TwNJdoXHAxZ9KKHGiI8252YOvx+Mx1MuIVW/WPs7oadR/9zuyD
wyq1KrzGZXoHFCzczw0E3DmZgtCGgdAVYbMzGv9Ww+EOrfLQkpNjxAcsKKWbiN/ODhAVml2+KHZ5
EqoW1HzeqQtkMpe19/kxQWQzoTxbs1xE7ksTdtWFy5c9NKAHoNxnFHJ7h445uBEWY77aQgkgFnmR
k3RntD/Kw00xHNQvmQ7iwucG5c5YNlF+84yilYvfx0eenGIpdGQvjUmdP06VKs9tGwwjF7zs4sNw
enAkk6Sred6sWQSIDHY7kuDTBO8s+cF/kWC1L2hxi+nPLpFGfgQrJP90aUHGZbKYRKEw4WlhbJDF
Dl+pVdwYrtdoV7tdjJQEmkcuN+pqe0Pazvd+ihxHBxsHQnsQZbA2zkKx16qpTp01N+oYv66U6V30
KACkhYjxY570R2ffmUdV0YtFGwY1JytnhkC/+iXyW6qEpO4huhtRtHqKDLIo4XRgAloNHONFa5zv
7MIFK7LqLEQrAPZTBlb7CRXbST+WHf6vhSOUYtaU8OkffpTA2pQg52XEwNwNYTqrCko31lW5HC+F
Ec8nLl+fp9Iv2Vp1VKAIBtOsuGHMo4KG/EI2HKFXg8gWN4RiKOsEttm78gp2wZ4jH6q35jIEABZ7
x2siOX7j4Va9E6GNVmTrH0l1n1RtDgqw9ca9tld4EUgCZq/9JLRLdYPEuiQVYSUjs5L2zWxnHzd+
dgpVKBV3a2e+lJTWWDgeGK0qwjLDYZQdO2S21j6brlVUpe7CDHtLvmsnofxYE74vHKeXhWl6S7tO
sYTLQm8Dlrh2QLslfF3PgFcFdDGp2hAw/AxRTkcfSQbUtEYa+rhy9WELZyoSYUVyE///eN41r3mC
224zZOg0he8Sg0QECG3Mir/Wr9rFlM7BXoym2pQ7EjF+OXq3giKfnej1WxjRzOVnjvK6YF1VquUG
x0wXOXSRU08KCex/lA9kQUsG3VAFpmNtGq9rVYmfpmWC2GuRaNCupMiv3wWWfUSr84cGwpW/sD4j
xXOG2urXxD8jTFil5kKuYXlLsRgAni0m8WUmn2/4kiWP0pE0rTgEilUziHQweoA/n0BnvOCmqIh2
P/j1hv0JKr0rB3G/SEDzpJGIjYq/NGWBvm8IUJ+RW6Neky1ed1mHiZkbCh7pggOfaSz8Lsu+axEf
tExqeRl+ARxHuqpicpBR7BED0VIgtu/n2LZjFJCqIrGlPMGOsvOzdD7+NkH6rjs2pWSRXu4ihsNz
uib1ah5MTSFCQjF2kbUoPJdQUDgXOfp2+1YGgqkeRyXTjQ2zkZTbfJSXNWlV+ZzNjokpsxHEBklh
QZJXeDwgGl6N1cBE5JRDapMzZ1uswBvYmmwgtYUZ0NJPvnTW8PyBANDLDEWZ5bzR082u2IFQdDkz
H9MfDERVubT2gKu5uUGi3GSRCQBQ1tfdnTuJ6AIwJskMxUKVVovfNYFsca6FFlwvvj5dAzg198uJ
LJCUcLdJ2GE0ooV0Xf1Sb3mlR7UtkLl2GZRr8AiLKPo+nJMQxqjzcRhnnE+FiBsYDC+p8mNx+ZWO
eHLY7ZY7h1Dj+8xvz05wrWCp5ZFT9gYeCK4K02qLat6olfluH5LVZvqTRIkwwuNxQ49gBJew0JgU
9Wxr5NSJ8LGV6WxdgcGV3yymf/Ny+snlBPy4CMG0TCAoI/scFrwS/st0GO/w/BAJ2ojJjkvWDMw6
/6gULAH4B8MpSVlHtWT1TKV+38GvJFpXrL+YBTj70PH4KMD6kByucRbSER/q/GROPsfRF0wO04e2
3txsDDRwqR5Wj9LKBHd1DwS5MrZeitIXVYH8pijJ9ltV3dEq5FooxJ+m353H0zYUqv9Gvdu86R1L
SRieR3O8TfM9EL3SdGigOUzmya8J+deKY+27K3dBvkLRFrOQ4kpFrlh0+cIUG2ggw3KDvKfXzXDJ
fJa3cs3uqUquad1zeJazB0TT3cCusfvwdMSJgcZGwMcQ0kNNXK9OX0m1R/fSK1lKtn+eCeU6ABNn
15JGDNjDiybr82bQFhkJzQkY3kK4xc6AGdb6ey34vVRh4tPR4f7KqeUbHunAAN2qGRknzqu65fj1
vhvlqaQJgJX9jbhAOu9DNsdbkMsYa4Q0LrikQnRr/GCDcoiy9ud0nIAUL67RKUerqLx5TcSRXgX+
mW6lrqe6Vhq+NnZddaBLhxT70uX/QsmscyaRzeEL1dxqqiJxIj/eqawViYBOldLiMKBCliJnE5SG
spKOSJJP+fNJnyxQFugk5cehXf0m/NOhk+x5na4i76YWx3cBYbJoKDkrF+TYe8pTuWwrX/p+aGHq
7ok2bdvFNsqY44q8UJ4oFsNIrhfFDPbQ7ed0bUhhO25xn57o+/lGOyW59DJ6Tvd4zgFOhVAt9Znp
MsL384i2YdTEcP/Z2YlNOaySypwqSxOsvVT2MMS1DndpLWkvTUUEU47dAbuHxmnvI2wn81zCz8vu
OiCQJf4ObfC8anM04JFNDDWAeJzqqr2Qjsr7gnanuD0gZBb7qBagMJpuBwuV9603eUOOGgkml+Qa
ywuPuEZcOVZHYaJ2Pd7O7IWMPJ6xNRICAtv7IXibAkNH3T/U0wfZaGFCLYt1akHsb32cS1NgL1bg
TXR1ARbKDmof3U2O0PFwUWi4VhVKBdNKAQBjVEqGOjsPhiOAaxPCM/EubnBmKkeXekE+TvQf2pgC
S1UAGQzLiXgzOAMHjM3djf+dsyraCjQai2Xq1l4KuGr2igch4WxZAKiEU7tEt4iiSxjL/Fd4rVkW
Fwwcy0LX5lebduCvw2aXHXnUYQhOZILwSNDMihQ/idWa2GFELTaJ+jQQH6ij/JQRjCpLk7Ncrlk5
vPaGLvgGe1vY9Or0x4/A9Cpdya6LlJrGmk9yalo4NLkQgCSrkv76kUmkv+Y96vO9jo9lmYHsSRrW
VAYw1JHp8zTZkmVXyI9FAo7HqhMT60iy1uTLnXcBidbljZMPOoj+B9nT9Ob6cQCahKDUOmgyfIhB
KzgVo/gq8Nk3gnhrSaJiD7D8ApK9ax0UPk8ULJHp6lExcDToe7XLbSxFshTiwHP8xg2ALCKA5y0x
MKKFmta8chOUOsc82elBxw9dYfXTHAILV0GBaDFGP9W7oKLlY3VmhuoD//u8IQECglWqUofKXEvo
bkZo9oGXvDogqvnTuJMIGey0ISqEClT0XHb4yZue6nnoNIVPmf1DsRDtvr8XYMdC/ENyFY7txWf3
QlaBysmGpAzitVhoTIdML+OeXE6ULZPNOUxTbbrTvygJ/+SptuxExZZVsXIYvFsgiI5NBmYhoc9/
um7ObH9qyEAMnOHXROW3c/lTqu9f2MZacwPdZoLoeRBTvQClcQmB5KN/oCat07Ev85csVTutwnl7
aZmT/TWqAhNzLwVMMkwMHW4gRUAN05agj4dFCwZB7FZJg4G6SaNxNvH6MiG/+zVAE5XuHRSiOZ4e
CpbX/PWUf7dCatf7pQw95j0mzluf0LBvQYsYCjcm7TVyPV03PzsG5fyjt/QBEbyPBSmqliXSafMn
vI6tKuFPkGzp3lOxi8is9VIKCM7H5fbJNRRDvPamYz7xyIsjhXHyK9Yc8jSq8B+khRQ4XlFCyB9W
kZIJ8fC1PDAGp71BecxP4OaYTysbHnnileMOtl/B4g9fCf5ggKOzmc6TSqVaLJcBflJyJVUaZt6T
ma8xUValXEaBvziKRazSyJiLnL1WROBAUSkCXutRQ7VXGlEQ6eVxXNe74E12o6tX8GppoHpxgU9s
O1qClAw9PcBUMM/R7SuaCyYGfHSfMnUT6X4SMPc6o+7osKIHrJ23jZESjpjYyU8TMGuiQW2jyk4P
NzcXvk4wuXX1Z9LLrgAnWdpJR9Mapuh64FRkFq10x+lsaKIjG97C6t5l/voVuvj8xb4FE70Fugqh
/2+ivt10xeGV++Q6Z+Y3lzVtMwRG9OAfJJ7wCKpx45WKxBy3ZZRMqTsz5Aq/V5kII2QkaTAtfIgV
7iAEzCnu00ht1AQbt0mFvam2jP0pkPfGRAPoRMNvJT3CWLNSVvXEZEh7B+QaQ2Z+6ZmIFvrRq2tQ
GBM4LjJ+gIwx/OiKp4H41oNfFGuf+K/J4yARYDYeYH/JQwyytKOTPDc3Ru2SgfE4DFP4RpuA9meD
UVS4Bo1kMk1aHY4Ugt9gHPq/LwJzZWZQ7xDelvHFh16dDdDB7PeAAtu47WY2IGpWpTpgRi2m12l1
FrDdqEfmNspcDtqBSCtxC/OmhV3kFk3mCbseEpcc9YeCNRd7OKdZBXmecpkhPMOWlyh8hJklQBK5
puruAvnriokjkzJho+dQLsVDWFxx6h33XRLxqI97gi7e2Zmz7FVQtiV6oZt12/MA5umVfOBLJUBH
JDs0aLlFT+7gwJndJrqgBnuI4d+CM08sja6u1y0IXK6tS/+EZcphGf9glWApNh3GFaaXu2u2IHnU
X/yRZVaoGY9+Y3n5X8NFXcn7kEWLsGtu5m3YJ8uvLVf1nUOBS8smIqBXrX1SmS5XcLv03RI5+avq
QG32LeoayJzpfWRmV10eUjj/Kz2vaUrTPKD5qno0gHCIDtIhZigMX9OIbzQ2ZOZIZrUoxa4DWRF8
ANHwLGVH8HDkWWOkW6h6hdGDgZWoVbnHrpx3piO4/45sHz+DXqsIiy9pIEQn44uCEhkBoykDXxQn
EccU+b7IC8aMNyCknMutB1i18dmSk0agxvcJMAeY1d1FDCcxsdW+/a9zeT0tga7ID9VPV+nFIZTa
KM0i2Xd7DmNyCtC3OqFTnpCLICJzg0ESaKovYzX9b3AU0Fy91ajArYX8+HZK+10HAzBKXpdkQ5HB
GyzlzrmPyDu5H6rwerh/RuLGUXaRUU2EeV6mWageYicrAJZk5MS4K5qS3+VFn7OFg52H2aRaNnoi
PeRTnmdmSXmIopx1/5fyAFL8QPQs3BC1WfB9FvcIUz2xMe8pR4HRizObgjrOlzYFTG/a5TxJndvm
CSuQHwTp78mbAlXFj0epPZX4Zf7RdfC2G7TY2SbaaGM6pdo1ycDo6XsdrXj+FvROB8fhV+5Uw6pN
k/jc+hCEOOkxg+p7sq0rbxqQCgHtrI0ite6AdKGS5+g3lr8yWDxDYYuQd8At+jLzE35pK5i+sEgS
bd7MGZlHSyBX3qLWRUHPHc+q0H64h3LA2P03EsIeQcEgHjX4XENQjHTcceqKAMSUGz9PWqayH5CI
UwGnCTWD1/XKmIWso6OA518ddTWH4bREkOJOQPHv85aZX410Xa0BDMzx3qCwJ512OT62VWMcQWob
M6cfQmejdC0Ki5g7IkwUCr2PPVU6hQ9MrYhFJQm8Lgsvfft2XBkNv/Sz6mTuCsdb9srtCDP0+hf8
JmNMDwEFI0sTmHVFJS51J9HYr0LVLv7nhp67M9g+m7kiN0cjBEJj5dhNav8h8Pd3rNjgPOCh9d5C
DXLD1/VlYBluyTgttXWyDo5zCZ2a4eIJPQb4N7WXr5m1IvCM4vmzGQpPdKOPyRqG9a62teoIj5g8
NBIiwCld5Ms6Fj50iTJ8DHZaAcfnVhqmMl98gOcbwgo0PMGn+VOhj7Cb8T+dIfONCCCaL15XLrq1
50+0hKb+YvVi0dJCcpWgwUbyOM1Hvuy0LvjctBD2AxW0ST/RhiOxjl8BI2gxlkhYU3y0EPZ1/OBn
Hz0+n3NcGIkoSEKyN5ZzJe6aQsRsrX7Tms2qzAilOnZerzNGzf6MwNfsE7MHqxJsFkKuOnspSd+3
oOiaGGzgE/41GJyM4V9qLkNu+atq6f9n4VELS4I4VdCyodtBtoyxDSUyCgMriANXAJmc7qDdUZj4
EATpLwNlsq3wceQZMt1y6jAjLVS/XTBTNao+VIQ3ktSxQNmfOrVXgGiTc3R+CdJk43F0TMBxALPW
+b/CC3+OcNnMpAA0VEsKTC2HpJShwKBrIHEz8DzC1BNpPTDsFD62QOQMvDhv36FcHDgcAj0zOvQh
YHubZLDV4pufqt9QbxTLVuLi87Seh17TpPrVG8hImG6BSQ8EgqNshAy+fgEOPAjKvFii+0bM0uUR
mY2lvBGqTSnTQkcD6/TQecFYOw6/FQS92gS4agz9tZ4Tk0aODx1vA8V4M62HeyX4Qz8QtCZesTUu
ESEAyafGMIVLdHehoKewXwRw34tp1K68LOmsZlKlTqwpftqkQZXkthmqX/2MiycNJdQbQm5Jd+LY
t6yWbHL4g979/62jyVaVbme0Moktx26bDjlJPKbLBzHDOT7EvqdpjplL0A0yuEJXXwNuQoKiMlTS
6LHRgL2YrWASzA+o0Qx/sYXU8mWYxb43T9JeEZU63sPbKeCsnLDtgCtidxcseNOnS2eyvG3sn794
Q1kCq48UiqMmtIal71FgfnDZulJI1xpf9dxtTfJVKfTRavNa2qelikYcm5l1pKSUf5mLYtiJ4T7p
W5mrV5WNF6x4FByv5NfngoxuKn0dSzIgdrIXobdyFPyLNUe1EZOLdCR1/V6IDNQmfH7EDR/jxMT4
z+Ph+1pBcfxqG/M0VMeIo+ioPQkBd2BhQjieXaPJubmPYsLd42uF9NoHOJQ1u6YX34jE/5LTh7fL
K21GTQ8yrprxCulr/eRufvSA8G5msOZ1VJmSQOEFFHekw7fyBC/XUlLluw6z39+SjnN357G5N2Xk
gn2Jynlxb0MSNqGHKABf6JUqBjuQjkRV5d5n4vgBEuuuEKuKf+JFkdDZsU2ej43FmjN1MAoSMCAj
DalAtDI5axj6v51MNv3zmk19PlsxDP2HvUJjFYvPSul2edrQ5HElQZO/6mZdMjjgL7MUjmh3d38k
5BQux818xB+qfYMBwZW/IjlztJ4ywKXzEg/GINaPaMGtpcdMqR645v3jtcHjqdaqtGxBhlo+gUtu
/VEzGFWppBlYgQNG/sOebQu+gbdLcc+2T1uLK+mcZ7R0GUgWP2WE6s6TGHR031CcWl+gw78X+rg3
woQK7IyLhIbv9UF6OdSpQzj2/y0/zEPZQLRysnveA1+Acpc5pQjLZ9r+BsLithWgXTvazJzBflcv
1v74cGff02Wmy+Bvg5XGPrwFUrzyLwocf1xWtm0ScWPEqMjSodfhX7lC/0RBnAQqlt4fqJNpbRSm
g94F9grT9bWFo6SRuHSOgvelbga7AQX9Hn1QpbGA0jk4JmZl6uisStBhDMGSww5REzcQ1mWVIHUy
2JMPC7lbDfOQKwrBLvVFsnGhcPkR/V1qelrAt2E0rYOG6meUyWAOuRdcdhj98hsejPHF5KuB7mL0
yg8CrngTP9a1a+lAwsUVW1HB9fqUwK2yr3ovpuXzyljNULFQ+ChDay3knfYhhYnWmZQv2QW/RX7t
qJhZNACsn1yMpbw3+sH/VIBGw7Nu6ChrAyTZ57S8aGOljsXxGhkNzA3IzfatZvr87oWVarAD3ixD
zd2kvQ0VO1Ox+EaI67XJMrp31xL3cFJcgIlv6+h/x9nMyuzumZ6Ci8ts4GCx1glI2EoJQAze83Xe
Yafy9vjcru3rMziB8XSB/tqDceeNkgvRGUHxjIZiZSR19gwdcy6EPfwSjSRlKN/gFBk8l0VkaoZg
ThWgaOWzRlVG+s/1wIIj8DCVb65TnRFYpRBe6P+Rkb5nKEVySLz8I8+94YHMjpLWjfv3PsDEXJLn
teY4oiSqgkL5SGfel9wQYyMglPPE4MOMr1b0H20gCoN6WgSP2tsznR4bwRxHseSpfq5YPnTskYm0
RdkzgOrB0Tujw0UoxYY1YN3zXnmzhkCmEKfbFPf3FCILL22Kid4moXjklR/o6RKCwsBTYX8A06eK
ozMjU8QVN6X3NJVb5IL1TYfLu0STgfhib9P1JZayGIsJGIqROktszTzIZ7z4ZOyrSNSKZTwsGlwO
CR4567QOwK3uRRB3AYSzq+gLLy7z0r+p4XtCM4NpkF1tOblrN6YzpX4tMfm8GN5QUqwDOX1fxnIL
+5r/1qazZopJce6bFh2V7quNwgWkSsekzYkoNMyOWuJpspI0E3W5av1n/Flk/bWKTliZAF4eolFD
kqh1a/xRc6aeaZ2zQ912laa45TgEYPGXdKVSHN/E/pvTIzHQ559cM6otVtYl5IeWizxzNPkfVQIl
/ZGvgfay6mbIT87Aq6SPuCncDJRjp0vBUsJot1QfcAqYw8YeEyo+XB0nooQ8LHVldavxTICpGt5r
YHnLQezACcrySWNNk5AmptbxGJUQqvccLUjcQQ7mn8OqVUa/mW3b9o3oL6xcGbXcqlPvlR/GoLhW
EQZPBdHg8PsYKi9kxZoxsUCxnJOqmKZcpQOrqweQvYU3Ps4U2jvLWpiBsi5jVCOmKUpSUFJ7xfh0
KmQP3mQl7pzJatILiFKaFTMpTT9rjDEPFkNVrNhdA3rHIuBzDQawEWRrDM1VYtASsadPuD8AwPn/
5Se5xtJpP4QGouOB3QL3Se5OGch0iryKtZSdLmJNIWKfPGh9TbJyqj3RjFkDVCIhCS7cD1I5i2aT
VJXUJ0ckmds56CXUMpYSniXmQAYtECjagvr6QFidgfciFkFDjjjoJwF85FRB1NobfiqjOeJIdrg2
RaiVnnleGqloA396tu3wQkAssrqeISM9lnlbDbukFlIOcVXUFRdu6r3WQa14oZ10+gev9I3z+kpu
swEVF0cWmXf2LllmwvlvR3xohgHSsEaSVRExhECkt7N+9deoGiHIFLZKM6RMemRgjOPerf2REYMg
rEhAy58d1DOH3GahxGcHck7VnkJdiWEak9eQ85yrfaJvQIOI8cmOw+08xr/7Pq1JCGlqXFmR+iPg
RwwuJEHPUM/Z3vU70JxxVx4AH7eu1kx+7SQuMpSoKMLXzkIImIty+57AWTveNHJCBS4vyFMDbEFw
S45Q/zxIiod2S9P2cKBdFwogL2iCoV4CzXghBwPMMqnMw5eNlfvARh8dfq9/aatJN4iGc7XlOI2a
Fs1EP5gXttyzQaTECrW62KHxGHqL+Pr6DxiZBTPqzGHCxZ0GVeR7/XRvgVaj7IrnWwmfDvcP2XQl
zGBWqQphrVqfqdQwyjjbo1SSKmN4EAER2XbBg/Lf4a8BRjlUA1kWK+sY6W2oL2qN/ZWXYmJxs9Uc
n6b+ERkkv+t4PtWd2wJ10AePzlqemm7I6xHObNj6fwejpHa0MsHdp4Iz4wCXlzw5QrNjKR/bSubV
LoF/JwSTlsE/t8fJKpdxAYA/MgICjtuK/IoWhBfaiT7lLpXPSRohTT35+tjncnqK1yumQaXityej
4XrlXd6QKx9kCH5yoXN7YgB6a+O0MBksqkyB4FRISfeWHm+hiDNPJ0B8dRKWUUNdsOTlAzCR/LuV
5v+cn6aHmmutJr9nHUIqU5nzHsm30nlpUnLdyv9ZlfF7Lw97HbtiDzGr+J25VotmgA0tRFX726AJ
SJonGy7jLqyS/2cbJDrQMVWFQf09WA43z5QHog8HJZ4rVT8Q7wf/r5kqoGrtEOPL3s9R7euZkc6E
mklS+SQyar6pJiTuxbvwVYKVRTS0DJc6Mt7QDvv/ToVtGwyWSd99EvcHUsoJ7hGVCZxf5QQd6+HK
MT0mF3w2UzivEusD9KtwzoqZFxPRUJgEDdlbrKxDEA+5OCSeaCurqkbqd0Q+QIoDmWnxvuYgcU9E
KuqYIqHCHYSNOdEy50CGz5f4kAVUZD/NkOBIXmytFGWXvZ55y0Ub7+XX0Bd4TbAsaKXV55uaOYkl
JdI4ZO5Xa9RXHZda87fB2QmuaNyiclmW/UYhmmBaBmIJSOIo/hFEcETJb5jCP6Y/FV+bjqjXxfGK
JyPsPpjWgDcuTEKT9vYsyDrx42jNpBLU5J9jFZb0H7lGg6moNXcWPtWkVZKLoShBSmaVcsVyNqCY
UhbY76hghKkGXpb2umOEnJegtI0Tw01VnGEC8CS1Kdwv5FO09kzdliceAbjV3T4EopyZAOSYzr30
Qfpf0UVpKddQFEvOZGrQzfn/L124lPWWudxt9Z+lAY+UTWZm6Hw57xC7B/ssfmW9xxoKrQLa0JAK
jJ/8/HcAIJXlzhRFqDXd432KWJFPO7no2RCVrMCrNGTYXk2dY1hvD1opCJU99PqpdnseUmTIHX81
eVbPclEH1u+xuVVXkrexPianSNxJvAI+7ve39u83GTvLMT1BJZ7C0kOoy23PYWVXtroPsve0Xc7c
n6/PWb+SFuF6lt1Z6yd11uuk+2v4JVpVuodyLfTSJssc53PNXJ0cSbZYTP5lnb6hOw+ZKdbXIEKr
nc0CVvvYfBtb28Uwqa9Eh9/IIxuPfM+8N8Rtmkon6MT4fHwmPBY5MoGYMWG67MZaR+zGh8Aiq5d1
jJ+fZV7/p0HkH4aTQ/hp9oQsIO0XVphC/W3nDoM4HI31rE/6kuyCQNGs1QP3vlW+y6hnbQ9177Dx
jJciPy54SZcvQBHVwr+a7sdyg5MBuXdZCuPShiOCa/6N6F4PbmJIgc6+3LmuoyIOaLvZJIkNSzmk
dJxb/70GS5mEti/sF5deOFveXLWsvO0FOrQnuiVoVA91iZZpoaHW3wzWSc+ASyjQ7/eurVMbkZJJ
NXZetgoIkiFooC5w0S86OJ3zkaOLbEp/4ZsDDjnRh5I6eBrF/P71+4HiIVTvvkgWWJt/5/ipER8L
q2aAmz2fW14W9OGWF/1FNDMZtCM8Ct6+YyvV2KICIODH+rNnWpKRchClJg536hev2JPGtKY4MAKd
3BGlBQfgixRfuIBDEn5/9RYojBJhQgwR0zLRI472nQV1ivzEh0t5JFLAf44KzsOaSnS7QF8iWGh9
p0y8i9x8d4/tTWVQ7Or25G1/UkskoV7ZNu0Byun7cMfwR0buoQDwgddp9ar2xCXp5m84bsFPCjCD
oiUYS4DemKODph075Dont5Z+954QfvBkZHPtlQHd8iBiao74TeixsOmCVKu5ZDpGFoU/Bb94q+Sw
crfH1MJhH+or19W6BQqzrM95hInbkxzNZTXhH59yIkQ+8Ac0QS8VNxtjTamKAuxi5g/OnxujtcK+
m1MfZoGMXghvmJmQPzfNJR6tpRHG2PNnOTiiH0dJKJXULTaYW6GI9d3jyCYRsG3iQQtvk8mOppJQ
7HC6m3zcE7Fz6Xc2gEq02ImsGCOq2Bkrjf9TZTKoR8/9a1jnGHvuAi8HtJUGLkjA6vqQq9b6e7y9
j2MR0vipEJQBh9nv8bgqry7+gxBCxCHFYGZxyUu0NvquWOQN5NGoAG7Ym/OEPJ0G8kd67lJ7YdR8
yQL7QHYZrHhuUvuqWPLtfIgOcEmFtir20M+1rkyX+3XRxI+h5pITlIJAEyEW4qTvoOb7+iB7UR9c
cgTt1j6vhKOXxlM46ExF4ReWfJNQeDS7IMUabkFzJqeOFJURKPwDdw1+5t5t59n7SRYTQgI9SyN0
+Zb4UC7vNaFRMxiJy+uSkz9RChc4Apr5JFjYw8C7/KbFu/YZtwh4P4ufph7l44lSb7zLaPPWLSL0
gIuw/IvZdGaYdnl/2iLp1PX0LANr/77+iUPRNS6uN0MASPb6k4G5/KHRVvjTSnKrcnWsaJ5w6BUw
ikr2okzvVc7gbvgqm9FMpSdWWZ2QvMK3nHT56CpCEzeFTqSgOaCS9xjxHD53lfZJ/X+qS6z0xGel
+vs1rYZY/KUtpIzugz3UnMdMnT6wT7ttXAQtBd3dgt3G7ltQjVORsweOnE/tB7kzFtPFce58KrMq
+U4gjFkH96Yiv0iNjsMqiXDcdstvuvXmNrfW1HYhoG2oBq0A29jVV+SJgY2GFJW4uuQS8vQuyzBG
cbKZTvfphQUpk85Xftb/hD27T6hIrXcPyUSrWli7pPw68IN9kkEM7VjjCXS+dSr86OhSsxXbT6M7
H4AcBB8yQXgs1WdfudAwq2B1B/ETncavqDDNd24cRHF659vScIxS8Lq0JZXwyaAYczJl7O6ODx7x
f2W0VgjOUaAU1wyxmxBho/zuhUFexQh5CgFDxNVn/AJn/fQ0aEts7wB2kbEfgqxaLfcQDSIbniRZ
6IUYciQVJbZGQjnPPoPEiS0iOZ1Sb87rLuQUYI4KPRtA76vmNnt4eVfUQdsnmsSnvS8sWfpZygW+
cHG1HvBL6r4ZztPGKLFeQ5ZmKP3nhvHl4hH95LjjC8+RlagH4ppd+ZP2dK95zWY/SSbCnfcD0DXB
ONfkUwk9VqTxI9WXUOcPMBzTYax/6eaDy4KhxJGGSkKzejY25c1A99jDS5a4y8eSZaUiXGnfdahG
hZb8UufSE80k8cSI7l3D4QLi5mReG0ElqcRhRaLEZIoyLCWyUBHP2OWz1mOyQmgmX0MXnQi87D82
E8FIdi81guARGVTlBS4vmD9BzyILQ8CQYlil80eJs5sPLVnLQy9SOhbF7nqZ/+3GNugFhSfbVJx7
Rc+s+oEQqX9W2P6YEu7b3bcgVaw6O3Bc/8KpUIMMyqnkrb1hKSe0BflD58zuGWHVekgQiBfv4q9+
kAo3KQqY3nrQzPx0zFFmv7+ZySTrFhQFq59X6BXN6Q1d3xYEdMBRsDEeiv7ytuRRdipLD0y64kNw
GT2DgTKgEtB1ZCVDQICw1on3vOKrPqw0yUS4yjD+2O+EQ/Nb/t+NIz5Awzq+3WFYlYxrxphXWYoB
8GGj95p5Thbj01MlYF91t0Y2YfrHSMf/6XwQ+OscoUUN6TpugSi3/mF4uwNSjMuB13nW4EHQXqQL
gxdgZCU6xyW+hl7Frk9JtTu7/IpmUdRFtOsQrv4r4gbZsfL4kJUs4g+VDtwuZ0btRraJZ6/77R6I
OHx/SvxB5c3BdfFIHLkEsEobyzQqopEnv12szRslIaHaVxI/jTKhZx4FLnDjPdLxJGurjK/KzVKU
L2i3AtC0Cu6wgvFQFouKadCvzHGbGLnhHj8hYsnc+rgyhAbDzlDWkg6aOYenZ2uLYfkA0FEOouHe
9+5B9/DFTV0uqY8EYUPgEjTQjk4ovOhFDX3z1rxjmTkeuG5jXNseB2YPu3/2z9C3Ja5r+zDqdK7k
Sj33WYNFZl1nI9kO7GdR+bLT7T3m5IlzCCwOdO25YpREcCTRsD8Y8JIvqkXLm4Cpy2vg62TwNp29
rGnBLgxiLORefRgOm5Y6OgbnoN5LgymD6c+A5JsAVhtMaBDAPiX8JGu5sOg+psVN50h8OoBUUh/c
NK1/K8LgOwD6Z17dYjXIP5lU/vDQd8B1Hyw337KtJQ32gvWn+Pj3t9+UcHcJywIebvooaLWMfJzi
31acJ15FXtG9hZ/WNl3T2u+8V3zocDtyyQWuzKpfMbWqd52z2HtpVLQoGLV3utjECtP466ot9gor
LyAFD3UHy+d71SSAZGGwGikVHZ9LfzoAzFvh/JKvyV14xj9W6g7y0daoD39NauGWnfw5cM0iV8y6
8+wEoFCG561L7tCBuVocOVD+pq4nt87lUOCXGHe/va7TqLLZjGCOPsDWn4uzr/sJ9/bov8HzAm8z
kjuiw+inwbk9CT66Im89TG33Yvuq13x67jAv46HyCuzwrrApiR9EP8gpmy3vdWkUFDb+OB33wJq+
YdikyuBsHmBd/7ZX0rQfFR13WIQGHSMBQ8onSfO6rG4eHjHLzJ+9jTQD+dJPL2CGb4ZYFpKUncOv
/cEvuOsE1L3Q+qsbV0CScMMIyb0FcXadtmZOtbGh5xqXboufDK8nGytRPSn6e/QoP9py/Y+G9mfJ
68OAQw4IDkBEsS5QbWa2oj5V/GefX5KFGDIifhiGT1+ZlyzP/DrjGFIqmdHOgVbcIDP+/7bnoo0z
WlEDD29PCOay1/kgf3cIbQv9GmKCzZiUizzyuhgZewFOVyKfNyaE3BPsuX9zLCOLNoYe21drDPHV
UBE0HiOI4PhLNjv9bHnNQpgu5/vn3HjWeGFOY5xWOvtsiOY6ILCMljUC/ML6ye4cTTmbsoW2JxI8
hPpq5Zfu+xn+q982bxOMNTBW30QgDyZ3VLpLJ2YhlrlHHKyTUPeJofldFBJ/tzA+bL6h9mqzA/YG
96DNDBSKHE6tDa653IWpv4wAcB4EU5MdeGezczIIudejzTWUYOEwHxATBjlLDseb56pgQwU41uXk
w/qrN/3HeKUqUuWXlDzPY3tmRyrHCpkFIOzmMA73CSxAVBmYZO0QEPM2E0kSpxPUci4+s9iulfeS
29riDfGRLP9XVoVi0gkRt/NJV4nav1SHGyygZEh8tu0AfLalOBVvM/RRSQkYJqVwVulsUlXFMEQE
9LeJYfAaKfIGVExEjZrRPzxJHi9Fo/Vue8KRh5wly3r0aT2jEmEKVfL8RZDlO+UTZ0nxSA+GG/gA
Mb3ziYQvAsjZPR2bygSRcFSIV58rl6yRnMnYofPvJRqu/+W4GHH7b3gha7pg+KBtUOq/SnvCMmN2
pCfdz0TUeCAZPSPfsoNtauaI9LLfixt758cRX+bVC6H022uZ4b+OgZzl0laz/DyMnfeKIwdKzRIN
q9T/y0lvxnpFxncWGcn/8ZtPvyG4RVsM90OrUC8JpRMomnDGWkXosePOU524L8qKYZsUPu7lSnzA
29jNZKSQ8qWTs2QlNDCuozrEP3uCe02WZlbTKYoEj/f482Fe8qQ+IuFLIQepd28nWPlkcHByacP4
0mcnHGdhdgkVc9NfgKwweeTNiJ5dWx7LwOwv4GAEiHDuBu+xJFCGV9Vdivt1qtOCaKxAUBY/uZWn
p6HvIt3P+PxkMegr/AJWhdihJbg8Tli5I3wkZZtIUr5KdUelRu9jym8Xr/ABGJBkQKIOuojarZIn
HwTT+rB+yOoMdUbGaFMTNIZwZSOwDdDp6bNPNh325c4dp11W8qur8leZo83zWh88ar8kpC7yrp+o
hxkxXDPXOdiNKC/vN6BKNQ7wV6gyy8ZAMWSePOLF94Y/+tSJHy0YWyiTCW6ufKP3nWAAq2Lb3u7o
dp3jSfkwWcTR5RB0zyLRqoQP/3waUw4fg/rYLDhCt9b6JyJWVkWTtNVJFjd9tBxwNMFNsg6jT3po
fwMirZyvrxYqJoiKIr1YiPuAK27vZZf/Uu1TkYPv54+gULluS8o54D1RD37VriX/SUZ2G2oeo3mV
0U7ZVmpZdu+8YppPF0QkCNFD+hFM6ciGrzPydL3di69DoTbGwn8umhNWWT9NkVMHT6HdzgPXT9Hd
xG9nPOpVaQCle1lC3wrjU2ouHmzw/yRnazeTbU0IOQ/lRE8CidsBjw2PxPn5mYe5PLeyQNFyJ5P8
MfQeK9qtNpY7SBuY1A6pv57F4CRzL7vX3e1SGrFBTPLyHrRsFqMUEi7YcV6dmntcpM4gPDscddZd
CoxdXL4u15FumU/oi1EVi11847QxB4J6hgiw1lYz5+BN3pvlOa+FAGluSfYwqxNgTyFbY2AzFYWN
4MEclWwBbEW1jehO6YQ9xMQHHpxUomg/ONIxNb33ElxjW+sFjA0/dlPK1Vn9hVcPVFSL59YAXdnU
8qgVb+PsNjkomdobPuRMi0A48bjlnxV0lgReiyYl4PndyzSH4D6dJub6x2WO1l6Hnyx/Kui/eJjz
IZVkZRdwEHo/MhdysSBC4Ag5Du8R9cAVnEYSgnb/L4XJxGnnoOIRvTQo+K4mhg/aCDyRqjei/whx
xHQ48xYmJLKdqKivGw289KLkgtcl/It1SKfQN6iPIR6b+y9O262AUQXK5X8vrllVy4sI6W3YezNW
YZ5DD4l7FZ0bQ40T/OXVQ9r2rV3ZTp3lCXaOeIXU6wnQKtqwYuUhlJhiHxZ5Evq+uKHZrY/DYysr
Rw8zHbsip3HSmXK7V71IpXLqSk+7bDuSyufrANsamrTtsCrRHUm7edS3RdQJoHfilxpccByS+Wxb
p0xMOsWOdMMRQXQXTnPJLZ03+NMjA+oyFQyhy3Lue3R8YWU7KegY6LvV27FtpaFfovAGJa8puqZB
yL+pP0PG55HUgGI1XC3OCcpdPgW0JbIeQkKwiAQeaGJz+uphSp70S8p79QsCENxHYZ5c4yDIPdJ2
UKm/5BPds1Xvs9uUDsGidYSORAvzROUwokLwvRaxgKnONWeEtKD6cWaPftqs+PFIdOgw1lXuGyfP
zoq/LhlaklSvPut2bC+rHdSOazRUpf4ACGjsKbyMuzHw6/SPGqTKmAuV4qFBUjOBJybIIU9pCSrs
kBjypmWY0YhFm/lOR7dvBkKQY3H8x6S588pNSMb6Dc24BRzN5C4OrWjDetNOdiahpIW4hzXDlqku
Dh+TM9jwl+99nTlH2g7TfspICRIuk1NgSENjDXxTQMgmgj5bdTVlAvX3+6LE00z9GtBgVhQfbpFD
Zj04D3AOejXrhtEwd5yCS+zbHIv5iLowwVKUHD3SfP/atYKjmRVuzONOwGmJCjt4gUVgPGch7Veu
20/0jy93n9n0fNSEcSOsMMx4PGo+nbr/dFpa26G90gL77FoY7pnBpvtzUnBu2JHePglSg5Q+aN7i
kI8019SU6gHRHIfbIk9NkjxEfxKxSxJT3/lRpwPXRbmUyvr38DdH1V0aA9MCT3miF3uNtJTZtXAz
qh6Ykk5cpabxINkdJbKs9I0HSQyOLJ3YLVIL7Pb8qIqcGQXcU+V84hXAutP6mYfqkhwXDvxRs6CV
flax1H90aM8iav/oZV0ukIoPhR9wxz6IzRfD5N7RCSaWts42cP+E5V+VIlUCpgxxIckRXogJsIhY
D1UiV5L/tpGuANsOpWoNduOmErv1/1mV2aSHw/w/TLW7U9xLsDvYZaqq5me5HPKK7bwBlEKQlHD4
aQMBbpHQedTlbgv7//45rIK3IvKjNBEhLGYrm6VlJDADBHM1myj7QmsKr5eFECis62Tf6xYOv5mX
fj83kNsdjy3q2YSh+q5uPNvmudvWL79ta6/4mwDeqie9dR3O9RUjAcDhGB4NAwi+ID2/M1ptgwFO
Hyb7pRMkufMLd+BV1O1jyAZPT5Lw8iGVGrZI8eKTAT0AkQVDWAQLN+1YHrz51pysHREHTIHZr3zk
eDKl1Wcszvinf+qpPHRpCqH8kfCMSGwhydzCiD4qOPgg4z5pGvv04VUmOvPjv0tMRasFBRDP8aP/
cbjqlhIc19NvnT132U2ASYlpQdr16DKhZ1gOxQ845jJrzBGzofjFjVX3SQxEZGE+cIJ8pnYJeH/h
VkzFkO93ygDSEb8wSiHCbH8dvhKZA20J5+gfh07Z9TciOf9tAJcpSb/CoqTPgJL3jCnyKG9oeH0a
qGdbsECz/CU85k9o6d8RlD1KQdanIw/WTUpr9M13XJjV2ri5XjFA58etrR0ce7URRBuspYDXUAkM
huhGmB1/amHJzmnVbgqgr8lj3kkirojRrdtpcuEzipcDw+MA5t3++U4H/0IBaRL1CZYk8eMdxxMi
Yh/GoBnyQHA2RLZWiMxh34IdSaNzReLFJi0BfpEzl+Yd/YMwX/JiRIEe9bNbmiStMgtAHlrWwTG+
mQc6sE95n1n5CkmabzxyLripCCcveYpYSVv6hZpJQ2XmtfkKaWzs8yUgmJVFWZGtpiFBZxcUkpIU
FVNdtt7fd41mjWVNnUgwvch/2LA5h5OG0fUj8xpM7m29Hwws8B5y//CL/sqJPfO1QJxbUA77Swp5
3PpkUmhj5p4Vn27z568WWNXaBWTJOkpGuW3aPBuNvitOqNVAGTHlmej6wWNjs+8lK2E+W/nkG5jd
I/3MHh3EqJNamYioMNhORMpszhyxDGWaYWTIRcJI5j4HJyK+i43T6vbwBHnBbJF2U/jNGRG2Gunb
tlEj5GbhZOPG+W/4ddCu4WPRVtrl45ISarCfHuui/tN2KbbkM8caz3gYSzNDIJfbfRuca5ycnRxM
pd6Ei+XrRvN17ZvwrwFcb/qkKL/YeeCEb3IsvkIaaq9Fvlc/e1/dabstS7b7uClo9exdjfMQmntJ
KHneByX18Jlm2JK185uiVAbWowU6waBvZuXpc+n6xormWx42kcIDdYmpSGYLNzFs1TUD/vSayLr9
EMYcCf87LQsU72yWpfYTU3qJwdAoShb5e16GAavKeVXdriQ1huORncAsifH+IUz8ByWubzcWVBzq
tiXNUCdUiewF5gOi/QpFN46j6DftdErQim5zEzz+RnfJ79PPh4bwiPDS3zJcqOJJNb4pifoU/pOI
sv3pB53Lj2Js4kpsiQl8kOl7grS+A2LnKgrfmcV32iv30obSQFvIhyOH4pzhDAs2r1Mz/ZNzWZNr
n2gSKe+ot4V2QLq6wIRtZlkNUag3h5u/zEAAZrlXZtCR/UnOdEZrepzJevPEYsScIqfAABLjPuF1
z8+bouHOm+vWxDntnU84DL37AHX7xfM8DeAXfInfNGOPYI5B0AC3e39hiQ8vu1id7BJLrwDV6584
e1WXfZgU0Ms4AiAUvn8BYHXAH6MJ1Lmg2xC4XQ80iYKX6Iht75FJeA2CUoZ0iZ3pvbFGzDhtmmxS
ANr8oD4cccy3FvhxiX1H9s6Weupg5R9fQZ9RlUAx56MFYSHAsHneGQzxhXlnpJKVgDBzT8O9U58D
kczfu0TTocX3xG5Uq/DgT0ZKyIoySboA6waCvbU5qYRcTcwCW316EQxeLsb5AE/NN158FmBsyJnh
8O4aGLvhexit8Xe0WuCbJxrHlr+Cl6Srw57txECw0aSFx+NiwxVTQgqW9a8fSbr6RBeWFwCElSAD
1G8CTYLskFHHz6oor+AZU891xP5lu0J6tAFIjikS+CRGFIjY4IyxVndKd6L3LREpI1nsEEtjWdVF
vVslze19rbrxI5q5QSNxCnhE9dRT9fye3EfUC5F7x4lSnivThdeT6mSzW63Kn5b48N5SJTe5iboo
HF/MrlcjiDo5tR+/gSm+SUBjyQtPiZg3/54FGrOw0xbEY+Sb498wy/oayx4dtln3QX6hi9TjzDrc
gG8mg1Lc7anCq+zt3kFhecYcu5in7EOHHNYo2GC1Jh/d4vFdfGJyGam5FnIilhBQx0RrIwN2s/jh
4ejCNQ8atXPvItTA/gQUMy0NOT/IdsrdFj+W9f10ceS5UJc3HNMTpbTZAgCyYEHFBH2XztegidmT
mDGQlbv9Sf13YmxCaBvPQ7ifnbQdd7h27JG9k5xK77yrGSVyJzwKJPZkvD5ohcFvkfv35/thcfan
o14+54Fa6QXhCzr2XGYhVwZ17JFyMZN4QGVEOqifNCFT3dG1CQv1CvcpIHBP9XsTYYZVHWiRXkvI
aKoYj6J5GJfbw8mtqnAVEZdfyDWzp+oZfdrk6OhZo3+YRtGCIioL5+fC/cXGC0H+V4yr6usip2Df
O8hpqyS+9IFENY5VJDj4In+ZCeCdnnwmC6xiFcF0ZnRQZ7yWeDMF5wwjZU70zTWAzh058Zk+2k2n
gwgmTBjj9jWYILOY7atBlos5ksHZCgSF6sFoqDfrnLe5XL4OluTh+icuGAoK9Drv4a4LJky9bzvl
TzcXycqNv/rEk34Eav1zyXc772BjyfpzTeMluiB5bRZ9JNQCFzwrFEeMnLfbxzGofauyugLWAcqF
5bI1U7ETt6LfXI0MuCF3mah6h2b7Lh91jTdOh7MBglzZLTftldJYFa1I441ZRDXNLpYQLB/iRhCY
ZZqfP5AtGqMH64yF+jgjdlhdBg0G7dJzbnsha6z7X9dH0kH3EdOXWIbbV9mwB21z/5aySyQ8H1ZU
YKDcVSlwCC/hhLZd4NnH88cSHQB49de/O7g14TyDlzmRQOtbF9Bshmc5CDVwvFoZcdBKnO5vhqun
6X2Oon3sawalgPURBg22BLgEYwWwqH/JozQPEiV1N4aTKj9yEXjwtnu7uGR27fWNaewrDsWMRHPR
r7MYC8Urfk3X1F7Yb3uRMluZg3J2d974t2eirbJV8JpfeZnVfWRS9NOCfzH2zz1hzgTc+03fts+m
68r0z4Yb3eQfQKmOyWPlZsKzVHqnrWdzpuGHM8YPM1sGFjdO5AnnRBb0d4tCBTOESHRsqWwfo6+Q
TmpwpPDHzeZ06QIFj8XSp9fIf480Sotfnb3ELXUVlEucwTnRvdYf7TNfUTSzsaSyuZUAwB5Z4dlP
8b0pIfqK48zguKvssSboU4HGP55HrAsv/A8NGZG28fCoVxAFqWNzn40J9PAaxVNWnf885OEXU0vw
pni7GcLENYrRuyd1uIxDiKaW5VE0696z6S+9tK501s6N+v1TRoqSYqJatYoobvCYlIEi8PMc+ke6
r5BVggcGPsgA/JQJa1wKGlZDmK+VN9j+O3aI8BU91bScjb16Cg68LuMtHJ7tG/nijtzi5jqb6g8t
1aVFcadpH9CvegUG3AKhilqPPWIrheDskE/g2v2jEmvIFb3qMRbjre8Vf3hELl3E7wbfib2/M/Mi
Z4Y/JMhH4kbtUzdumwNDg4a81eqVY4jpx5j4d3d1I0vPimKwD4gpFZwyhhr1xSvAKEsMHxED6KC1
+hS3k/dGSOHhRKxNI6u+XHFjnzt34OAGigBKi+gCQb1vonS83n51Ii7v6w7AKEknzLuur0P8Ioo2
/bW/VB/9Sw/MEVhkhkuCAzBilcf1FIOTdYAPPORThfq4Y5RRi90ZCHGuM3K9sIDNGwSly0IKuPJY
ILgSagFvnfS/1Zlr1Di2kaumx6G/zJgswp4oxDSsHlo9X1wZYSEjTeI785eqblntwQ6efNsTxX1O
O0fcBcvazc4IfF2EcBSYYUtZ270rHUoQNnLbM29kaiVXmdXfGLabbVSh34i39Myu/wkEVSS6mTkm
HMM9hGcDnCsVhnJeNcQa1xcwZn21+6m75zMeYNuDDH4wMv6SRVejzpqGDfNpb9IPgdaUChrwRXCo
SIUgBw+Tka5+VZPs7Us3rU/bY1gYoYzdFbZCDjZCtX+tvGa0+NgAqEjhajqf96l99EYzy0NsvOV2
FHcv7YIyJ66dXbRLR4ty5VR5bJVBTqLfNYRYBRaLoeA7K+yFR7favv3bdvnnNwYydITJqtXYGKtm
wpM/tobSienf6FaXYWhT8f8z6rzPdL4gG+dcCvWo1Htgl6lFociM8RlSw8jhg+vTQ8GXSFZyQ2+a
FL3grUB13/96JN++Kgo81jOZW00mWDC0blCkku16+4lMHtVuducz15IbxzOQ/OHg3qF54Pt43q1E
T3gYF1+EUoksGuGVcG5GUQCWRD8zz+aDgHYdwbL0Y0cPGTZ61Y1ra/lzHSNmuT6E3rto//HjM+Hc
W4SEIJzeeEwfWmXXY/zmmKd4ma+BlCG0sq9ppB+5Kvq+rLtNuMYtJvsINfKQyxiqW/9HrnolSHfX
1EDMnLh7T4kGLtTv/HupDJ9ZsSXeY+RMMF0nwsaqmmbci7lvPeEMWxq2TlPUiNheE+h7MG5k5LlF
FiDNqjnffXl70xDQkd05aX7RGFws69snwJRxj9zfVw7jjeX9GlVEQUAfcSBvniT8MgksG3x5GWhc
48iDooa4lhP9jKLxAdmS1eRbj1C3Y3P6NGRlXivgclO/4nIYV6fPsnqRucpcQWIXO70YqMyLlA2L
whWVl7prw6EwrplJ7VNGR3uaYi5PVt1wzvFtrai7nBYPWqH+2/aaxzaAU1NIqGgOafubenTcgVTf
KhqHVFuzxpgLzaWZd3JwVpo9qZLmgn/3TQcutnpfQLlVfpFIU9HO+ARFXqFOMGxFSdL3TleuSgQ+
s12KoChYYmxEjXkT/C/BFm9BEaFzSpE6smkbHCqvqtgV4LCcdAcWuA6QHHRYaPqVlLqBrgukiWzN
8Devf9E0HmcNoPPiKj+840SQ4QxWn8G5PE5QKbnXEYyTLdZP0QHG8z7hWtXB/v+qDLppNKPa2QDy
fVoaaCOgXSaMs0zXNtlKl35xGYOjVUJ+i5ynKloZn/mqOfYJC0M3GyqYmHQXcxtneJyt01OXfWPN
XnFj/YfW62tIs6fhBP+ufWmZ47mloljGUMfn4WkQcmp6G3Ib0E1I2/yXkC1AQcv0c4cFla2pWExv
SzM5aBUo/L2+RpcWJ3nmIkNOEmq+J56gd2MwRsyh8rM94J+WebL3m9pENYZBujmFf9clwVS7LElx
GtgbQAoeCa8XPXKTMPzSrJQ9A9042d16F/f1mEHIDzRoT823VDCvdx74gAFuVOPAWeHR8PFEgF+V
LR+aBd9ewceFgE1fHqV3SmsbOmPGFu9zQ1PWM2TkufSnpjyxSx+zFPQ+8BG9EctMd1TyqNZ02oGP
4byh56n4I2yPwjGBw+51IouIRCt6GbauQmJG+D6k4hxrZBLwQ7zJ/I56KVJaXeJxpmergNmoLZVg
DwPF5aT3FjeVeD7IFsngWkGnT5ZxtbH2/vfwGlDamrQU8rwomAj5YOvemkHoJlwUyvioyFcV6rMV
x3sjcGQBuCe0TPktC7uR06o4d+qz/ZPOabLohKK9OE5RE9Ua8uhmaLvRssK4UKbyJfrQ9s5ltJ42
ru8ueND4+JP//eSz0mM20QNEbvQ7FF9Ys3EcdXQay/VxHKgurA6p60LU3PtIqW1lkrpYvbGR2LOf
MnM9PpIRiObOClESA2jBl/3SLkZoakN7G2ymw1b66I2SJY3dFTEJeHT4UF4lId2xZDuwSatiyGif
2xDPzWvB/T7gDyb08OJd85whiNpSJMiqAXYw0Ufobwp/x5dsqHj+65jmo2my4rMHgLEFpvw4Anfj
H/W+1ibCJ2zhDG08eW325jqNTRe8N8XmXZYaJbLZQ+0q4orYR4dKTHdsaFz6PMEvyEcBJwol960s
EBhgdDs1bRog+/wwNFOJIlsvujCt0NppybuNzCZYeNALYAEPvByiEnGdzC0zZ/lU5yv3yHWMgk5m
QxxruYkVoVzLso17Gy23j8FlK6xsbDV9csqZ+uCeHuCxxMI0axeQwumVEbstqIvRI2hjzGU0epsd
M4KRuZ0Lrn20v+xsuRqn8xKgAJTJxqhU0hD1ImTgYgNjGXnO7Yxzq2wjbvgP1fqtYfli/p/VumQx
sBF4m0m2BnLZ2rDGURlcesbvOm9E2ImG4R5n+YBwDun9I3xsOh6Fl7P+sOg0PRHossn0qJd3bJQb
+dsJ7f2FcBxkrFW5QC5uJqitVmf0fNTVqJ3nnaos0IpeljO0smhQADYnPi9YAZlPmt1/A1BAlaRY
bLMAxJcJ6e97auvKS7F3dOjLZY3M3IK8fuk0I1kz9O92Cp3wBTkDMckPm1/iDYrWbu4RNK3wxTwX
jIfwlh3zJ20sXdGDbWrFvHNJ8ECmmCf9BNAgZHhl24OgIszWUNkPfb79OFbEMaN6inacmvI8KAPr
bpADi8svIIdyvu6yZ8/AQtrrDfoNf6wai3zwS9ylkzOGtU3OtDSt/dGg1vO13HVhsFm+mN0swdGI
QNChg0vGco+9Zka5OQ6zJ9de3Py9voZ0MjOxYgjUSd1+bhMemHFHQ+IBdqcVmGEhLtFh8+SPta/9
I7KwLoQkH8PPjtH4dFRTRuxHDy3Lp4WXV3MVYW3INt5Twenu2mhtjN7MhL21YsclLKQlYhK+40UY
LbeaI2oRZKWjlFfa9COhMms6miV/WiMnHR9YW/dVqH41xX4PVTPhna5+9Vyk6Rao/yBCF2x0A9b8
Q9WJmprObzIVhUlWeQrSH0EhVoHz2iTANIlspsrEsLajsGtirf93UsrN+F/z0xzrLiiEdaZ2JZ1R
4u02gUWjyBfwJxUMJiLg7GyKs8TEZSsNQZZLJ9HqljKiTEyAvH4IwAhsEjRo5OH6wqb0v5oB0ejx
bzzqhMBS25HjNWsm+wY1+RtAQRR2mHuu+J3GbiX4Qoh6nRSlQW5Sr/C0uFVobsee2lmE4VmXc1vB
PNhcLS97aOHkBRerWtNq9pznyz/flfONJddGeZWgDVtavgWEIS79hbVAMIl7NPitakqGbyytIZhY
sUwlIaA8NOtKQnH6coHNW1hWbFV+bAzCkumn6RqnA05QU0OP1WwWvwtvx5Mfh/g3Re5v/4RYH0CH
5DWhM6z8MRCyf2x4qs+36gtkvigZs7Mf6R71kp1ahf7ZIdGtSi7MJJWsUBDPVaAroFAgCP3Qdn1W
yGcN6CkzFz6+kDQzqdqA9kw9WFcYN3e16AmI2AHPONjrfZkrHwSnlmBMcBWh3rLKhZ0iuQ4wrTEq
hahkT6vbN1KVd3ZnebD2NK5oej+XovjeyIzekhUN7wPhrSMnVgi/ClHF+VrRIoOIVVl/iSXgBRmX
edo0B3wLBogY1ggzv1eON+fEVgsbZhrnOvZ5u2PqwUsF38WXe2QnnBWiafrT1ESU/1h7llYl9ZjP
EaYYEBb3VLORY3S//qE8zLXfls9i0YNU0RycAt1wRTSh61Avht9pHvgoSFVuoIN2feaVDlwTpr/B
/8Z0mI1GYn7Me0ZWmLZSnUnJxh6upjkIunlzv6Vd1g4tROKHWwS4KsMxvePc2x57F56LSDgWV+Bt
/U6xlsloAoIda34H7+VeXyJzYanJP1RtDe4Pg2PLVY6dxGGBUm0M/Mt7jw0ndHOqZYNqZNL3vvFh
5hbfq0Nq5btRq3JTmsBKkHt5sjXs738XTRBqYfPX9lm8vElsijXrlCQcsVRh3FOqxd60f6OTPB7Y
QifGg7gRRoD9gp+fZMZ0xbvCzkcAibJ8yxq6a+Ku3LUCXA79xd8Rg2+yZfRitCQBSyS6K5BsuV9H
wyt6HF5ewYbL3g7PRK2QWihLPRZ/fS2MvtbfY96Bv6oDPsDa7yCyRRAgC8MONk1YhrxzctibFq/o
6zL+p2HIfcLAlujMjC3ijvs1ZeZrf+sS4igUMtJILuqv+kH00zuWfXFAVJ3l96L+RhGjjseDL3fv
y9jXkxW5WRkDR/9Yv+K4ClyNPrSAGxeQmluYrnCl7wwR/FosLvS9ALWYT+Bzqj4bPicZKwUVyG/S
SSP2DaHI+f+KqJuoK4se6vyGZrnP4nWlYCYc0uFIvM58d5Fb9W+UKc+e2lwAXJbhBrCob++bFyze
S7MwtnnMpXTrMLK71KXLQu7DmdX7M+/FHuSV6fM7En9DBOHlQkpLF5OSPcaoI/uKSeaWvo30yI+/
G5ue24F1Po8g8QwfJYrsQq9ZMD7G23whNd9152QfrZTVOGISFzjtSUYeou8N4rmBxtyTVPf7fMK0
qaFikObztbpHphsmYcnOyhx1mDC4J+623HB2jdWR3hdFwLxLy6iEBIL4KyvG2k7S12/FbqfNoB/e
5pQ+r6jizt2NkBY4GYjhSXwmLo7iLZh+AgHiEWfJUxjoYNXSnXg/fr+GBJY7RY0B+oV2TzXopKAT
APfJSyFIraEiUpQ2T1qXm9pXb3BWwffKJqd26y0uog/vWIiS3ZKh0x+KfaIIIHeV6JlsvxvwkCYy
5CPQsw/9djFOlNf+WN3Xlh6Tu4vVSf9MgMpXrMnqr+bikaNFX/HHqTSf0ok2JloPjTs1bohz3Uq1
ajZWZnYMPN86NBIjNupLMl7JSwCSjiO/mV+KUQJ8UtNG6nEyKOIkMGijqspYVd5sX2hXR/P/75Zy
JqpMykr6VGdici4y+nYbHVOJX+JtRJ+6TRia6P8ea3iQRBGCVWDHbFo3Temvp4t3CMS6mga0XuVh
euFgiURWKgF+wuWM9aj3ydaCk+H2iaUN/hNVGtr1tmzR/JXzPqFJJJ9i7ZatW8nONpzx6OoJlGY0
tOaKfqbolsvfzwws0kB++/ZamjWqVvb+d1PmQLHGsFY6sOntnCsq+Tvjl8WdTVBcCUmZ9vcIdclS
+jR5wVQQk4bJEhajZPh4VDbFyZkqTW90sp1KS1oj7wNnwZ8dQhS7KCjQguoNkhU+UbJpeZzG1Taz
PUSdjiMca1+8MThtbXPU798TzFusFcQuVRxGrtB0RcH0WEnwkeaZ9kSyk7T9srCDja3hODEj8fP4
7oSORMvoGmopJSL4/fw3nL7DsOsSWXUhBYrUoEC9ffY/i5G9JUwOYwJOYLToD7mNTZ5wm9IcyZi4
seAqE4dKiJF9rzmm9MN6Ego3ad0Jbe1JvPB0TeqIoQFpKih6fTV/h6um3j5EEDwXZ8Znykbmy8Tf
8vutTfQuhZ9gw9dRVcn1/NoqlJKPe8yMcOP14KfNoAVTzu4YNDZwy9wqUF2W4JFJxzb2Skm4Pth1
516dirKkBIkM9/FfNY8L3WXm9PF7IpYntiYuYiSj15FA8tdnAJMz0HnS8FKwG7YKfrhcRodGI8rS
HYveg1X8m5ewIaZFrYBtlt9ARS4CqTVNW9YPSSca3/q+ZGfzyh0x0q5Ct4dJ/hJSIsIWHME0qnZj
Rmb6c26fI+2mvLyR4VWl2oGFg/FD02r622ELGftKI0/kjIG1RZJWrdun95j2RkWTfd4QqOWvvNXO
Utbv4Ar4EnrlaLYgwv6COeGTXogAEhaCvQqWVCtnV093wQZE6E5SIyc6AeXjSyrVFLfhlLMC37f6
nTHo0BlN7iLhd3FqeaaGAUxP8/7mngElMMqdTeYYno+OSiBmnXBO5L5fyYITGUTsA2AnVQxTwvdU
W7+9cNEN5MiTv/Z0YnQ03NRvgru2KwJK+3jv1xB4e58XvLFZy9QdRGzP9Wv4Z4zCRpUgKI3u+ogd
5Z3onjshURC+QrOzvJhYjmnTKV321+6H+ChXfXvCDpwSsH2z0cpxYH8fSJzbCoQMYpMpg00DuW55
9n9Ab40Q7FP2n4+HZmk0CiWf4sdKvNYpDs1RVUH0ZuYAIEfD7ptO3NFvqy56wuCPsqcTDutzGqTR
dbkejuNZ4DCI7geG/LA7Xiz3PvxDBMl6pi4LhjqVoqZ5TJtwneHFHnnMz3z/IZ90WC1HxwOItKW2
+6+ord3FQqQzXzbeJIuHOv6WbXrZkyX+3ew2XZekW/uIv88uUapCQq6nEG1D8NavU5DgbRgfwcHb
epH8rciDlQ8pwGai0dXFd5dY/oCvjVJiutJqtlye/NkIgA9NWRgBq4I2mvftemCZY9P4J5hT+h4/
RThfs4Ju3MP5mv8bUkqJ5aFHKM26tEYi3tW18wRlCODtYcxe2nIjQHMD/cPPfg0+c8ASszK6RMZU
tEo+20uVfdWkrqFH4izsPW0gfV3oaTLW9KUXHknCEPrixQqcFfM+vMnTSTgIIOHemdS0vY5wf7Mx
zwjz61n+5jwYeTGlONeWxwCWheCO89oJX7X/6hd/4VX5pI2z/OHdYuhL/vhheuY9s+tu+CzqZ9Nq
/yoy1F4BASo7bWh+d/yRcdu4gYBtJMVlGmwqwaiK9OP/SMo9zmKQJuMtWUckzdMFdKUGSxJ5SS8w
+R/Lj1clpi7JnSDKborWWrXNwPLyNMkFzvv+8DDLu7VM+7hEegPFDEPan2CDxf0a/qrDR77zBvct
WB7fx4vdYB5UbStrXOxBATL7bCyXaG1kIBwENIuGOR3N6Qj5AOwPJiKceP0cQD9X9I5leIcCj195
QsLrqJvrd8bY8GgBHSaSpLCUO9+auZcpzJKO6tO/GYTp3CPiWBRXKdtAaBCN8ixcfbJfJ8pqJdc2
y7gSXCjjamJ4szNRsbdFFceMTombWuEZ4AUkdx+W4Iu9BhE1MAzmepRI2Puh6KEJgooyLwjdMOnS
qLn86TfCxrH4gCLBW7e45Vso5e4WkUoGrTMR0EWaQF2BnuZPxXu+ETlnXHQFGsFQXFLdifeOc/24
DZjpyYkURPTlUOw8NMM7frKPCoLCLCwwQBInHpJskcheadYZd0DX2+zxTgYgek2NRpY0bhRxiQGr
2xJViQhtEjLkxmDXD7X2QlXIRPGkf5vCO6tTMqKRA5cNc8RaL+LLrttdAp0xhNAev5+xHYm6wrEq
ynlfE8lZMA/N+60GRJkUiOKcByBnjmqtHlBnrTitbLFJICs1FaoV2OzHK3bF7W9LzF9NEQ8osV2z
unf+8bazYTcX4LPw7Rg1rFwnWFqye0XscFBHSwTzmoW3j4dUwRtGw/DiWFzQhrmPJoIida2prGIV
eKlXBGXjfFCVfQQ36RDDdGWqNQAYSK1wnuq2aFsKa8APHV542fQdn2zQEApF2id9WoyM2Xpe/UVB
OsYa5bKCG6RNrDaPTa4MOLP5voyi2MNXipq+obO4HH+sAZ5A+wKHnJ8VImttU+H/eSwEaczJo2kF
W6hGnoSby05YhKtjMD2gZXFJiu/gmjEKPRU98RGD+QVa1tEib5CMaP/ZfpA3ZKJNoTrToggdRDvo
EYcFKDjqxj2oJvRf7mw8ZIwbePYjysjdhg6yRVjFP8rBejCucZQEpIRig04ghQEfRovr36uyDdqM
Mkj0AFZ6SvrfQ8RaG9d5Qo9xA4P/C5eJCBzT269CL6X8WQHIturRP9ORMVVt1jfmg4p9n3eoPv7h
C/PvZ87yu1YKOskq/Ldzeae64yJgy8Ki2AFT8+qmiDkm0VoHeZj1xHaALb2S44V7XLeA0A9cMMDA
l5uQFHZ0TYQM1jkEhEp18fmsOsJ54xxea3na5ToEav02liTKOcRq3k46DcHjpe9b3hb15j6LJkYC
f+xCn3YU1pvz+q6uJgmVbu4pgJAwyCKTG3iE+dWfz3AoGXwI/WUltNtJ1gTsWbE89VVom25qXxGc
Ahrwf/iqfX1MHfT2OCwF0xy1hDCE14PuAmqAm8Ewk3CiZS/CSPTpQnM1e5J6LbuSF7pKeTJqjZ3m
Q3SbkfQjSiGL3SsF2Tf4gMxocEkeYgF6ShKoCpPor73afkmqMmvJx/KsbAw199yMdzKJqHupIrYo
UodFRrqCwEp9piPwhBgL6fps+8/DvJd219Ex2DT8EZ7Tb4gQ1d3tW2mMvYDPrkYq/I9IkrHtt15x
nhbrt+zhtqij2zuul+gRL/hdvjv+uUl42RYtF9g4xF3o1Y1mKHwfu1KWM2zC5KWqUOLJfqPK1xHO
ge46JfC0mxh3fPZ/geW65uc9SwXPfjmYw36bJ1PdOIUBpGvugsp4zXvVCbjx3YgWDGIX3eey4g7x
eNofimr//i0tDfm2RfoNFukcuGmr0SE6LXbruCkWwSuBh0DRhaeAc5t0dGtVvelXNTmYkYJcNx4X
1ptdMomrLoDtXxymElPzXYRmR5IsEs9rZFQZgL7sqq+NhNydX+Shf29Oi0ZxkSnXjgjY9IaRpqBm
h8MjINKG/PDxnGBODa9ipmkWBCLBFpZOUG0W1KpF3ZqA7R4mFnUg0T4vMjxSktJaMCoJHEiV/002
nZR+nrnnX5gE9h/a6/LzdRR5JzI30D7dsB1kQF+K9Gqq2xo67ATVzej5KxAJB3SZRk3FihYIMLuU
BMQYkpvAWJP+LxVQaFJdoUAJd+36DRgHPdQGc0z/udymr7/P7FAFCyXc4tLKGwd+PXGhKsSrAmcG
FMdfv47iWT+BdJ2+TMlLOJtIINcR5hw3ko6bc8TbgSTtfsO7QtnivvXvTlUCqDdTlJM3ZPIK6iGw
8644qYLeyt1eFYYqds1XgCogmBTaLdlPp8uY3MW/Boos0mAZmAHOi2sc4/XQayq9PtVruhN2fVeE
B96ZRaajCTpCOR/Wm+rOt8NOxMxr5TvSHMOlCpZLybiXIqUYYe6Jry1nCtjQBXJnwWpWMwJaAi+L
KXhNa/i8KU4ynua1aaCCfwt4NhPRFRufDgprrDFwTG68T1a7KN85i8qEZ7jNSpt6RLxjxmMFf71K
ExIUD24Gv1bepbn3LYYn6aO66vfXuYocti6WZ+oL3Ds3+hqBoa8r9ujWCiwfhkXbN3cvRzb5l8XW
Jk7Xk3hXOnYo0bC4o33sdZ1nBdMGEwLat1cgcAeuwLvp9tjKj2sowBxrnF1H1AkFueFZTbtcfovh
MPjVBdxyBdPfkqpS/++XQRJkxp/nIc1rDkTBenNuPuqReVdeu3WuVseXikUIJRmWf+l8GVeOaxfz
bJR5ATcJN03GZiSy5uQlH77p9kH58sA+TeE9pQHW5ZmMKTGrkwvRJ4gViDlva/BHfgRJxuby/Kxk
NZImGtqGRnCCPlMVt4Em/3EgSadckBBhoRkxnkGN5iySacbTwJnAq/BKIFpJ76zS1w9jCzYxrsME
PKpyk+mnj8ie0xF751V8skpXvpj0Nd3WtZJetE8voGOwIrScOzxVvnugncnfzWli03HPuuvPqPyu
jwA8wNLAjh89Dpma4+0cC7MU7DUYg1n2ndbNg57NrgUZ2J7W6Re0iwSJa5o7mb5vsaK8qdLqC/4Y
xmvlDs7mVqrrtSEwRy0GVWJhHWTWBhIcP0VnOP+6Cxrccpd4idWHPa+bsUPwoDBaNQjcXgjmGHaF
nHQo6KLgRAv/wIkRvS5SduTnZmDQNwH18DkTMljungR0NFH+jVaQ0VYqv5woEruswXEMWEi35lLi
YJSXKJhTJgKaWVNfpkDgunkjyOgbdjRpGjuRk8FwqGMbSMAsZS7kO42TG0JkUJosjWp+lEqUVJAQ
8nbo+IvD5SjlCNIsz1t9D04NOUSu0UO8+ePvyXF0v8eHDcPtY06NS60X48/KRTsd3rTJ6wowXaJr
Mf0kaW9YeN8qa9MSr5S2CCGuRt/cAKJH7qv++hVTylL4+uRUndyfJyL3fItBJuOxn3FF0RY5VfAe
jT4BrTUeY105oe9hbtxh10bRgKi9CpRVWf/4JMI4dtMTnFPVoxS2OA45vJ/CSoSTGoO/Vv1Uqjyr
4OVyGz+cOvGUWHvxPg1gQRq+tT/TYFXtnmR3u0HCHkw9UOOlzLYI5O+xlyZPQ4zjTNrclME7kwGK
bbKgvXsdt+jbFGzqoZ022T8hQ5anJMBE8PGUhs1/lD6vyaGz4RmoRkXeynhsNnaqT2ivwgERD6zK
8J26I6moXyJV+jN6VKdOVsneMi07bEWO93w/04SOHc5xmQN5Ppt0wuV7kg0Gkk20FF1lRYXSCCop
muNcYNc77iu+5ePwAhCef+w/0GJnQeWJtaVDdYDFOId53zJqRqrRa7ik0TM6SfvSTXMAxHGgsQq2
sY3x3xuhP5J0QZTVVk/3wE9Klg6yel6Tqvxrw0beOa0awE9eAKx5IkOluiJH3vckAgMywbo2P9aa
qxDCzebWN2pfzlzYRIRZ7QLPt7xPSwthuTtwyCvNem6xjOry89orN8CBpy6DlTp9vb+fiHvtmhkn
g99hY9xd+xhz7JfwUuivZRViNgYGuoFUVUEUlYA2XSPEQE5Ak2SLUVIUPocuLluLzpX08ltTR8jw
N1Qx4ORRqwQp0+kXUj2rBN42K9OgpHiiDzuIKyU2mpML3OtBZBzI7mvAaOcArlIRxUlbqmmOs9gT
LFbFmB53Ar5ejaecXilROHGkjnu64BbPMzRdMCrEKt4pq6KvHE/McJetZT9k0GyYJro4yN4xfse2
6zxGby5zUzNqkFeL8rqlFPfKvQO+2r8nKoRcGW1qHXY4QQHCP0PsQBIT6lp0zV3VNeZG3oKF/kdD
KfjeLwNQNhaldicHdpl8kth2a3gMe/tVLP4N3oIIPcmuEHVq56zLP9mwKz7bPgo8TKyZtUAHOdgj
VVHBakVMo7tSaqGsd/JbFhVxl9PjNXGzZwbzPBNlFHVpRpHSX/FkYbZ61XTybYAGjMYz89Z2U9uy
vRQrUU9TA7iU8WMQ51Xj1WonD1gT/YTOcBXXdpyVyHr0/tSqyszozJEpkw6/IwdwhRz3lCwS7Gu6
K9U+Ntrik2vQaSODpY87cnrAQoBap1rDgHNy/o2w6ruO4j5CtYrdhQeTDKW3XpdwbpMlLP/hT1k0
fuXDmkkIqpW9rqyHeF1wDLUCzEwEfqjy9hN68k3uIfUp+F7huqJEP5mYNHgGLY9S8xNR0KZij/UW
V0EYqEpD5JI6W3IhYz5iC6l9UWZJwYCB5UlZ0W43E0yXxAu+6oReRioFF49ZFsuwhBmECQMBOHLk
QKT+XReYSj+RlOAHz9si7vANTCKJS9UDr9Yq6KPgUX3V86ZWTLmqPJBtVEdl60hUYnN4Q7Jfchju
PDvHZTYZw4/Rq9XpVl462djjNbN42aUbWfeFH4skFOY52/rZ30OLtktqkhFdB8sQ2KbqyBJKedth
48D1fIqOe0cakuJsAAuBUXwxDZ3wNqaGVysuL1PMZRmTPFfOfDGgfICU+ZZOihQiAZvpmB2wpokm
/u0QZ6fdMM69ZVPyx0EghkFSORFFXjo2vciUj6Ndqfm3BAVpMQBIWz3PcR6eCbkCEg7KEGog8DHX
qqNdrx5dnoK7NaQgtjfoiKX5xgFtbvquh6mro0yyIiy3dEJYl3neaLV0l3GuYhsZ4GbsKC/HUDNI
WtKcTd2FW7kSlp0eFg8Hhns1MqBU48x31g6iULxg7YsUMw/oApA/VpDkHsk58AvUvHPosot6l/BD
ewGQrSGKjrdy9rpr09Dq8wYWhgPMJmmjJXcQ6I8Ezy6ciakeZZeem/Hg3InG+nplK/Sl56LuZ7aw
1h2fHcAKMWoxtr+LOVjhP4YRN/pFLQjR3Hic7LB9CTn73we1BQyct+rltjmlLuEGfnO8rjbcGMDY
3nv/F4bQ9T+3HmvGMWG6bRvOmy6oONUe9pMImyDjOyMQxQKsvFFjfNJpTJdr7Q/rW8kz5gWS+4n8
eBvEWH1S1AR+j9idFLuqHqzPfCYIFPyZFrOAUJHExCWQSog+msOB80sh1DguUEAnkzCrCG3gBD5v
7Dd4xkQzeomut3p0ysSYplzOdo4wlpahb7KjH0ViMCn5hHXaYvYizjyZc/7v1zBAzYKbTT/uo0ho
21dL0qssL3uybhhpEAFR6qVBUkcnxGtvNS7oTNqQOAzRFi7oIogdiUSFJOyjPW09wonD9BpHhTMO
99wXLe638vmgxNF0clW1B/ul90ys97UEonG3XnugBo12Nb8FkO3E5tnCbuxFGkWKJbOk+m3MnUH+
QAbSc/zRdqIG2/RJFxIqxT3iim0D7fHdGq7n5Oe4kXSvTDg06TLB7xbSRmupa315UsxuutrsYjgj
piVcWU+/yVF70DWJIU6eNPqTZhWDR3twk63RkX0uYPwHUaDt2eTGJGj8md53UJxP/fXDMLZMqDET
v1KVjAdurRpYvEGyMVVl41g8p06rmcCZxgPGw++Nh8UMAPkmN+sglN/Wi2wSNuKWus29Za7HPYgp
Ut9hqJhixk3E15Hpn7C8YNjnx7g9YN0hM+hPW+LKqC2JXJmeAZs6XgApYvAjL2tEDO5BEancXgfH
n7MbpNjKO84dbHBuEfVW3b8WMjEl1zkcaLjQ3wbHEH0Bm66K9nRiTu8up+qC3HJ/04/9aLYPyN9h
iT+PAzT3+IYQ9ngCwSDQPLmklMvyEQoLQYt036lgCyUzyC6d+1wVjR/WG7Mm54E5CauOqO6ofegX
3XG9MkHqilbuzgK6MujZ6AY0lI8X0ZHGtzi4B5VyOakXM2ybRUuZ3WtgN2MUSKRlIejUvpXoqzml
QzYZlltdVD6CepPVoj2ekWXtskZ20j4NevBQHBhIQ9rok0gZl7bQX3TRu3TxrwZbnaj8XJB34AYy
Rcyh377fNc98Rnwm88BuNUKMWUtrBNeiDfY0RUNzJLX4BHobvfzpb8aXzWVe8apQb4VJSLUQ+NPQ
PQReOqkicjUp1hs41f0ZRpSzC1rOBZspXkDyKyqTD372Dvv+e0xMpQg82ykkDFlZETrhjXr4ZR8k
LZVST644AY5h4kKPawJmvRwe244myGaxzZbbCNofwlsLPloUnDoYftKXWxX4X91B4CnJ85aZIxVX
lUfqW5QVdi1l/vOMpt2MbGakDqMiHwR9l1EwutQrQnrKrxFEIgB046+Xcb/fD3S1KxQpyYIGANkJ
d3RkUr/AYnaSlTofHy6hxW189Q7dkTwbkhGOPT719+0fcV6fuBbJQl9Y3UlYEsadV0skGnmPVdn6
qQX3o7aD19xvEzMMxwQ/gu4gQY7pR6HwC5qAVfecoY8+9HgzhZsrh0n9mlTPuuxAV9jFBYM9hSuo
AKuVKbPVV7gebcvV3duDwHqs6ULpxdZyZYZUE5ZKABhnN/GCdfXxa9zwD/1SfhuTZiHw2S7L6KYP
4ywjY+9/NAKo1mp9bQ6xmteO3ae1AjtrPDpePlt0hvgxFRUg9+Za318YF94FkmkVvxnUe1aj4UwT
0+6YdaykWSVvlGvyEylaeV+9XAg6Rds71JcJ+sJ2L7zckEcd/m2Io+TsbXRdsVTOlkTAwnLSXXEP
ZKdJZj+Vv3rbVpffoTlxhmcSdV0xPyXKH3LWkhfsv67G+1ttMBxudWEb4TVv8ftnnTJtoWTIaoes
wOyMgGak1Zw5DYXJaSdNfCFyOuE1gYVdVedFjp8fLVDBpj/1v67sNssbB9OaNYk9SPyg13gv+waM
TvfRiEude5TF8B0MOAw1ozbbTqHwLGzCyfS27U4QrXPLmfOoxt8gYLo/H6P+jc+1/wjMeswdKSHU
1mG227jJREgTZ4I8cE72BFrhqYGw5dWnkmZ1r9hBSBqXfnQx7qTUqA1Ni/rFpgdidgMaaXKM0XnD
wmj3wg49b1Bd40eW4MhPUI7J8Q0bAkqlVvoN6u0k2iAeDE3vVvBfx7qZUmh3ZqzV9FNQESfxBZii
JIY/kOGtmqe+172NxxoZvLb5jHCDSVa2g6YuE7FETmSDmOItDNyCut5dsOflprJe8VF5t0kicVAj
pew4YQ48ShJkx29PxLAM+k1xFrqPOFSvKkKR+OSReKgQn9yFvfsFlJ8ox2N1x38gzn7+vlvMXDer
XZ2gD6BTYIPyPGn+3PiC8vuMolgV1Ql9bPFE3grB74OjqbK1aTDKOYs3Bns4M0QIny76Esdi4wXr
s2htOOArlQjbPA0lb6/MmVD6TiixVCqhqUAkC0f5fo6jseVm0nO1gxcnJzhBD0/aoDvUJ1X7M/UY
aZN6nBKvYV4+eZb0KKgFE+ia54RUGKzfEx1QP859a4HuwQJtygrur2HjHe534MRBkAfbOt4WYVtc
MfW4nbufKIEZvGufCuXyG/B4pC/l0whZGqUzIgYKSot/3EkjeKAGoMxQDOE2+3DBSnH3b9kYETVX
+XzcIBpWm/BB97Znwqy9i//gFIv0QXWzASAp7mlEnGgxh59ZYHr9XoIirEwhDnAB3RlNKj0ffYj3
UieQfhzYsdvcNus7qwjBEYRJZ63c/r7CINqq9kHXPvLr5zZnM4oFbRcI5bH1yVFFDguFqSuzJp3M
zX1O6Xlopw5ipIpLBGpzDXgvEoQbMprY2i2qBK745/LzCeqkUZY1r3fbge0EonumDdE2wpf9q5Ud
hLEVT8MRsGr0dbTRA5AUYA2Pd1vEOMlHimK+Uc8pqANBmktkO0ZgMbQKgG569F9GN1mSHYuIvzXv
Gu5Fpzjnb1aPHrwED0dZijVG8lEoPvVMSd7r1vQXdgmo0w2vMZ9es3o1U4tqjCG/G27tHKuDrhEq
1PF3mw2gguSOZo2xtBi2/6B9AwiA7wiwMxvgXbFg+UDhdybWY58Zlm3dUbWB7bgRXLqcuW9gLRPV
C+Id3R6D9GKAVziDNuYl1tl54kztF/9uhmzLoGTGSH/Nk/PjTKDmWXth2DQ1JxmcHZJ1gdQTYY+M
8P2Wbf7xRGF3FYbkcn/rdMvs8lmM7yZkkQUYrFyEjsb2yW3l+U9sqiDMDbroZQ4Tf9d9F4V+S+Xy
ofWmVquFn2x5EuytMyQxkYE8hWjmB4lJRGrSquT3PEOErNF21DqhI21ZWxb6SAzuyAEdMk9OuhBG
ZaYinbaSPX4Yx2ZCrPzWl2ts5CJ34Xgsk8tKjDnOcoIu2j79m4JdnQtBNIKDVYs4cjhPFlnAFtsY
TrZHMe6V2fGInmymt0gBllrr7ZKWTUsPHpqWk7MyLdy5qL1E0q1VVZfYXNLUmdK7E58cpFM1uBFi
3nvEWXGapKr2oUnAOHt+cm8m5VpIp+d8QnK3FWdEKlU6bv6th5yl6VB9dhEuLp8zgGgHCBg66F8T
chJ0G2Gq0rUZF5dx0K0BHPPcb1/xNwKQsNywsv1LLdmc8No+v3CoT0GSkFCUy4dOqBiQMrUFFRJ3
wd4q3BWYerUJK/JQWhavaVE3tgWkYPzYCRizym7Buuko4HZjGnAePXseAxC06H4JFoZ0jFeKz1Ea
Q6NEdjHdcHHVCP/rFZsTe9Rfo4BGILfqLRVRFWmZoEX/JiGeZgAzr+1LM2Dk5B82zkGgEx7VGYT4
iB9P2NPNiIl6BiOQuCbHSuMsUn7/z5B75Os2IihIL0WyvNGPJktlitnLM5iM56KabzvJANwmXklL
CgZEs4wT8wK30do7NHZ1Jd91U8721gYTXgLfxLOSdQhPtKsQ540PiBcHTQaFidq+9BWp0xNnx1kF
s2bqb0riJEJakqXBbMa95a7AYktk+vmm36zG95WmBGfRB8+9/Y5NgjGBvnJ9GieUWxfypWngsvlI
JYjOa3vnlwmaz4VGQSC9HmdU2g9RaF7JyEhCk8m2g8sg1MgUD2lmLH4cZord+tHY5Fv6cYOFPu1T
HeFCuuYMAlgaUYP+XIho63yXzfC8Zd/68cDTwNiZ1RqqzAIESmNdHwcIo8TO5QbUzMIWyxC3Fxyw
mz+nfKj1WV4VC3/4qsZGe5qCCJAmBM8bhL3OesnoKi2e329HSUUi8Ou056GoLRa5yV4mEInecZ+M
KcUqDE3bEpHKPU++kDV9+94IoaLVlw+KlgdC1ILlbMeTuvNd+AOymtbMhxW18ifVA2+wg53JIHYg
zLNAfjtNBrmoL734kWA7HPoyH4mty6YwvUZDHuvwlBTZPQfzjtaKgLAmg+ntRDt1FK76pIpQURG2
yToarrDnWsDidNt1UunE2nlK2m6Kc+sz9AvNnVcU75V0NgMIA1ND5Z3fNfNc6zSHfTGp779Jl6X/
Er7VCW8u/GwtD4YCLi1JNKkjfJlyxbQ82YnAxWEgoM2R4BDYdoudhOYET7w/m5HhaNqX/pAov8A3
/VTM4zjKf60XWMyQLC7GldiIjsmG/vWgIToHnIKFGaMtrWv9Oh3bdS8+D+xHHqiVuse9kfC/OSQV
eZFmeRuNyRLVoE6xjLf4PHAtxL3EBmy+VwGvOXsV48qF+PYDehOE28bb5dNHC2KVTVLX2xbFiwER
yqfoPdqJH8GmBGSJsvlC9+TqgIXXNU+VheNbpxXouC5AqxNkbOo6ZfAfDBd2OdL2FIgRGP2+nE2Y
8/DHJAmVfcsGkpFW9dO7JCy1f7Q6SQh+pbN3dKOPrIndH7RbyLlXdIM8DZvqhglBBMSe8cUOV0fh
jasNTORRm66MeE0bhe8+f0v5O9LqMYJxjf6mHIMe0AWxfaYzoueCRcC+rS8AQG7xlraoVnltfrA5
uLPBNQWn80KYhGuDLcJT7VDs6GFQMV6+j35/2i+re/ybyGjodE/ScLSMV3ybgZU0wzln8rmsHQtg
9bQgLvWJXsKO/+lsXn36KVGAjjVWB31FDAtKd/XRgDpHbvQFmv5pEvCejnESxJvs1whAq6Jke2o+
nbM4HjmESXNbAfRQ+zoLFnTPZ+WmU93M9lys6FZ7npl3dSPom7mfJ/o+JHCBjs5pqIOyy6Xdsstm
ZF2HEPwCZTkcuO9nlp+zQHSIoiOQymRKQHdQUyX9npYu1Q6NkZhuhZlMZgpDXR5PqQo6+mRwt4hM
FLFsDQjHFNTlp+jEymb/o4cpEgt+5ToT7+NXK34yw1Fxb6pZwOwv2usp2mMuNwaSeEg0YxJIcSz4
FzDMriUSXYOULQ0sNUk3d4ES05VQtbV6e7vy+jAvWYzNyWVfK0zXzVVgzyfbDL/7cSBonqLPa9Qt
DqCqnRAcWpq1h89YAF9jWEMW7zEDufVPYZRNAmJdaNXQI8TYZOuC5EGSkjg/mWVmrCrHc6DibsSF
VZZXhLSr7I24G1GQd4FigPKJBD5+/YLZhCf0OTr/ju0b/R+Kg3TycDMDdpUVNrfIQA9PS6m76X/F
Lakti+z2fWyl2MY/E17GLwDE8vmXmcnydJHxNkUID/kFBNppgiQHFKDbPZSSiW0uwjONP9+yXbyv
knwcVLO13lqdH6B0H9rPirznBeTTjgTM8yW4r2q7V3z03nIqnWnd2ZlppNk1nknBzzsSMYM+ww6Z
m11wtxD/W0m+CQvS72WjvBOgdvuv0zqOTSgUycP2ft9GSkaEyrCRgIiUn8OcjqoUJYQ602NdsvC+
LatN5PbN2humwNJc5yKHVbh8SPY1odMjaHKORS1dTi11qCbqh5ti0MEgKm9kgDGvdxQf5qjaX7FW
driNb6lWYv3PBz2zNYAMMkZV/H1aMEN9XWB9aJV7g6lFdxDE+0MBl7G2ZW7kj0GCQ+7BJSqa8YJy
DszwwHLa0/IbRFUJD/HFbCwFaIsuSl9xpxYLJDKp3zoPiPwW3hTfvB8J1piWJ7jO8wVMcQROSP1I
FouVlonMPuX91MS21mqK9ljBBygaspXxh889DwtYfSRhbfk/nKCffU+xJQ97ordDa/2WFmvE7lsG
QgTJE2YI2ES4qMI4mnqtW46GPALY5zyXHdciIOx618M1lp16SMps/oe+yCA2Vj4YSBMgeAUMObpG
wjPdsuD9vbw8FrXrzuOhpTWqd03TeBQ+SQT4lwCjZAwD2DiJV/NfUCuNIqc+fjm04uJqOA09i3/2
r8B5cgz6k9VdWdDGnJMmasPSOKurswQBAsUH+q52lWCTE1yb0sQ10wl/GgLdlzZLxl1CwxYvL7xA
lIssThzfbqwSi1oUYbATZ3QtgCmEXXsLvJJrs9J5dAsEsXNRwIrIEy0luomSPtwdufWLW9P24hls
y1xufzjAJ0IHKmCb4/+VUOFs8ENX82YvGmmUTFrtT3ZJUZFYbDw/shuhQsWigxbpsZjQXPAUE4hq
KKdZpV1p5VFPQ0p170qJ84PLcfK6b3q9Cu3xLNKlty+d4a7/HslnF9Uo8HkoDpoHjKVDFBD8DR5Z
EHfdH3kqhm3PuN4Pa8QDGEKLaedJPTXPj6T+s8GpUma2mebJLsv/JYkzGLeFesi77+YRFHRWMj9Z
YHtdYzp6c0J2kUUu+lNjCViqEY/TfxQMQRJQEqFqAYOLW+urxV4dT3xNyIOMreZe+q191VrO9yQ5
HgK/lW1EWpJSkm41piniTXV7ZDPmyKJPDuO43A93FkrC+TZw6X8oTRP7Fo8RfGAkn6Q0irDGyX+v
p7U3Tt1tB2UQcv1tM6k6uXbNdAAqGnIDZbQRmciU6q/m8AFVZxdYQGGbXqB2Yol6CeCwMqqR74Gr
+VazHseR1u87XPLm7gKjQKizTtATN2lVmwy3+0WUYZ/kKB5hua2iR6A5xqxE2zoKeLZSUyYJvfmp
jNw7uq8801K2r6LOh5O2/ivB90XEaaYGq4ihIUSAAHfX+uU3807skACOBR2jxzK6UzkLA75MRna5
2CX+pBmB9w/y0hNymEdoJt1xmXZUFyjMwcuFcMm5wL8apwJIy2cQgyJuKTE4yGmABDzCSdXpUpC1
we8kRVc2tviKlSwBDDNDFXEFa9WRO7VTaPEYGQmEYoCgioJanYhFuuK/x3Ujeh7XCjI0bN8vnn7V
roNFFVwvjtePPAvPB93Nd7Aezk+Rpf5DWHS48BgYAamrrfqP6zVN48xCG8Fw5lkSyaMfEymeWW3S
9Psq5HuxZ6f3JHp4ZgjB8vFnTLGi27GwCNvs9UCOBrvz4Tsy5JxA1cLdipY4Nmux5a2fXqzk+oCs
5OXcE75NWPO99r2X17ywdzqTMmKLXHUu8v37FTU7gpOSeKg6dYAKsSP+zqYwHnidq3HDSZstVkfH
p9CfNFo5YhTZSqvs9u45gKLJZsBfFHr+t0NWIzck0/BFbxFc/xCXegqrLX0efA3WI9TLcqo7w9cQ
XY62KE9PuDJPL/6TiHY6hn3ZxNHk7dhgBtkWMMQfmuCTi516tYZAKG4JS8vKNCoguLISaddoSvJ3
f9ENbGtdjralOArmRrvjGgikiEsQFX7XXB9aGLWNwO2bVk+ZyhsSchO1VsG+kAazVtZH4Uw1NXIv
qo1mexC+TcJtU0eOUHlX2Nm0QD2yLeQhzCAaKsfLmj5QwYxju4LTQdTSK1Bk1lZM1KqLb9d4h/Vn
l9OfX4pkc/gMiJ3ca41N4y2z/d2AxpuDp4C/36k8c0VqBlxn7mGsSbj74kZK/9KcTQtZuDSi0pWJ
zSS0zMI6p6JwN3NuN5wwwRT9gJJVpZCEj866mtGTTp9p9GduE7+z6PZ99rKHoAS3y0aAi5WOIEg3
Gl9kTzXD/L0O+qsq8CFEN90LfAHZoDz1lT4pTd1+gblk4wC2ShAPemRDeqOVawtWvI4hxvJ4ao5g
l3ROpxldwcblLSzc3eUlPuv2CzJzVxbgTcjoA5Pj1qB06TMRJX4nAoJsMRoyoACe9OcAfxUiruDj
xRVrUQ//oxQEMjAPx249LnOBTfYnIFOxWZ5GHjvTZSLXaZp1NnSCQwW3S9fn8SJRuc1UGRX3YRBE
NZxbpmg/1Tx/EOePw1HwkUKc0oapwWAWmKfBbAuD1p2n85TSHMZbunEBOdzpg9dzPz8oOhq3VnWc
4ycsC0ulgqnSUQ0ri6ESNHdT3l7YquwKUfweo+tv0aNiPHlt+Kuww2pP7ncrM0MGCqNABelWwZ7J
JA3Tl0GAGzr/HiYB4Sgaxz9bbzWA4nMbZo/5RcfndEQWrKYlLdQYkj6umrYos8ZoCHcRH6GtIaDN
ZX4wZojGEfpsptxOTA/LgR6euyWnpwU1wfIxnhKMfGEJYGFLfO/MMsLaHTD+jvUUAhj0qswB5/H8
i3cMedg5ZCCw7Pp1oGAD/QImlRoRcvmQYPJV3PS28MniE+StR5QObcWmVO1HasOFJcwEt4FpzrDh
o3E3wHHkiA1Oh0XlIbgQxU53ZBovued/sadiAh5GPer6c+OYHWvODo+o6yaxpz+iXSWXX5IlLFVu
ljNQ1/bAr7eLOahBaU/bxccn+pGzg9HtLc5X/mt7/BPfJ2Tn/8AUckr8sXbWJ6DqTCUjCvYJY7Do
ztfrdqae+Nc75MeKN1orTs1FgNGsoTAToqnD8ZvnkFITPAsrJhyVGuj6VkW3CdO42YJf+dO3k19/
mcr11w4WeBMwrAgz/s4RDQkqn5vpHJT5m9gug03J6/C3JhzL8vWb/rK0F9hqJuTmx6A3zIPUDA2i
62Sx1zPh8zIqiye9osWK2mRmTK7msCLKSHjxnDD+HW6SPYOyqqa0pDfHpYs8YYNP8VwggKNpTtrd
KDbBJb+d5qBlCKMpy+MsoJrFxTgC86XxKxxwXIudawwJc9YgXop/7t3S9jIy/bCilGBbiD+Aft/E
hk53ZdI2XZGy0LS+Y7vtyEwWZQnYrbLA370qY4sJmoCKWi7dbnw4FqjJW5dCH3OBZNPbWOwuZahj
WIQ39TfvoSmBKXF/hOAugjk/ujPbNx46DDXCgQ//hNnfMxkAbu5B6CGa/uZFW+87BS+IBQX4KP1a
iadP6RcxwhliV9ud10POSKeHnVZkOSiHbq/7qdsieT7Z2bY7xkSqenZYoYOkSOTGzEu20PfIVSJF
q6kdU6WtY5vUnLw7YqkLGxVe8LIhST2txO6tSo0QxQN6fRWQtMXCLGu04rCi2+RebtraH/K8ER3J
+206yuetE63Pf03c6qd8hVrcC5Vht644xq0r3O7CobqHJmDbGgyo+QUTOrDc3tycWlUuttVohQTw
Te/JXoxZciLmXmmUeHSE3oNwKiqFy0JQn9EyXE9zz5wCxi0PT5LokmnGfFnUpzxSuLfpjHZWBe7Q
DCuj4ebFd5/II8jnwJLY4z7q+CYw3g6HZAg6YMJprGILnpkWSw4KyIhaqeMtPsz/REQlTtKhXSTT
QRypNKbDRPskL9DCc36YGvxg7qLDOozeIEhZCkwx5bCKXnz00TdPGBxUgPr91N0WvejeZey6S0vc
D/UUwXUJOjF+7nBauLlSlBGE+TBXuHNnPnjX6Q1/IuJYEqkK73I6jJJwxymABgkFwT4C3DyWKlAr
tfDxBHoZ8Rnc1eG1WYQGhUhLzI3rYWVq5NdUnJzPv+eXconr+8JyOND/8iyIBPoSLOOZ5Vrs2p2D
ZksZmn9x4Kdzu1IejgqRK6FFbGjeSY/NqVeixbJ42FszKL+XmpQLOALOG30z5pPfZe4LAN8qgCiD
ZGa5+lsVocZ77wGUG3Dt3DOEC7Y8oCwRCDaIAiBhOmdw14gWZwr4/9AxJNxR4iTGH3TKtwFSB6Zp
7Xiq9KYy8z+A8xvIH87lyozrE3qiF49PzCNMK77nefWOawscRjQGdkxtSFayj6T/yamJJ8x3e8Yh
IF5VVRAqV/VOCjB4FUmTbfgY9aJfjW7b8G0koPRdlNNmsC7rtbabtPXp1vtjb46l/dphUu3YvPp8
EDXdMTPvmpqJrHvu9VCoHD0wvHOrjjyYCthRjZYDkqIFOb9LMmyBGQQytmSoLt1Hs3H7bSRKhvFk
9M5C0UAB74N4krHp+Bbv4aE1xSldRub5vHvqZkFyHUf70RfkCW3pg7NyWX4nGOshZ0loamdRhVer
2QD2XgsIZGDUesmvMAckFNqEdlB/8xHpWGKMqEN+jQ5mLCqs8cONdC/kOWJU0gqwOi0zWiKp1yC9
e9ISRtqxOAE8jjX5qYB91nPWa07hJk6oUiZpCRBPToD3xFsYsvRd1WHOhIQaGX6N80QPERJ1M3PE
mhlls3+WbO6lXPHvtSkeNgc+5xguoXHNYbdm1YrJNUohEs+UWPcVyCdrqPF047NAjHjcT92eIXbr
xswxgS+C4d8j4r95Qo/8loAtjEBR8o013OAipM9VX0gj2B4lNTS1JIaT+tDsP8RDgaJLP6MVl/xV
hIS/ylRJEo9xh/utj7u/2MQkLb80OA/357YHXtuBXdmkycIQ9vhwBuNwzBSqdydZDP45IKUA2ngc
wNsJZTuqjdHH7r90IMhsfJuFXjWX0IIqV4JFNOre6UAZOAcioITk/Aq1d0JGDPSEXFySELNstodh
JPfZzMHoClLiYq2BmfLyOL67BRSDiUDzm5ybLpQxxMIEBDMVCJg7m97STdcvJ0EJwjQKS/MBjYiF
6O6UHUzHe30dcLfpms+3iIrQWJxfqll+7nrmHjV1ipsCWpZapDQZ9YbXf4rGIFoLD3bQhFENIt7l
No/PGmdCfjayaW63bm2sMIVIWeJFP6ttzzCJdziYxqvVPoZnJ8XX6Y0US4z8qsup/n/ensljZVlI
7x6MUSjCuBraE8hAmC3cHRp9+PCJMcVXCnIsRv+XOH6DIyWA9ip5acr8K+QMrjegGOUzjaTh4l9P
iXfQgxPJTwBndFPrXH1jy7D6Vaf5y2q82dIHkXHFWWabwn3tKL74a8yBD98n/FgeZmKm5a7EtIXq
xjITl1QppL1so+xI69XIHxbQDHGp4zsUF65uQkm6OjpfbduAlNH66CguLWcK4T7mCGZw5d3yaiD1
DdvrmTdqwYsKSCHVH9G/Qj+SN2UZMa1aEMapX/42a4KbkESVic/pUHrdxRSBYW6sxlWHmjHaOHuJ
GoS93TWgpnZUCGtlvz7uWQ7oe0TYsT5G1+3QACFyF2EQZJ4GkqX2dVhhRDPBfbheivLgZuvmltT2
7czUVfv+oWPYbeh8/zeH8D3hjKPv+oUMZC/03FsRMQRCWFAbmP5prCCer+lzIlnPM64uD3k8gsu9
AZ8J9nsA/aZctYK2cOKCWY9mgXWvk8VCttj/S9WSUZxculpxdAtZWlD3bLRPKKyH+ov4tgA7FGfF
+q9mOaM24kT66GaMXTxbPyApOvEM6jmmSX4LdcitTo/pgeKIm/T0CDwQ4Qm0JWaBnBri9x1OYD3L
U/URbiFOm7JnXxwql09BSIpT9HE9kNtk5R9FgvnAfyNAHfyndLfslSdTi2hVJVxUjJeFHzJPh+C8
pA3WtYFmwWCElRo2/rhM8MDkDuCP/EEnr7mjqrvq7BRClHCco7DsTvWJgSiEzq29R/oSGs30Wum+
oee0z/av3JF6+O1eiIxzysJQIDc9apCCC/UHYlKRVzPfuJ2dkMM97RQR5NArPiFFGhbdpM+Y07NO
9e6MciR2k/M3OzUd/MSmKAf7mXt/T9r6xvXWVqZN0EwmcysP7HPZ/AHOSH0dgeZe5ZTkL5n2HIhg
EXf5OTdFNFgCcZf324E9SHJslR7zn0hTJuoESFBZixehj7Rk/J9hyovKrdiDGBStkqrqlSnBp3rV
kV/m5zvio1P1apEf07age+GWGwBn4ri0/l0qpN7xlVFL66ACufXftyYMJLlkhI8kiw9aZ7KndYrq
+n9BZufUjTUPY9KjNCrnAvB1QngzqmlYMDZ2jyt5MlinGZpXQdiU1iLo2vS4PCaxW0AItWSevazM
W3BAxRG/WPSHdPSreklxzKgu9zJq7wNzEj/3w3ja+QFuKqxt0QHYvkR6H73UfpHJqIUJdEpH5zji
V3DxNI0UK8KDPsnp9lRKXuTF/aXaRZiutSHWhxuTtPfMiBIN80HFJSXR0PfjNX2VJmQGzr5mR0eq
pqXIvZfSxLpko5L2xhJNBhAEsnAJq2qh/l+6r7A6X2Z/U9UDhdug4q6Tt+STOLiKHBsEhYnZiZvc
V1pSNmGA5qLaCxQBtfZyUBzNvtXGHx8srAlCreunRZpBXDq3dRZ8xyCJMHYFRC1Edd7N5k/Me5z7
oQdSbJS6rlIeMCW0dqaXczWDdjMQfceqlne6ZsL1bvk+vlzhalWjhNVhzwJfNOdEBHU1kdkTP8zO
XaBSLz9bbxlMiD8EsQRlyKyy0fzQqS/TJ+BqZkJdmbxZUCo+tj8IqRiBVUdDrOV6pJNHiAHdJ/4O
vahBCcHuWtDeoaubT5UOO+AbF+KnrNOBOJDNjvbuKcZL73Or19Tsd20x35D17GaKTMmAntXC0StG
3YMRo+AD8/pvFZfuOEnuNse9lbtN3jE+z9p7m4iTYq7bo3zMgkQIhwtTAmRTOaw5KuU2bavXs0pm
IC3eCy0V+/jtNbOv00z/FUK+NIwlErobMytpFZk1kjCrRJAeuahwNs+9kmAvuGrXfAhCPKA291vF
zh9BIYShEZGaye67H7EixHv3d0ez16bqq4PhJQg/Z7/XCtxiC3J0jznEZ18WX6mX5B+08TD4LWa6
PWaJ79TFenht2fOCLFRY+FAsm9qiryAX0jRdBq7z8Ok/bmcEe+4CuxYL5vUaLmPh+LRCRAyYeb+k
9lxYnPPhdTgvDm3oYD0PYqxj527c9WeOk63oIxUYObsPcZZYCnsq1Nzh9NkTKfNptxfyt4ywFtcb
bDNLVCa3fam94Vvio0t1P/yfd50rs7FX8U1rhgKVDGdKlEi5fPZBv99EIy2z0fx2U8w8FwZSaPvR
lIOJ+MEzV9Er4ZqIf3hAyZ9CU4zmDXkBUChRtti+XKWmkkklk5qQ/jezwaox5uq7+NtDFkPX8Gxu
k6gJe7dppxYFoFpz31FOvEtxnepbwzaXmJSohoO36MZDdrRPcx0oeCFKtSn1zsHzrCUa8IlCcHcx
g/Sru07nHTS3ke8Fz3qcntHFLPI4ClX8gBX/0wk0pf62c5jzEkWj7jmLbblgyIm0me6iJaK/x15t
PBjbMAoQhHwhxzAUbN1bWjibE3G1qZEpWhrqFTz6nG97Dc2QWRk/MROzLhSRhOADAHxaGyEQRGRC
V/DVlIng4LvHYbthut5DFneRJ0nhg5Wa3PJd+4IJGRJ0FtH0cwZ5Hv1A0Dz6cY0ccYZfk4ZG4e/r
wVRtBdXPVovyV+RvWLKwRw1PAK15t83VbHE/1wjThBQkY/uCl8fs/zAwF+48sdCzy2Pk2YOHpbnz
gPVe6BNvfxXlRD5OriYrrxvxIXlIVnTidh9DNKhFiBYRQR/WD2FeoZL8/KnWHbQZnbZDSZW25U1D
KDWtsZ4K1+BqIWfaL2PNK2amIyEYAaKIuwqQz8/xKpindoMz8s1wEJ2z/oZJ+ezyNLBkafR5m1vc
SL9+pbKb/1JyuGRjaQN28NnGEYtq8aHq5rXHwOYXrd4/OjXsCaxkgzqV8mt0z+c6FnA8APybJyoh
yfX4iD0rROdZYVw4wWmYdN/Kxmtb5m7JoHisfo7FVp99Sd1PdzARVuJe0HBS6ZSuXyrqlWFauPV5
yja/slDybD8KO360Dzcr6h/AetgU+hQh7Hy4InQi/FkDZ6EGrjXDu6paXOz6uCZ1dPTs/YO98VnZ
vJbSDvH5Eij1ODexke6KHx4A7352L7flDdZupqIWhMlaDMjW5b7OL7v2D43TuAjtRxMV0GKdz/Uf
Ee/q44EVAZUJrks34Rdj5rtDuRYrx2RqkCNfWPP/QYm/9jbW+dtrlI2zz94624fcbG9kTLqzIdGC
l93zavSl9/AMw2VTUK+hV+jBgTOwVoqiNxp/ik8pq9NC9TVBAnUDxsChE/tNLT5X0DSXh2upKRpW
9Jfd5NEZCLQcNL3enc1aR8cWzXRZVvnPT2eQz4aCEgV2wb/Ym4TuN5g5BfIy1cqWk4m2Fji7ajzH
d5IdJqJiDbNNXvTz2dGYgHUpPrLWuCckmlyXT6maRL+6qzxqMsXtgYhSKvOa5+eMIpQQ7Tg4X8bT
hfGZXX6I5n+NzY6FrLBL4dZj9+n6TgzoWiTrEkUlwY3Eua6S/s6U727afyHlLs9SSgoNc90IGXjV
Z3vQJpP7+2TpNH7J1MOgbUW2GkDOTt8QVVPDUJlbIVWnWoDXIYYT/CaJ/AbvmlF+MU8BZfRavp23
7pDh6c/JxNUV96aI2H+V/um1xqGgSuRUmg0YrIiWfXP3GBVWcwblIvJg8P0TFSus2REwwoFMfC27
ZtD0XPql2xxhKiDjBv39gNfBkiHSfZiAt4eqhuJgZN+q13m+ksTuabvybINYGEXappMhAc6hC1WX
OoyZtH+07fZ+Kkk+8a1njf2kTcAn39jeUw0bw7wfQiw3LL6BsA3V5zqjUm7W4OK3oMULzsV6UWTt
bhez5ZwbuxAyhIfoapcoYgq+CiQqiUtG25xTmnpQb48uiPBrkeVhRS6/jYNxS68C0WMlG0B+kH+I
fLm6WoQqbDagVkJDXHDiAOmLTcBQG4+MiqzNOIU3hH+KkfP1OP1EtKpaTjvTARgi1dv3HfNH2cM9
GYeXmyGPOuTYp9gyRSWaGmpF+LF7PbTtFw3l9lp9K4ZYqdzRyZDzgnOTGy6idgDGO0MRQzcM1Ch0
gAIZMqkZ7ZRiH5zVzltTgqf3MTSeuNWZGfXHDQKdLzsMhQsBiTn+oDVw4tGzeRlFqGVYEvBts/EE
lBzfJjWETU8PRLFwxqHQxygY0Jc3gPWpWIBaRHvhcLAz60kw3ZKdSWORX4vBTQo73v597PYDo+HJ
mAZG3EXWf7ZAKGIiw/h1MZZ4zV0RrszViHMHjvsloe1nYVhUuebqsqV6BcDw7poKNa3HWEGHVgVO
GfJr7nGwcOg6ar2z4o52/s8WzOakezeVpn2i1YUaAJ8mnc+yfDZcH2fHMEQ1JYOwMPrP/c6rM1Qi
+1wxVwO+JLCV/4TcYWVW2HWt3bHduQ2dwgirW/LRO6P8kiXtAW0/c70RdqpIJg1/oFi/CAa6ktxv
wZn5Cc/nd/yOeh16aavu7AkxrG/JmLp3DMdgpQUF5C4aS1DBT7mfiVGs41P7H8JOH5gwBt3diyft
d4JEWTcAmsGsgpRToZbrtLZMbHgxjuY2BAmfoqG2MiHUf0PQ2WJZlVcgdBgkEpFTup14BOpbDvLl
5PXGdvdQEXU4tTaFVMi2nANLVRF7jkSdRWFvFEGyGi/mIJ3ReotUWV/+LJPQLjGPMFfPR7uwVtvl
nbRypYvgkJ8rGf5mxnWpeVcfXBBsJtrpPVq6i0rbkZr+3xQQLvCRqdgpppC8gjQdCXQMturKl+oy
8RkTkso9qnDBzaOMl7aob/nzSi1bDqXr1lH0mvmABkWFnZ8YZyGQHK8fKg4X7PDmjVeAToi+v5nw
6bbAD7xcSiDqjsd/OXtbYC4+uuAJL1uBlaGPYdoB+qEhJ8Pppe19A+ctppiXYBVBFmdRg61ruL6h
VI5eL6X1jzDAPWQ1sdeU/UsEaRiZLomSHssfEGt7bi8Ky8CLrNV1Yz+pEQXMlDzk5gDCYjAMd7E7
fE236Ya6Yqko3JnYm2Kfsj1O2SC8Bq5pvn3DFhOWswur2eq7Fjq3mQrM1oRI6SEiaNyYi7iiVNRR
lvXqPwC+DNaAfuKmjK3dSWwL8KUIFEzkT80F4BODbKuXwTkwfKVpSKgwsf+RLxiPqw4w1ZIjfKY1
iynCdLN3jRdrXlsLAgOLiFc2noZBC6SDYlyjWNI3FDdyK5As+u/0oBSSNZ6us6lIIGywXiNedlA/
bLQg9/HzbLqUphbSCbu81hY3RsmUBQ3YMhE7kz4JtmZkbBhvp+AI4EWt/DUj2UXzvrUo8A1413w7
dRZKba5uFSMu73gRGKULRmQOLCggcaHss++UZ5AUDf4KPNhJshg5f4XNiN97F+BiRQBQa300gVre
bNz9TMN9TIKz07wELh5lruCq/qCSDFBt/2p5ldnsJTHEOHdjxNxfXaI3T/bcmipsnKevj5UNSahU
wrYMs+sTEXTNTX8l7a1SxKDa4yTOudcW+8O82hAl0IvjfUa8XQt7YRy712V9414Ycz9/XovBUP5a
8BGy2FDpt8Uwt1PwfUzv2+3zKGQRUstoCvT5yvxDSuhkW5d2qRcyKgiM8Bv4BSUJgYRYGv75HnNk
xZqfg4yPtR9WSYl+Rr6AWxK2Nj1egeuZfBaPHiMjDkO+1s+Yu6zrutoI9h2n/R8ptkQ1r7/HMypT
QINbLcFfYOZmhAXLw9CNlAlFFKkh0vghnkGjjIhvH+foD6whEXn7CCrneBVPeE/7h352NPHsD8bv
Y8eElWT0vPrCCwKDZhh9yTR4UyXsWACpO8Y1IGa9cUNDCB8CV/C/3VJnsK3oD7qgmOmGoEYmcu5P
9/REgK0zk2cgBODckhR28rSL+WgYdcrIcK6zokR0bYz/sWL3AQVmfO8d0zv8F+vEwDKfOmg7+iPL
+p1GERi/58d9ZoFl6fo+ZrqKA4wCKceN9Cl3iSGYqYb6J4v45L3QGdXg8d1rSBV+0Y+gFD4mxVqa
XK63zg6HIsMyp3ysk5PU4AkaRCQeuY7wLi4ZnyRoBPJjhpMcdBhpEmfVxZPltNfAFkDnjRWm0rF6
7vyfZ4vEEQOCuB+XICtaMA1K0u3NLdH01sQpg259vgLU0KhXM7jXuErVtXA47Uvu86ohkBjc5Tg2
XYyyF0q8Sz1Yae3hH4fWf2d6b0mEo+aFLUFTVWlMJPrLNglyDt5uAggBs+gmI+5Hav3Pt2CsmaNM
ZMwqVrCpS8fvW6uFYZyE1oMwjgj2mtj5ZammzDBWdqiOjF9e/a6Hh9K7baN3QDyeWJbJfcFQorrO
S5ZoQrGJoHh5+KbaZHV4lkMsuKeQmYBqFXrBEQAfSx5yY05TEIZ3FdRBS7/3bzQTf0uGa3eU22ln
/Fbkmj5kr5nd2fBseAYJIwA/r6IYHC5RrlHLUkA2Al6ZlgF4Xn20Ms4CEqJPTG17+OYlIS9SaPf4
Z87hahPXbmb7CHkzjrv1XH/jOT46epx6nXTa7Sg4+odsJXkdfxC/QuyWryTkUODmom44RcKfZdIy
OjYGGUuYg7ZFY02e69DJt2KqB1SZnajpHZwlIQtejTwGL5kLBYX+R+V80k+6A5av1OPX+gsMhe2n
6IoaHQyrKL2o2nFPgo2Bd1exji4cKVS9rOypPASHn9mXad/3LHoVlkEhAj/ZzvW/+zkQgBz8CwRx
dZe/qMNtn90cBCADmv2hlZ2vT+d+gEZrBi38l2B7KHSfugZu5E05MnQB0lObPUDLsRb3fA6tlmfK
KZLdt/FkUHsAIckKDnlxj+RABhYnhw/F5jNvFSNjbxqncTflb1AhQZOMy5MAbhYLyxX/oIGTDlfZ
pxp0I/N9vebE01PZAaxYhA+oYWkdHTGgOPOfqyEg2OzdWxw4Mu4fk5gPlu8d9wWDspAbFoNOAC8y
1szftIWv7+2nPjhmg0Y+cP5/ouvpg0LMs/5n7fWO00GBU71A6BwGJPrE49DdEDEyMELlgkKiuCCb
uRikUh1gKGK/lMOHqYHzgyDg48A5RZgsMOfchkMlkYKrQimMAdG92CdaodC+N8GSHyuC9ayYQ9Og
pIk+8xcaitF4XY3QjW2s99RdIZz6TY4cAUTUgO9A4D4IXWgjL7WdTOi6ukjAQmjYOCptxraR3HBw
t0Mc1Hac1UNBR7OIgiGtpYJJAx6DTyV8Enl/qAmUYAkudafWLmfVH+0dTtHLIs85r8eLRTK+DBxM
JCcudOLQzwZGQkU54Lel9nT7uYEBsm4zqRfVfpu6pilF2byQHAUFHbX43K1CpCIZ9Yk71ZvwIUsE
JUmpvDRYaFbGXW/6QN/HtHqKHqjtbtK1xT5poodn813qlhc2WW4QJ5izCZ7YaDDMKAlkoU+K3AQ2
HnKSZ/vZ5QQKHepep43SdfCRs9p5z2uJjW8LboBeRISLN0/HBSYjKJfYUgRFsUHSF+Yfmf53Pg+K
UbhCz2oD7ckRm55AMwh1PyySMuYymUypSbZzGzywW7xCg6WUylWK9q6ZLBUKZ1VVGZ/1STZc4NnV
1TQPzMtrFspwYDOdAoTjrU5io5gbYQFpG7BTsw2bSbyvTZ0pIKUKEDu1UGfVnPiboaxijXQuDHe5
MJvS8m87ACX+MLad7D6xnEI1O6E2g/ITuQq17isO5Mk6SEHql1zKDjM9Li5k+ni4FmuydsVN8r8A
9D7m01ny0FvgmjKEyw3J1hTeIc3xjTSyd/lx4savFH052Moz4eXqDDV3ExqjH1p4x8cGtKS7eODf
dpLgfChEDcDOzqiMzOVHDU9axaRbBVsSFOF/tHbiI8LOJsctyptdDUsf4N22/5xwsmYz562DdwcA
0A5MnPZSll2Votbk4skf3rQKLO/ZZxOlFrOXeL0Z4uY8S7aeifC3u4EUUQJA8gy+GB34A6SnN5F5
HzGYsjQ0mi2FSR3oMkUqIDX/TXH2JHM24QjeR26Mfyp9KD2wkDuv6O/aduZ5rG3/1sOKXr8fJ2UJ
8wq1I5sN5TYesnIixy92WtYZJsoHs5ba4wgDVPeV4sGR/lU5IawYy1jprwErcKg8jbSs8PkgDN6X
QD3pIqfATZMi1eKvkP0BoKCddU+YqLvc7zQAA+wBU595Nk4KYUigz+gznFsG3SPoLoqhxiU2xqDC
GtsiY856NuM4SPapYfhoXbMT/CpSCHTjGQKZOFWGktWFgtaZfv/fQMAr+U7FwNSoeC9if0jCCoaf
5pECBE+LvT9J7kXk5pHU7JVcbosF18qAnUo7EUh8WDwmrOvEojE8P77pDTvm0+GVdwy1P5jh2ftn
rfSDZhxD39Z8RK2bPW5dwwjkIYloLghPI5RXZJYlZXgTlLIfx23apnxMVE+3aS1JdloL1B8efd62
LotqOWXs5kKTYrFsFrVyznKg3Lf3WSEI7Z+acpCm/yvTV3wjx97QegEBbgRm5z3bNuTJo5G3Yn6s
4tOHEfUJwpAcSgCGNt+ExWnaNHEsZKEfjfhU9Sa+MlFQ4ivKuIr6ehaE0P75/llhQxCB2d6H2QqF
AKhIpS6cqbKlOnNCzN8ZqBV2Wt3B8z6Juvkr/hOpq/4tSqeXMOqyVcrzYtK94rd4KG2PE1/NBld1
Tx0hfwK27WMc4MIruMu7o9aDizQ0Lejw8bR3baq2xEgPz3Az0HMAfhFHt3yEIamjfKBwVhnuEJe8
dMu7iqMXTpcuPy+bMhW8QemmwcrClQhCQ2/wV6+vZziyq4Ol331sO8Fa7gVkdh0wawoBkKSXbJHc
9Ha4Jnwl5i2temHODlOfGyh0EnLA1VePmgueHcle93m/40Z4MIRfr4MCtGqvBsY+9HOxoi3/mAbd
6FOTm61ik4F43iVK40PDkB2jMLr30iahFc1jxd4BVJXsOZoQEAapZKIrTeunUTY6BzzO4Xgy6Duv
V9MlAVJJuGEc/3O7LIjQxB7xl/w3/bs8yUHbTC2CqEmdfgs0lEtfx8iHGLqFFtYwPVKfgO/fccGN
4dSUjFwrf52i1VpkpGym+MdAZ+ZLaz2G8GVxSzPk6fZG1w05F9nDO22jfgRnnlNAZrnkXnCBS6xo
Ipy/zLTpunEelFzfmKKS2IdjjtUgF2U4WZcBEKh/UgPzZ+ago0TkqEwJ7c+bcJjF/9Njw1TV5Hw0
JGBg735CkWBP9aWC55dI/Q3QeRYLWvff0BXgC4/Og99bp6KyrEdHHzE1uKsRasbq7tmF9eXrfUIB
4FiY6mHf7j/7n9Et9bVCi5KDDZqEBE6AFDg3M/VmP/63YRiLrkcAS4jp+GVOFP/5uPDuJVF1v1zI
RLoQaXdgMtdwgOq1p6ggvbnOnVXA3C5Ao4krLgejtRrnelNVbu93P7xUZeXO8aU9CpSbgXqB8PAs
uCkhYwCK5dXRX/TlhGDjj/ddTxCP0xXn0WFEEJzTJ+Z22ZTJ87MCiX+wWeJHL1VHNq/0oOKXIZY5
qbsstT7oVz4Rg57bb6kCQCuud0sTwxuJM47Jbip20fSOIbvlxhBRWQYIAT01+/h+jJ7GfZVEBNFA
kqIVkTvd9zg6RgPL3SvzV6AymzCyTHVWjCjUdtdgO80npyJwUl2BAZT926cG4Cj5KNPg7ylgzHM3
LiYFkCeIMOJyqfz0V5ZmTJ5LpRJwnGiB1jpgaWiFvm7Qn7uYRYa14ThyoWJ5mzwNSiqRUyKscSKJ
+uMWXP91pX3qnCxRj6sg73ryAkTqbb2mOfmGdezcm1p6vSEGtV8/mRPiruOY6d5gMPRqqe34OSV3
CZb95+dCSjiksCHQB9I9pjbHaf8nJjnSwFA780MBilVAf6XzK3eWfrjohsaYuvAWqGP9mwUsmal6
wNbdbUV8nOX3pLt8j6wehBr57VCDGOVLn18GTU5feLdlbC5jqQJSRII0R2F5CPbsvkJsODECBjeN
AZuPfAl4Si34UOGIhevU4CAxjfwfQkd2EYemxRCQinlC+1QAkZ/vqqlwbxeNiukVITdR7AWpEPVq
6spel9Rpd1DjTgAnDR1nHsrk1dUF3IyHDo9baYq/RDkLyd9FbPjnptB5hB5VrttJf/Bx/eLtE7sv
lC1un1QgntrW/P3rsSiF6aqQu5mzQf0SDGqa5zc3J/aYwJOEle65wZLqYDe5OIjMF/6EhDUlKAJr
GwtuLvXtOpEfrY2IWmWgjCKEAjju2F+6TRIbMWQEYbxHYP4CaKcIquNzx7KlJWYpkUtvp2uUbhLb
Iuq59AxeJ+S2kpS54k3PYxTEljg8EeUleVPpBtcrg3cuAX7/LgaQS52YiWzMn6xP0mztoIMI/ige
nJ0dSv9oDVdbI+0j0gh6ZgWa/WLKfiSIZIJbH425+WarqHuXeBSRXn/oE5mPRJy2wJjGZy3rGt9B
VHaOd1lrC99m/RC2S8G/7UJWbcfltadMff7MEw7sxHMDQJdEDLKzLKC96YCPw9G0gXM05d3R2CEC
f2NBV3er9ChQDZL1Ztk0BYJFvptKyhXn5eDKg3aYMM6DhseTrocit7q2zxRz8qHyWb6gKnYNTLSv
L7FkHEr6/eNzpVy3O0gAT/b5M/n6MM2jymKs+AeRF2eZlIh6HvPxX+rShULom1aRaXMXxKKnHcaB
zAC+QH8QuzLYojvuj+ap1ufT4lw7WOLyqxVmNdlhB9uQnoBwKZhlUB2eJhs/YqosBi9wegR14Be/
n3BYDcMxEKcA0FZ43eXI/7rPLQHVNN8293GGLNM/TCoIPzMC2SE6BzpfeRo+TE9KM8yCuD0oobSm
+LrPidvYPEDMB2iluHhSi4JufuTyXsettfq36d/Dv93VuN2wiI60XGgWcs9Bqm1J5wlPLPqM+xFO
DQbfVDUa1n8Ksudz6U0/GfENFVZYs+1TxggwwmYGnVqCgU54SCk9Nie3TDwkDhWxjZpeC2GruNlE
1N9/Ub5PecfcTCQEEictUiFy1onEU40VWQvyEliX1GG/6HQL2ateXjMj6OTgDp4TQ5DsjUYxUYrT
/Uzyb+tJZwmzubNgKYVLf1288vmawbZa6WuFpabK7Y9LxJUZuWHkPoVA4+/hDSr9fybu0dEtgdzs
2Ja3uZQTC9UfK27j8j15Hwla0EyTU766LPfHZ3zDYycYmq6WMJ6GEhRi7uSZkeXZnbT8ZA+XVieR
B7R1KH6Fa9E5xD00IJm0wmTitiC9g0XwYMxu/l1nVVey8It+oOzZvQInwZTwyjhgFR6E1EiHRTTF
N6/EHZmlqAOQoU9kOsy+h/fMsZLod9Cezm3HmMEAoJ6UggiAkkBRwtXsu5d4klzIwk7PiyKf+zcA
NP3SO7KmOl2R1E6Trmq62un+LTiDz2I+9K9pmWDCK3pr3krbLKVoMgnxza9Kh9VDUC5JFEeXG6rl
9J6Na6K6zQASj07GSQemV0FMixF2zNLTPI2F6ZG5n3Zghxk66Ltga/j6atbcKo7iLuX9NkdtQ/lj
QNP+ABVB59G72Y4ejTeNefflKsLSObB4ZLwIyZI4/rpRiRqeg8IsphYRuYCvRAbECcLV2yYVs+wj
NOt4m/cnx7fBC6tDbix7DH5tRMCnRnOpgG43D4os3TfjJAuvv9w/STbciXwHIJbv2gLOzzSTthJI
LFp+YWcSGV/wAb5tFSTRTQoz2R1RIWTArKVvOc9R4mJTZQhz1/lpAi4hYz8K8MapR/DC5+pIcOET
GWunJz1joA+b2486YmfBBNOVgTJ/eQd9J7Ibo7mmMnJhsqWlaFJOnWVdSargVNnj0N26DPanCSE/
hMbq0jRRh8OcYLqx4x3M66Y1BYZ5rAXFRRZz5XHzgFmP4TGd2yijpCDP+X55wAm8Wg/PzxM4sxz1
mufClU0vgeCejZFqkMBKh36RRdkWMor60Dll+K5J6hBhEbi8+9qy2jBEYHPtVkG8V0iqmQrqwE8h
XLnKQ5Px6AJRG+uLfAbO2E9mjPQXuOj2KNLNCXxr9eVnzHp2Rdh5dL8ImffzYqdoHybxW8Vqnl8K
7OaiN0TVyZUOGzeog2k3DIWG+CVW53Sfi+OyP7gjJfNTeK4qGh3E60kb1a2q7CVTM9unoD9kXiFJ
4YjVCWWxxf7Ytc6AOkiI+37UXLutVU0lTF6WFSx1mojMSjrHtsLmADTc7+fZwn67Pwv1yS0UXn6I
sZlOw+hdSp7KYoONS26VEFUJOVhC79xUlUSElm0quuE6QTBzT9oc703+TMCNOsOuGKfDY3VpRMoP
YPmkKM0tEWZTN5RnNJhS97TynKIGLWdPd3fmQeeG5rr6Kg1FEWzfP1FzzQ0/C74Y0ogH5kwXZi0C
kS3aUg4iAn4r6LwwOTYPlgR7jNJcPmKInHIuRSFsOMeQjIKB5xlHRH7FT3AbILju2SI4THaWJ1zy
tTA/MZlKgRYK/ci09nynLLJNzjvvLR/kwfiPe8SmnQLhv/zX2kzSyIpiuq+8I4d1GJ1wFyDN4/+z
zE+SpxNbmh+YvF5LvHdY+kdkQiKduGLe4mxc/o4zxt4IL4582SZHD2O7W7FWS7h/j6DmssH2g4Ds
v3Vwxr6VmMsv9ohAo+LveBF9p91HwgWHklqf+22ZXNXpjRTIeK3NmAteLq37LKNBTVW2C/okHgTu
Im97UofMQv3nwIGt6oZK4nPcd71UCkohXagzqN+KekJR8xHUWzO9jjm8RLol/fICb0t+icSmhse4
0VsGeWKVMDqjMdoIpK2yvOGYnDMKcp3wEl/BFyE8oVjzwgY4Pw+5+T2K+uLdUXs0JNPCKBOWvaT0
Cipem1pH84RtEYk3ESvo1TuS70+xEFZOLtFHf2yPBIHsUP5oS2+bHDnQMB2rEzhTRjnuGaxHV1W+
ggpEChzaHeV3ExsW/K2v7ePgkBFuKEQWqeFigTPmy+UrtpvgyTsfj+H0nfLnw9cJk3b5r4OgeF3w
RHuPaKsye6L8ZUP+PFbP4M+sCGU6UAObbiBnf5e1CfAIEe/kNd+q09mOG4iE/JTfBhy3Y3Z9HW6u
Ufsu0qlFz4R3wCp7YGZhXa1HEF+45GlQC0EWWO6OX1Jrk3IYFlieyDdaHL/Twa2ycmn0xFL0qjMk
WNjZnpOWwTGZKloz3oBWOvRtIwJ1ECJ/YAGAGHzIY9a7BhAZRgh3FbaPXQ+twcmm1aZVMY38se5d
HMpiICG2Jiv+HeDaI0aupXePt6gLhQ51e8ezDUfp66cL9RnAtNB2ymfkJz+umnAUHsOHUIUJodx7
1TjgrrYGJrd3gLjs6zltQ4WprHX0zbIWQbFlOQNtFX1aHQXE1EyKzjUB2M0E4ao+91uJ3Wj3MH9z
z7dCNrL3IYvwS2QZZi2+O/LywTg79UQj/VGCZfYOE4qJzEZluL8Fpf2Y2iGA7TCGQ0Fz9Ulq4i78
gAjlV8eNtVnL81H+If15E1mRJKKf2mJKJEUypd61+ZMkNLAHZUx2DajFeOu0kqoCFF+ULgOtXeDk
XyAuf1FGyt3n+hK9P2NsHU9VZNW47M4eZmri6XgU37Jthg4xWuJ/f2A21iS5rdwm8ETye8RvHuu5
VbOUsr36tgGCR6BPWQMiLRlUgHjdA9pvT/BJyvt7MQoFysz/QtiroKTKYSvlfkmQHup6SEbR+YqF
AFsh8EDWQhs3gUU0O1YE7r6Wrm7AbDQq7M2C1n6zwc5o97turAgftwUb5w9ZgL1WQl2QYhX8karX
KY6C2aWYvDYK5uiZOsrbY+MwnfgKaYvrxZDfVh4VYBhQaNzrHaZDfIFcd3Jys5Vk/TqPXXObGCQ2
vU6jz9+7a5BaPNVK2f7pgb3jntj5BH5LSBBsLIxgE2BNMMHzygqkAx4UFFO8+Oj19Mz529xMTbdL
mK8nlHkxqHb7Kf9UiYsmuBBe5AzYQdbXAnH5PRAL/SgBRPF15A6HeRb3d5Gr+O5a0y1+uJd7NHQs
NJgAO9bpjhla+3Ajhj4Uhst0s86ciPvIkhU0ZNDkZLELWOeLcCyoInbTnISzj5uXkb8LpVYMYiAZ
4fxKnJ4x3d4uuwr36xMTwCG/EYo/wcLkVu5ceeE3kpJEDCgo/MLMwnB8od+BG/Z5qq6XpFPgzqcm
vPXdVziO/4nf07Q8MSGYwTV5cRRKow+07VmxAXgr8RGmu+uLflPDGrKZ06becIDK/pge5Eg1aqc3
EJKkAHYRGu4NLMDQ3bS6ST8IDXJZkxnVVFMvArDTa3Gy4RszfqQ+sZtQ523LqwZl71R6AIQ8cOVE
mIFrZH8ekRICpDaHpn174DAW0s5DU9Z1c5DH9RkTZAIlt1qs2vYl+Eo7Vd1pvCuY9n/XmMif1jZq
UuUWpg2Brnjcx+wWUC8qjPVOuG1WfiNUe4k2mWmWw2yFktEZrNj0gci20uEi8QHGz7diCxtIaJSg
5to54BNrsDqPxkVH6SUSche8vzm016x2xwChOTTd+psGhmHJiyEPeJwodn+tNKZQGRCcLnnleaAC
4JmSz1Z9ASA7Loh0DPJxEQKHp5LCjBkX6s+6EuauO09B3pdPQcHaZj8pBPdw3IMZqeLNPW1cv4G2
v85yUkoE+4SUB2vgPlG75GWLjn+FcX3qSbYElbxYv2kfuFIYJv0SyN+R2anzl4YRrpsida2bMYMO
srskMa4tEjDG9CKlUhixg+o6/bNhJst0d4cS+pnKgRBxXF8Uv7JuTJB/J+8jzPlb9X9qFZnyjHZc
Xq+zHeLcARXInkFq272Gml3gP1yy6tP/HVGtAOjI1U/GV61KiJjtFpzuEOFXXtHXh5C0tbB6QDyL
/WrV3baGNoTLSifI1lk/eeWO16LGeH828rRsq+S0rayBfbSxad1S7/hd/yjRvd2XVpaRpkt7xCQu
SpcRhcqm+bNijZ+YIRm+ZuBVEg306oMSqMd/kaZNvrLzrMweiWfnPorvEfK68uGuPiuIy9zhfqVM
TYpqFrqGE9w1GdlQt8xN0fWcR4I6BzL53YJQfrIIKJ5APxsZxYySNH5+d9gd+LLfNdyQDs6b3IIL
R8ivR6sFlWfamZPmrGe/sjFxmfGRf8CDiaCirUXjDP8oRE7/DZFYBfQ8IodwJi298csBq/o3qt1j
HESD8ofOUWd+NZ5/IyTBk6KAwl94KvEz39O7VV76925nEqefKdiVItTHcDtyqYpLmRrN5mFLB/wH
IOhPz1zZD7TQwAbGKOq2GHwepSGgUsU91Ks+Sqh4AlruUH9WFOGMHJNd5ZmlQtNw8vzL9ek/PoLK
tMZqA2NcGNNCmowji5PtTfjDhoP4NygrgsFtNBQlormgR7lsNXJvaZboq8NiDpWaPT6qszrRG8cX
ujJrcPCkY4Ewd0tQz9dEYpJuo5EC0MJE4nIbogZme6rF22YqOlg+jwXt/o3s+sZ4lvDbvzIrB/8s
ImngWC2OOCe4ovb7SGLWAciTyDuqQR1VMbNkep9sI7RcUAJfkLy9kG6+tqlYbOId35H/pvopBX1s
GISXncmsSIzTrjNlArk86aHw/o4R+acp37PzfPOvrK3M3VD8LmSTkJpWyjXt9PQHZh7xNiiOeJWC
YszpOWxmPBPdBhht0dIdoQjiEYI8lDLDAqy4ase67o317NFArHNyLuvCE/qrrg5BtM7aXQfR3/lF
SMOHbfaYLPeLdBUqV4yfj22mqtleIVz6cGSCg784AzhOfFeuafmat0o4ecSeHey7Drh7U62RSUx7
UNMVBcgx57UMRhKjI4JvlUQi+/ZNbt5ke4OpST+LnDnO6dP1CEMOjmNvfaJPKkuQ5LO/GQd3bhGZ
7NXl232gNEGClG7SoLnZZidTVVBUnD+QAOb1pWlXZfKDlWSjNzoMDsnIXCE/2J/se5JrXC94fMVv
kSbClc7L4rJ+nI6RqFktrF2JU12Drb0n/RrFBemxZfeUjZiwUjeOXNloMNP5zGgDgoAWOmaDxHfH
744Wb/S3kSjjmBf/AbQi1+gdkJCfpaV86GQlHQ+aNFyzRVZ/lJp7Jzhrbt4Ri0XeBaBb3MkYND3t
N/djp8PsgwWH+vY4agvllCUbaPY4n7giPaiTRJBtubqWK0QP/v52vpiAaEGgvh9zBb4hyA7CWLsm
HDxWPLDkbzxlJTSYYTQHs7HNf8R+0tTR9kFReo/lmYP6JX3JUM1USJXFRSPSfuYdJ9aYMJa953QQ
IzMik5IErbzCmSKKh5RDTCGJoZ+cFh0Bbs+lURnYbF1QNxvnCN4iQ8svMTjmtQDvxB7V9uethdzn
yo3tpuRf5graWDaKDtjtp5+0GUdEEYpXy06L+EJGVfuG1oGas3ARSLf4BE1KhiaPsX7dRVpCSgaA
UPUNOZLPxv6X0ikV2wcu4MUWucnvEdvOLXWPiYVpthDqFy+eMyb95da/tNg5VjOmE2tPycp243o9
M+zsyM+gn/YwQZzVXph1i4UmMsx0R1gkrReefwwRhJVU0AA3yWyPsThKCFQZWO30ZO9XZY68Iu1n
bbEHwxHFujyql/aKzwgmgQgyef1lrKXDY6JDCJi+sAPEDtZBqGbeHkElGZykI1/ou+Rlb+5vICfh
7SjG666sg1INn1+XpcDsHPvLo8REvbHiDrNVX/QFXCwO02MPr6czi+l8Uha4579MRcfWxtg6GsQF
uEvf+5XXE+wMSumh6vkk1XwAG/QA4dEIbJafk7gUvujLsx1qUPojnlmhgLCFwVMtLtU3v7hRCkrY
96uxq4l3Ige5uD8Q57fh8R+lk0rT62Ak1+CfwtbcibObYpgZx9mco2xMYf3b/g3ivw3RH87yHHib
n+zKthwGAW8nbC+CqNzMTGQFhZo5S8yJ/IBUoWFaVVx9Q6zDCAKMu7nAwrDVwpPZnzYk7e5JRmuJ
fw82ofnioSJ8/E6GlBb9FQyjAfEOK2a0SQ7griFcUcNkjvos3pYNdJfy0xZQ1bszDEbEPLTv/fEo
NBOebwc3X/sz+7p/Ql980INM7E9j4gMUNC0PCp2jPPwiorP4l9kC0TXuqK7rs9+F/x3qrDZB+vmy
1ZSEoDaRik4KlYsJCtc9KivJv4lOnA7PLB5ap0hWtLHW0R1QXPx7BPsZAtkPEIopzeXKaUUUh+Xx
lyRdLABkC0RwJX+YMzzOmVoMxzMbYgGL/qdPK58xELR2JL/YyOz4hVkwHgN4ACwuKf7Q2ii2vbhm
nnFOzSzEuUQ8w4P5p2arTeXEnqGUdS0ANI+MIZ9CUsCYeyxCmgECssedrFsm0qBx0Rq2mWs0/+DF
fJeI87mX1cbjhnE8FKnFYvWVA7GdUo5XrQOzCGISGSMowjXnheVNrq8+WsTikacF+Hh0tVXLGiTM
wR2Q10so4O2h0U3xZv9yENc544OX/V6kY/faxER4Q0f5a7XIvAzEzSOcQREcsGIZrGe7wTdMb9FX
XbPYdku78wmnlLarfSWlPju1oxvUuBfkcgpgN2Mn11Y9BFiY4cUbeTk6CSGdeVkUBg+V8UXLZdY+
eBCKH6zaD5eT3ZAM05d+fPnE72p04g5rOmUO4bso0lD4BB/10Bo+1C3Mv3nfwKL/V0VjJUggSskF
Q0X3DWKqNW9e14zwGUQ4PtEJJEoAmJRvZrASClkCyYd8hRXoCEN59KiuKaag7/TxE2yayJzp431s
obcA44R3lMzQeGh9XM/zfFAOnlvWx9gQHv+TedSHnhkE1raBJkNMdQVhKQ4m0HZxqTgReUdGvu78
WcXDomzAlXzsujWdT8AtSYrX4NuG+w0S7xFhlA4a4cHzddxgma3VcxgOuiUmNq/AlAmfKsLEzUAR
Ffb9eXKimA1Zbh70XNJrFM4MdZS6ewODGiCOxyaFRwG8g4rAhep5dkgnVmrQNpfDQmbUvC8CYTF5
dvFxzXZJKeQW5Eo/33o68yv1aMooeCaK3gFHH238Q2oI9JOoyHnhVCRfNdbO/FqBPuttgePgs+iF
QzjXZrIvjNU8+Phg03O5aa7j2YGu17QRtTtoZ3AVX9cdKS8KS0btbo/tmy9OC8fqUWIe22c0LPxK
1hsNuOZdD/6b7a1QO78s0c//6MFc2eIc4F/uuKeojvbxtCHhkrelJohqpDP1HfJdqu+EzBupx21t
bsdAsTaqI8fO/frRaqN2Bv7be80klTYsQfXmYZHOEU5meQ8x1JSW0F/K6VACY/yVa2RQHs5oyzHM
boWfWDyu/o5OCvUYV7u9lBAD+nEbsgCEctBz/8kEfBhw3sVxJ3vy3HElJsSMunSMKJLXFKRA6ZrK
LHfEb6N4ru2WF3UdbfpecO0OS0UegZB73qydmDpzC2MNA7eRPpdJ0lH3TB/FLFNkjCe2l62IKgnX
/sSR5uCeXgwgYmSXTYp38gb81gHz9JlqxDzUvqm2dnGtHu+7GOmejG4Q5hZlt+CVnA0f4b86+b5F
6zyAUHBJzGkYfltk/R7vHa43wUte+vrCsNHgWiqXBo3bF4fm6S47MwIq4kNTU7mGXT4af2eZNJVg
D2H4oHHec1nLPIhtUt2m57tX24Il008imYv10JU4v7+bZI7NHMzh/JF3tzY/lKZEO9hxYf+4EaeL
QzLmKedzua+2CAzqRJhRX9SuW4LJfRTouKbi85UODX16t85zQP9Uy5QsXDDNSGnlOmmWrYwwRCC1
S9MTi5iTTNpHGGH0/QMKTruhVGRRsTuDbdLMAo9uqIXgywhuyeQ29DIhL6S747MhFll/E8DesFsh
O2DhAKbsOzlGl/yyn6eixsJ9Ef7p1b/ruS06lyV4GVzVi35AK7fPQ23kj3giJvPr7llfBksONs61
8RPjOExTSe8g78YhYjJny0ZXK4lJvsleiVcMTDyPJZXPYsPC6RHRB2G+4w4/U9B5OGbhCgfH+0hh
AHIu9RU2743kw7Kj+fmZ6IccDOZGnHsWZ1+em2g5O1AwQSnpnMMsHJDYXTFWRPk8L4kAcuuayS9e
WlDkSM8aoELFyhzyCYt7zvbmRwA3ASAJVZ3n87887uOQEG3RJocGZnivHWIOjhqJey18k+AVAOcx
9IVXChGJvcq4IbiUqMyp6rHgKiruTszFcYlGDX+HzlTKWAuJ75DRooz4l1nVny+XEkC1sMvF2v3I
mwgYqkbuCBpB2F977bjz8qK1qdTD4xuGCaRIRVhxrbYwjecAhBon22d3aOI0e//Lc2uBbA0K3TP0
6ov8CUWI+pFtFN/zeoLeriEYhGr/WPbYxTH7J4kpuaNVVOHvKa82Xoit/n9IUIdE0ka+6LMMNaPw
X0wzVTQUTC2Zo9Wcx9yMPLczjUwPfEX22N/3O6JjxF7iNILlFVfvpk6QJ8O7XxTIzQ6OGM/SHBmP
hKWDTvWTI6Vt0a8lKstYHV39QfxmPLhYPC1BvL1zKZxdfjYyWfK/DqNJHHnKRyzeKfNkRB97lDtH
3fiRLIm47VCLiQd2D8BtEkeJhv3PcmEW9J8UP3/Veiio77wgWgZHs5YqaodF74qDXllw0TDMVAQg
ULXRRhnj7hSLNm6PJ3LAT8kDlirJsmlq1MIjjBpeMrgyfycji1lH1ZfWMwEunT50lMHk/n3Zr9W6
Y1SbnadHQugG8iCt86R26MgaBp6rZ5GjYSiXHsqJz7vgf/5b1mRQHtkzR8OihO24oAWdg4QECjR8
MJhkHrwr1Bfu7llSswNDFEbvw6CRl1NRXSfnVjGXAu/9UMindyZensl4hBS7kDt4izF1T7YGY+zD
2vEz6ZZzOSD4YMUnFhXeQbXHD0PFYyORaKBMWorLRL+IesRxcKgqR8wFZF11cPXOtwXY6SPtGZj9
EsO9VCIamv4ieEV0TyL2NtjQYsyd9IRuPLe3TMwDJChEIsJJEccBErh7niZqAgt/bxm3BtqXhhYw
UECp8ReKnume+AquOXt1qFwbSM3CN9L6BBpIRdtWcb5psvodhxTKSSMo+zAGXX+DRZAvhfB42Xal
57XeGUQv9BfPCvWf3q7GMm4AZv63XOAgPusn8k/T/zvGaGsl88rjIG3HgccLaZ2aqJfK0iPOScHV
w8y3Z4hiYdeYJw426bCkTTOnhWGTONJ8goJ8uZfA6JcnvxksJio4ivgv1l9Te+FP8VaXK5HsASAH
Ovbd5Iwm4Wb/x/1yoNyc6XuCjR2MS2OyUNnAyG6CmrrITcBTXATtezDYJFOxl7MDCheuYqR9vXfJ
11hrfDnN+YG9aY0R0mS0WBdlt3GPOWjjA4pbmcCqfjI/1h6XDIKHab54V/6GxIicQJZ5Zznt7db3
mVvIGeKnqlX34TqdPKbxxYjcBiwBgxPNHbnIB/SRsbTnCPyYSz6UiWElxIJv3acP2lZK6rpSWHZ1
yn2/JKlXHALUdx9zfR9lZ+Uc7bZpPSUgtXIJPJ8zMpJud0V3ZrEst+Nqukv486jiH8QGF7peZ2nv
FjND3gQtZgEZfG9OxgkBO2o2ta827Lcr0qBtLG8Px3TAgvDzif3Km+2EzFH3rC8+tPrnOivilwxZ
2dUIqik3cvcxBhN+CYZ4PPw/Pn9/8NK5KpjZULcOycqaJhxXl4hjBJ6hFvwLgvYb2PWi7N0SedpH
jKhfCJ4RJ+H7nGLI88N2h8+up8/THEMX82ANCYNC40PhFT16Xoh0ExFV9OLYEk53htDanic75Blq
7oPvXYVnrwrs2cMDXMh8LZL5fPSThsIDDzSe4ndTWBG8TmfwLRQ49JXI7/T9reXWFGtlzV1GGb18
PxrdStXGh45TnpBT00SmVt1YNsshE7UVFahq3a4YVrPjZFzP+2LCPhMBtxuDeJhTUFblZovfJkHw
rEKgYxhwn25O9VLHsigIFpz5+iclVIcK666SA/dhMFmuMwkIaIwiz9EKhbDO433O7uOaSR+LwIrQ
dIrn46vnaDZiEOFvDfVmnvjYSfCYrtRZhfqLSVSU+EzBfLyy7H88i3eEjUxQMGeYD+MMLXusE6PY
Nol9MqpLZeTlSsX6UykbALMtaESLHmWpBMfhJFrR15teyqp//Xszp88UPioQ+dKvwAtQn3pluikq
5k3N0zZIwIOdWvmnhs/zYtz0JhROGyJxF+UMtOySIxzV6QQyyROzK96yrw0ssZUKwEGwrUiV2nB6
ef/GsnVkrqJyCTW0YEJHexU0uSx2cWHXjsSe3e/4zdvJfyCuSWLe7GBj0Se5qDeOGmfSMwYfu4Q9
eF2jxh+IGn295z0kXf1xNoA2xH67YGL4CI5zc+2pbepipTaAAlV9RSDNpxdnUODdSqu9nfjtFfqe
qfc8iEUn5834cfHdjXVAoLCKM90Fn+jfIyAjWnnm2jmMwwdodILyzNVOakHt8wtY76OUbVuMFUvk
j/bb9UmKclDRG0/eV9oYachcCgam+cr6XStPPdm8JhrftdXiU3ygN7eSPho5Ttt0hLDNr7uKYNxT
WBANfri+7Oqihm5DYNxuyUngNDfmFH5woQyLSiqCnJ9uFqIDAARDggYuOI94/gNay/q1+HD279hz
v9m4eVzu+/7gOIKvC2uVN5k5zsfsw3XfddotyxLsRuIAadZs1M00MdWJ6hjti1jqnxdELJEnXqPA
uOmxDLqUbRirXEbnWoRBd23HibEhzVORSRlJU1Y5a1EXdQ/Gi8xs/fUCxADhD6hVZmohfeiVP7qQ
dU7NUT1pbjf69nPHJ50j6/yoIq8Qqrwbt1pVClWG9DSU9zItqM6EB43qQQhhil7gmR0aSRVoRdYF
1R+z9MeMfokGKD2RD24KaxuebfvAfyBP8L3V5ZdF+h6IJfMfXBHlM4PdB7LgsWLhLDnFX9UZVdV6
Ut2UwDRt3TIiJP9q18mTaG1Ldo3drkTPghfR71utljKIuYwShGOf8lqBKDc+sLmjIN5S7aluIf8M
wFNHxX4dAtWCq1IYSZeqOdZS66Zw2H+o3EJIYmhGl6YAjuTmHGF0lZpw3TmN0T8F/MQa48MISuFq
lDXD+NuQz4ml/bbwfvnDNQp0uE5K73RKpLVlVIXd1t2raHqqmkfn3uGtEaPmhrHXITMjFPBc0VV0
/NNJkLa1T4Atw5mywGxBDPeWI3PZAgqH2YRMLv7dGRKnqL4bmCJmyIzGksgKhZ0WAYvvBzhVVP5n
xOmHhqzQXecyLioX0dIiWua/drDUZmxAFmvZBzCaCEY+TsCuFC5PVAns7dzzRnl/AdrKOhZnRlTX
WTzWYfda3yUObfuhQlzN4vIRIHd//3E6mwZvJWn8RZzZAuctJhP/q7GB/uDuicM297KvQeN0Lk1z
8aZs096jak+C8BDhsoUpHH1EQ5y72cW0rV0oPHBu0hXH0JaO+ihXJs9f6pCAp7HfzVq1NjX2b6Qk
YrW1AcLHOmTgQC/0wO6tDa1BM/YjtHSOw5NhXDNyoP1PffUBYXSP1BOuuWTvrGPx/V22FNgQqsAE
2dtdpyFe0xOh9YzIAi6pbCw1kCPoDHIq6G7Of9pRbPGlTfVDh02litmgJ/WuHsYZk/tSuxtM3b/u
tcWIuRYd/YMnHcGsL3mbXTWD45eHXDQXYiqVKAEwmwaDai492dSryaGXuLRwZdr7SStZnV2gaBAl
kQYHgqFH78fpPW2NnL9cISdZXhY9VX3YeBgoAWTweE92kA8HlVJLA47G36hQmQYlhv+/r7HTLE3l
83VOEYp5NHjQSc4aB8kdAR4N0y7PRaUGsDEzvzCKdhUMukqLLGnt4vebTGGX/sVA7NOVR/vfZXc6
rPuENBo7kqa86PzOXIgZEyBfPX2hyhDc0y4NZgscwsfBlHdjRzQlhTOAk+w1hA+g4A1baJI6ZrD0
xLJwbX5pXJ3dkNE+nYP1BgVYN0FUFcsahbMcJRSQQyNH3V5RuvH/VFKmlN9x2VzO2lQXa5WZpRTI
/CsdLemqrVB9uftCVY0caBwpLgFqaqGzsoZY4UEKWtn3NqpDhLBe69OxPU5d6WJ90GU2MPml98wm
PxjIAqCE+wTKm/IBihRuZYUfN2SyveWltDpOOFNE4/BFkjEYy3t8AoBagDHoarT7Vb0n9/pOA9bq
GsBCBicpkgXJ0D7H9Fon7q5NjWSCBj3onwm/yXwwTCoV4zS5s7OMtJlKq72etY98O+YkdF14tps0
35bDPJqMbC24sMMee3m7z0ptvAhEOxYM2TTxLYrJl7K93tHzFmUKMh4A+0RavEw1RR/Cv7TXoxL2
2wW6/wQPIEbwLzPLJd+S47lh0r+re5TGacmphu3GzkBjRZZggWt7pu/kx5AKC+8TnvH64uV3JNMb
Lu0e4OIrqUViQwy7ckHFu6C4qETa3AXcQPvBI0C8a1CmySRTQRPTqZrzPlR+VoBQgagGBncqIR/q
nqh8fIvJAFTDyVZefNdX8ExQs7qBNX+krBf+UsMcV51N/DT5qnm1wQ6IHnhjaDafqfU2l1KV5c8K
MehwICIBTLfcbqF4Lc9+cG8jd0dIrdS3ss+yamFD1wjPt2SWLsVd8y1uPKmtMDBdxfqjr0kGnL2G
l9FRjkEmdciLTk82ECHDmBOnWPfpRNC1/Pw8/dkuMPs/HfpWT5UwCDUGPxJHDtKNSYyGu379o5eu
azjkOzdhycqcVJGiEDAgzUEtsFSmPmQatJJBr51xsQAI9eu9eDvQpJPfC10MZirgD2fmDF13ym1z
reD3NjMWU/B4IGCO+Ccjphotet9Rh0Cj44c7TsYCoxqfHOanieI3mYI9iODhe6m/zP0JlQ8B5fAl
aVEXfGMD/oK81lvpjgoGtZKDwW18sn83So+/4Yt9n/ICc147Qhi1F5GGWlpV3RE84Sy4Q8FVRQS/
AWL7fuprNIXkfhHqqiJUOT6zJRjPCGCdFsslM8kWYGYqghjVr9lUdetVoSc01Bu6X73fcWzAnCzO
oAnB4hJ41ta0eQOW9+lElGJd0j8ohGKXjFKqLcr7rSK+1AEsFHRr1xDmEjl4AoS32xFjkidkEvQB
+hqtVoXwLcfjByZZR/nVZzJ/spYwA1ufaFF6nIbEmOHMFD0L1kfV+3bGOCdQ40UyEuheMgSCuKvF
AiNszgYDZHN8jki/90KocbWTEp4I0cys4hfc9Dy/YpQ2RvEIIAVfksbb6hqmHK7cf5yTen2Dc70c
dNIklTDG+3P790IyWNqmHrCIa2FkUmvnNwg6C1LMUzSZTXqCqixo3FWcF4IWy1dGC3fa6FgV85dT
2qqKZEieqriwYAiltqm9CeKZ6omS3MGfYfDlsqbsNARgUE7U9vMZtGbs/1HBUmYj68/qE5iS++Va
LoG0rP9RKhTUeO0+W3BVHnlsQmbUxCKy7e5cnSMKCA2TWCL7enssr6Qflv4VMWeRlIPMlSa0wuTF
faR6cbi2esQHzYF267aP+umJla0G56Kl4jqIZkNwLn9x5gHYw0L8UAKkdlZx5wrvQgJgs//+/UWo
Za83iwITek8DCfCK2gV+eE/URjBZXZNgGkdGj9uD+fU2OJOGkfb/bqgbrqvLTi3WCPyaUFJJIAvy
UWEIAdqGGZ7I+FcgwZE5pThT+CBPOhvwfTyOPTGSzinmtd7uGDSStMeMWOPMcNoUSSaCjyHoCa8U
YDu5FwNg0CnVDoqKkZ0jCQRbASUtROd+HWwSrjcGt00e467Jz+2dqC/8wzWSrLKQub8rXMUolVjZ
RM408GdGCJQyMEtxxRlHtGx5CWh2x0Lmco2SzpvDly2t+Pnmz+P97XCFJw9hoo5VB9oYest9PqIP
qLtdmGQ7tbADyYH8zHpjFUThsRTmUNBR6FQR4ZhW9xd+4aY99tRtStPXhfYTjDmob3HUJSAHNnaL
gvPndB0Ew1g2ufd3QXOJza7T3s7wa86ylHVSOH6QyWM5tERXjBddwRlJwieoLvHjUMMcWp6+3yyM
gZAlCueoSB4iqdK6QOgjfp5Cvr+Uk7AmP8Jomz/SyH73jxP9Ieq4Xe9ud1DSqRxmgybO+Gpdklax
aU2R/CqWq+O15Ar432Ekw8maTkvwsLqVJWOyEkvcOc3a2KmgfUe61gBloHB2AW+u9BaOIp93qomP
RX99QgZTZsxmjwL3ZwDmFjBxc4lJMeuue8fuNSmqbvSemne5kgnfkUj2iSh+WAJs466V7gnubgQo
yxv3NsPfLXbjRa5SCqbUMO4/mh8nx3nE2L/L6DQxt/jacISmwYv8mCpGr6vaAaOiuBMfyjzyhLWt
IgXpjGLUMGABbcwIPFcw7PNDX6fRj9VPLnjrZt/2gmNoYmL8GZ88veLp/cmag7FwKSJ6mNMaYsa/
rtjUHmSRokY1SGfLzuGBTy1ncmeOswJhKhyXCdQxCUbtoECfv+OG3BH89xF8C/nxwHkbuF1lE9Pl
JdXHfIrwmjnzG6udrwEWtrzx0BjSyOZccrSS6n8/gQ9jyzbef/b/Voj3mCkZWKYsWIi8/29454pw
LHC0+sXDo5v4vOq00172n3Piv1mtnJJGVgnBGH67H+ZlSAueq+ruUI9SzHtIxv4pRh/qXjEJZHSO
LquJblorlahzBA1+O6h3gahtb7D601Zcqc5exSmbmArg698G6EIKNccK27PA1afFgnT+lsFhbQ6D
Luy9P4On9QRcxVvHh62hqfQEOMBXIeHbVfFGqLzZKiSLOZCmUR4Rvwc9skJOt1VtvSEJp+rtIBBU
Z2XvPy4ibzMmG12xFoQ7JWKg1E/nma0E2uFpitwZpVVn+vOkpRsDGwtyNd8Si4wCI1y4TiziKQaJ
qy9MM76mwWUgItQW3mR28EOpkHPzH8IbYX21RrcqpSIoINz2ngBfVH5LF5+uZoVkUacsFjh6EEux
DReASGLsYE1tagba1MeSBwuec81HwGHB8Dte+xj52BvpgKOdV/rbrue7gWnbVsR+7U8h82RCR5Bs
GM7BtPPOmeriu2B4uDHKG/Vins1z7NrFwkxjJ6r1SKnttO+s/5eTY7c9x/MJaDV7LDRYjWPBF2G/
ZIMn8UW8m4OvpUwTW+DyEmE8u9u/DPvVznKN2zT3ZTTM7a4o9yOHZOqQVU8T9zP69V+Y8/p1heVW
MXcVL8L3J1AbaKpRZ1Hf4OoAZV+Ognc8tpyvRa+EplwyLE2C/hV8hAYvSv2QimHSC66v8Dr1sjqm
KJiHS3/tZ315QVacd/IvbU/MWfbFmb0NJLooQXtUOA1+EkEDgJMnR6vb0rF7imC9omf/Mv9YfHse
iw1I559B+gDhgnJSpIBiOur1YCr9kMOetknsoZuNazcu2dwKDuv6lACcHkYyqwp+7RTSniA06bjc
WCu9FsxK2xxXFgskqeX9E1iE85XEZX0md6naT79bnXeGFn7AfrOqT9AI2UBBl/1iC+lgkDIIrcXY
Y1jnaPgkKMGLkxdQYkNQ8VgL0IApK8fHpNuGT8tfv3qAYtmgu4nlsGLXvCApBrjZGAuwZK9eHAKN
ZqqMkdvLeDl7jmOWktvwM7ehMb9A0AqIpYjbFLaoB+we1NNiAx30swEQELfkjgcPI6RK8w1jALpu
CMpg6IhkthgqYulF14+KEVPPH60gwnT0Gn+bxEDHqP+IzxRn3dXSaP4TP9X195HE3ir3WS1oy/5I
Od0FnT7BkTFGumaojHOdH3tn5I/KpOn22PKNyBJW1msYwZ6+mgVvQ/nNKHIrJezbMMtQOLjTkJNK
NjnU3Cfa6r9Diq1myBVg7LfU0zfzHbRUBjfsczppZX9TwKcD7MtfAShqXcdXIixmUneJ/rdtiyVj
wNNGO/sEG/4AsqOYC2qaiYZQVrduRcpODXSwyhgoTBUuSfIkIUv+2Qsv0NbeLtIMqN1a6d/ISmNP
8vvmvJl5NRZf1+LuIptt5iioZ+w9SyIkyUQuKAW5jzbluibcqRBlgURqC48hoEV9hr3+BivxTU9j
yjBYoDo7cXWw+aKE5SvTDSJ3ifGHQwUea8u2vreGJY+cLYNrqPzH18mBr3EziYmNOICRrhtTDU4G
2KFTUDU2sTzZvnSYxZCh2Zx24QJAD4ZtMlxxx4UBFT95DOgRurwJX5PSyumFAMWQVXivvRzsdoUD
N/Af0bBstmAhqdjCfD4jVbM8MGCfLNrQ0QP/Ofy1orvw0dJR6oN99qiDuSc8ilnoIOGeRwqqgQQn
lCvVm0DpBIMqHLUJvMq+HldbZ/TLVdgG5PW38HbZSJXFJG+a62oHOLQcxfDfLWUpfmdKCOQRl/+e
S9RqiJfppRNNnUPmCpLmdS2aNdGr3DvUPiDeNeu0EogHckwbpEM7kEV4biX2SxN5UcUnb8LYK4pA
+6deDO0VZYK1Y3mDf/ybX+POrIWLGdAuCmBhQc4C0pxldWHyRhfASqlsitQcDU/fsTULLIV7kZeZ
iIIzhK5ioAsDFFacGPT5rwqLSROH6IEgSVTh71dsCGbYDVmZh4QEMXYONiVokfc2HB6xdEsOXkOm
CKgaUrhAURE5e34OvqlRK+84m0uk+G5XyFs3mpvJRPOP6+qFNzubuH0gvrwV6kaGmlO/Dhtnvcby
RAGqDvCrKtpN4Xe2MV29GL69f+vqibscI9SnxcI1z9T4I0MQU13+Vx7gFWNUvhW7emUu1sZ56Stz
EHz6YaR8bDd2I8k16ciBJVMt4dnJ/mcniSzefl6RsSscdS3MaojgSUWSjFhBNk2gudV+/Hm2W7Nx
hrx38vhovA51VqR8XLltsUILwrhNOtV+hmDN5tB/VPovtE7/G/Ap5jttA1Nw/eS6v4CRN8Eur7ML
T2mz8nI2RxaLnrXnHlkA9DADnXpIG94FN67VQXQg4C0Q9ArTeeOpaAQerUKPOyOafO9/BbaKOnuY
i1i547f9mhneIoHHez+hv/zQzwED2PRKmaolpvUR4+HyO07A+BpmL6sebRj8xwvOA9ZFDZpW/39d
0K02j6zYgJ878xRpXsU1525ff8cm/Tjg+pEFX/aeTXltXoWuCwniyPA+IcVoi4CRRgY0+fyzYIdw
a8R1KW2eETaM1bUvlU75CaecVUBmDQWHY6gZxfNRajCeKKoMM7D9GD5D8+hC/+kdd/zTxRXLttlL
vckNoO5I5yGrV7ZTB7GldJtZAF/xty90b/o1Qy9YRP/LZCLc6ziFs6vBmSP2HReIqnmB7BwRniVr
rZAvYfXEOXzoY0YRUYdH5G68C5uquC+dwNA2DPIFhu0iEUkGTbblltGM8j65fRgmTkszcRdN7YUT
ywq1cz6QLZdSB0eqLVTFH+WwZMd09/Ui/KXEAO28/KBcEL4IiNEp7XAoDFe2HcVGEmJlIUXftpJa
OEPRVK03hWy0qPZD08E+99TnC1cdeQ2RunQ7GDD1ZTFI1rpxM/UvVjh7AhNWh4itqT0WC2d5DRne
sbnGnuzIF5n1UyxNzNfmZdCL/aNSuuNFB27hUp5YZtKJy4p3ysEh9JXUSDp+462Y9O5cUntnumzP
xs0K0CFcqkXTEARtoSt3M4GbJRDDeteA6S0TSS7Y6/46PPFMKSrX8gWI8PCjKQM8a+4fy0uFlFcn
yZb/CjhVqbEMpng3VL0RPkN2+1UkCD6Ur3N5fFeoVz8zKtI7MckGknR2m5/ZKWlyi18qd6EZ8nYj
vzfJARR665cyTFmOsQeoqRWOd846H/EUUIepDSSQTyUhCFzuhz1fW1DGZvd9Un04LyfGs7/3aus7
/SL8QOqNEYdLiY+3VQy6suQC2vfU3Dm6ybmnJomoHurtrLSvbMvJWVB7NkmzvzIzUHYmYvMtcs5x
FIn2Fvqa1CmPCZJ9wc4aySL04BgV3qL6DHInRGQUOJq8PQBQK65QIuy3Bw94a9A8KeCO1qCjYPDa
puzd/KyOTrEEPP30bLJRuYtGfMFxBJzOZk1Rl3Tr4VSYNoV5uBjhU2XSwtaD/WPbUQMnaGRN0BxR
UFheA4gOqH3YyA12Ov2ILROtagCsAxVFy3j3UQyz+AsOskDiuFXLATPPPzoYHZKNYG6JAyNRi0fh
+/RbbekK7q9EoF8rYigdukE8e7os+15MtS+7PqDUdCLuqSX59UW0oOAyaiZp6Dz1YRNW7kTwRsGn
y8hEPzhI9XOCB47hPEgZVVNvexkpbFshnmlo3xYnQbdJiuJzkCdroM6NYxompXzYR2loCPmP73wx
m26BhIfDj4BBUXvemk6pdwXbSS5oU6ujqm6k878FKojWCygOl4pQZcJ15E9dNsTa990w5dKh+y63
tjjfpRU14AsrXyjBAGqx97VN876vC3kZHcpDH7WicUOvfA1FFdz4uUkUoHOA9TYOgU4TFbM77h9S
QDLzoUasXUpq1qgumsSwEE3ey3d4mEbShvOHltvoxpndkBJKeQ4ZSGoQ5skyPPT/BuFav+vidryn
P7sIj6L+y08tucdXjZQGEBihbHTHOLokV3ICSGJeVvMXcLlODZ6f5eos7/WVDhxlKbcIZb7SWgZP
3RKJkG3IUu+J/8x8V7fKW02vsCdaU3TMe4z1nk5H6wbbbjj9oKkBPYkM+8LHjt45gq8fQ9LqWekC
ojAER3pcy/9sD3JBcJHw7wQ8MzC1UGvQh7yt/SvchK3QtgNiopuf4oOnDzJa9n28qGJSl/KhLK+E
FbawxbGcnGAibk74abhBGFrMdl7EpHyMj/hcMLBolKxo/sX5hG2YJ6KBxaFC0MtUBrrr+Ue6ENRq
yqKfqG24YpwfmDdKC/WCSS59IiJZTwDoOSMEHkNXNPj2YzViM2JO9Ttcd0DjquKeJUTA7A7tpLwt
ggJT448kB2WrOSNm3yiFtghRvsZki7njxi4M/ZC0KtnJb0T0rrNZcS0dfZqv7GV9aXtqlRebs0W7
1+FvDEK0ocNDsXABj9Y6LU2ZNc+Rr/KyX5PFQC2+v0Dzd83z0c5rQBg6wxm9eQ/E5al97/0KDh1N
hqupdKXAf940GIMVqy54MpPfY9xKEpJjcC9dMtGj0/pCna//44NrUZCwv897Yu4rH6RAWbP3dn7L
kLVQtVadZgaREdhPaGe8ms/Lsv6GeagR3ktmKu0CAiB6rogTKUCoJ/n8GN+jOyd9ZvY6UicSXfVH
Bd71s7EY3T/9sPbBkOWSEJvjD6U2364YOgmsgKXoMtaXjPv8Ae+up+VvTlk/25wwrBsw3NbMnTQf
14RgtbZcWYl7gXzo/iaYQSWq1jkraGc2ZSSYrxFhIrKCsNqtCz+zwo+eza/x1p7Hzr6GhbjqHkKo
/ngAVqIBCHMJ3l8LakL7D18e12+vjg49jgLNZnr/v8UvWJGlzZvw07vScqRsC4ivcBE33EP61t6O
DOajCenLttZIMWZnyyWO4C87xQbZ+mEirhDXfKTjs0K/NRcl+duOR5Gx9RqnXR/xKg8PIqPv7yWa
5nGRs/YKesxUaSoQuMREZ0pw4StfqDlMN567LwD0TANTBkq3eoqgEr4IfVq4lL7gbrmwV8h2gNGh
pbL8UY1LO+7cTamI/hhwajpyYx+uNWOCM57OWvHj/EDCTlsG0bm48Y6vAF7Dt5E8ewiGzn0DCoj5
SP3yPhSEYLvOgW8YCM6JnnfnTYWVcjNlyLWo0zPXvWGeOCmJB0+ujufdxr5bdhYE7hj6pYO/hhSu
D5Zf+wZ+r3FynNPIepoI00GI8Yyzd73Py9nJ/F5CKL/jjsbJIWggaoJDO6fY6YhL11V/+Yyw1ud+
gVeJ+upKt/g8djee9+qHohn1wVkrMmuYjHz7go4UdJZPWlZz4lbl9kByUTA+GjuFJIUCGHHtBokb
qsM8kicjqDNs8nUK2j+HBARhq2QN/BkAXTK+oDIZS+DbbxYbXY2pOZd9IriQxuAP3ejRAyBxcEwv
7OUzMaigSDNLSJZM8T+HjT2CB/+ZKH3qBsFcyxRT52LvR6lFMGiRr6OXDhC69uzW2MIgrtT19yVd
+Fx/7kesPA3RUj6yZ0efEZHAbOMmQMt9Grl8LGGv0tBVd7qu8tfpLpZ0NyScdHIRf5TK1DoY1ZxC
awVHKbN1C+7tp3ddSesZnp61LcPCQ4P61oJXed08g0+FMqz7jBr2d6Lhxuk5Q5gFfQtC4Kg9fBhI
/tJ+xw3YacgtH+3Ce3AnzmTKiqUKZWOOtfK0Q7xgxnPnd0N/OsGDiPoP5UicAHp2gjbukuO1X6PW
JMvn9NqDPDQUjy/gyjxUgFxqPfmQ1X8SVl1r4DMXerlPRjpu49ZVsLo2sQ6NPEk6AfzuLwqFkFWf
fDrXK6Wi3IvX8lV5lruU6B5TFp0s34CwNYf3ccvxQK2JLfunyZZ8vC6FEmCgpAsvGGpTAYdTQZtt
URSsZCtWid4VKlWSMKWKxrT87dHFn3NES9nDQpSQkFpNn1ZKFuJFcLp8oOefslYUk3opp4UEyJ/N
bTW55n96WEIJYp24+IMBimgsaJrrRGdSzT6OCIUyVCU3/CmZXUBLRjp9fwpu0sfRjXShIzO3cdip
SVrAz5PXc0OdHJ1P0fEpwczjXjutQ+NNK9d6UllCARbEdlSAjCcTkgE4cu9dCVzNFpWuHjVHfvfQ
/sZpqu+W0kidHTavt4VyBguXWJHT8CweFyJrN5wXjpB2BVbMBc1SMhjGyXeHZs4+J8UrD0SMlrul
OD83kKMCVsA4+8BZoHNBZiSYqlp+WIhSa+PwzF/cIEfEMppfNOAe6WVXCTFOovfyJumQ7xDppme2
2Av5jKTLzML6Kpo0UUu5cpD4ZqIAWdZO5EdOgcsb85kV1ttLHwSFdh/jSGbPds75qHnFr4e1uS+8
Q3+F1Ctdy2+4lnZGu7IgixRaoVBI4K+n/+41H67P7YNZk49qLOZk5aux1WnZan1mWryz+tOhTGUt
NS7ft9KYFQ/ou092IRYvYf80gDwWKIYC+odRhsYLxr2Tvp1M052kEDFpHvqZE4D9dfPQY1BacYau
gSCaF7eaoFQ8ER76JSUOJA9rYzmPY9j5QRqBC7cvderq+V8kObpGt7f/9Zw4+umbVnkwBxz9lGMr
tHhj7MbGWLKWfuOMzUHdrGH0P2iWwJYvQAZzINxq0599KgX8SQNxEW1Lis8KJCY1HkvIxsBxWu+1
0zjjffJfp8g7hI6I2z2KxM99QWMo15c+vnIdTiHnBHLqRbVOhNSJRtdaz10V8FbMxE5gp+ZYoiEA
ttgCMWbHPAhY8zxCmamKm9waAEo3vHcP8MzD3i5PihEz14vSQX8nyalUOE9iFdcPdGexAd+8tXIR
zRrkSOI5J5Q4UgH9PefkWUYMlKKt8paFxROTPPILSX+ISIjEed/Xs6Pr6d9TlkwCB9cNAbiQZqII
Kky2ZmKRmRNv570rYr4p6f93vxbpiThGrvjtHIUDdtbxc5waOuaFvvOh0HmuKnWklxEMkVgBJOZe
YXRZyZ5WLUfg2nNCBbx7TBvTN5QOEM5AyybOXwihoXV0VJyKRB5v7D1K4wmydOvdsHDklBv+9xid
41RQov0isVyXYwXWkXxEQwj4w5zo7s8rzNkdOUSl8IMurYYEk6I9pSrhEAZMzrTGr7oFEpnUL2a9
wqCxb73F+lGL8LCUusxXVWi30CgEXjpfvicdUcJHVtKwN1CPmzU9qgbGlAAL9q8/xfAvQ8Vjmsux
fyl7Suh6cLbI4+0vX+9LyJFpPfhtpFBmMlFeY4JJw9/ExsXbq90ENIZYNXtoyiX33pwog9Hzv0kT
WVe4SucQbYWuZO0A4IjcvPKzm+6puZ+myD58C6wdplIgSTEnJlTP2pCGh4oZCtuahthnKozlqHzu
iKWUxdZqthsFBcOyCzN4GXdholnCd5WVLmY2ZF2Idjjbpizz6Dk8ge5OcHivg/mSRjH7i9EPJ/zt
iIrjNtAbqm5ambMFhQacokIW+sgnyDkGhHOC9lb2jp9ShnyWIZFtPOuFXOAN4l7P/mILNLOT1fx8
rwsEAnVLJgmIhhMN+i6+8wYOFehOqBt61VP0djZvDTtF2hSZmjaEAq1Jbeu4CdyTvujfAbqy2DLX
wozEuKj+Oy8ppf45UjCbBSWo/8fKUaEvKQzUJHOgwEEL0LHoRf+GugZteaaDezi57BbUqzWkWW1m
3RDlYAV3ZpcuapwlYKV4MTvMNo1NW0jiROMlUu0BhxRJc0sS5XkRJZYruJxXRTieSgL7z+q/f74t
dfonJTXyiCKHVstlDiRchkDWwAkQqavam43dcT3BXPnyaJRBNO9132afVWcqVn1swVHUlvAix5Fs
4iNdMO91iG8zV+3Lso9QXz8V42p53FfA8IGVZj9R+YP7pUOCm7dkA1fjcxvfApP0/PsIDG9E6chJ
g6J1aAzTxxeLI69uywsxdykX1vUhYkyfIWISwH5BNNybAN0ikJbGnLi4NLVKOfS8s2ypYEgmpR6D
YrZBA9YdD2MPhxVi6ZX95FDPq1jEaNu5P2YUxReOI+d8vPggQcOIgWwV51cOg4Ei8y4X8BNuZ5jA
9iLAsUsSCx4hAGgNj0vZr8briKZ23tO3iLl+cHkEimnz+KiasOEJ1EIkJJZrcl6i83Zmlw6+sSN0
0qeBY0fgUzMieQnu5dOmYJLK8NJR5S4kM48bH0NYix1P/cKDhSPqK1chvvUA9Fpjq3Z08SbBAtmw
IZ+AgoZKEkBUaEufoNids1W0t/a2+06LapgrcBkwGLj7h6VmR/Kp1mFAzn7KY2Ebw4jq20O4OPhD
d/HgMGyTYxZRZiZGwFAC42AJvyc8ycu1aCMDD44j9Fvv9wH1kjUJL8RENq3X/GLiJGknJtRwRwBT
tOZulPmD8o9GUh0Y779lH35fdbvCyv+7q0fN3r31XWhRfa3+xt42dT2mqO0AxU+2UhbI4Lf0vlNU
NbXD+paNqlEJcV186rAGXeTM/OyiwPu0f2CLflwgJQ0tj/s4W6JQSYIc/UzW8elFXQmLy9vhI/40
iA9qxgQmT0Lby18OBVOqLtL398bUmkq0GdqAAwXxJhvg2U8RpJjGtvpZYdwpLuS1b/XIyPxQKZDN
Gbsw59/VOkn0RNs/44h+2JZJpbRNa4pVXC/04lDf2ijKB1PxPqIcTqy+WAsQtNz6ZoPMbIhwWXTW
qeoXdnvck4k129hDdv3POzqe1OjLm9qvDNODTGAAfP9jCRbQYIRERaIdwE1ckSVu/wNPKENRrboI
OnPBeTH74aiUb3DPqKGlIe5nJlJGZ5zuS181IES7T0ty+amoi11KvoEPfVcg9iICN5FH/XaL+x1p
PIWlfel+afY2rdk/OgOMZnghU46mUinIDlc3q6fa7yodIWdHJ2cq19N9LriuUh1Ws/lNblyQfgT0
vFH3DgHzMvLIKkdckxmXgVIBhsngY6EeK5WJLui8YXCa8mNiaX3ogNQ7CE4eHYuZ84lPztwQV2h4
ktV9BOh1T15mg726FffOQLUWW6ENyBqSoDI2SraQvz8Jqcwlt78wNUpTTHE78S0vMCdBTWrQ8haK
7bDxwrzond4Fzbrsrz6YOZdeiQI1JteguOkwul4rz27dAqH/VIQlj5mrNBha5V0TUxux68M91Frg
oqLcTfBfsgrcj50dJP0gzhE90Kh46I4ID1422XRQdGNIkyqQuXS+4SY74g5KjcVh077m6oE373Dj
sakVqjzdr7FY8ZYmbnjMmkNAgyHIQEs9pr/jve4jljJS4l3Y6vWqFnlg+rkj5IJKuaVZ/Jg2vh33
BwZlKYyIzXQKtJLRlHwg/jazeHAhmgWAX6zQ/oRaDrYHZcfLrHmNtmJbSNZdOVYDnLxGEFC4Ja2W
8PFFFo8nF+PQfkRWsnRwiwAQW7xNkaqoL2ReeSbWt3QlKvobjVNOZA6oEmUJ9NpZp9n4oRNlQBKb
uRINsWCTHhfv6f/Mp0iJaSKh881XTjGhRQYY9UnO0XKiOPszFuwkXlhXTMdK/7XS0vXMc8nGK4ia
l9vEUlgwBq6R4WF3Hr8zGqIWuWrMc4BT9uevjqRQF7UxD1c9VbEQGJLf9/Hm+FC8xpt5tzdRZY14
QENzSiKFXhRfhwuhLM93ZhqAn3Qvf1ROaNlg6XFfguEr1pSG1ouFdG6dOVlkWUaavHPdPdYzxvc1
WM/lgqevnMgCLPs1dm5QQsAM3qkJXd6jKkk6Oy7flujm3j8GGe74Pnq05r3UdDufWOtL6nuqrobE
YJjTAG0LQNsnT76EV67INRcVVl7d5zhmDBYL/t/hRURs56RY2LQ0QV9Kwkt6ghSbLGCoBF33PK7u
Rf0VZ3hhaOMLXNCKMBzn8iU6cotHgYOYn+BzmOvKZYHPcFEhgK9gIzmnQYGr3GJDTMOXlJvrwwiG
y55uUwerNrJAvP/V9VngZdEjdXOSqc3RfKfSQV6GeMY2z7NJoWVbmt3+f0nO6k43fobz1ZD45Rw5
hL5GesgXomG5SAXSRDDIYNuvHFqURxDIv+eod/5Z89nrdDUiEOAEzFByEuNHz3T9a8lykW0NOGEI
W1m8gUMoqMy3xOj4pDIHHEbqa8XcRtehLSduOaJjrUhEWgu8wgXnSjX5RkzO56aX7U831wscaPkJ
Qzm770cChfkELqevSWPHkVDd18f0xWkV20JTDWwzIczZiErlic94x3d14UQS3teIJzcLZsKJpbfz
kWTs5PWc5OGBWayrygn6OX4uB76gePH8EYZKTOkkb+1mzJnnvwChb/Gwzs//lFDqzFio3kBEX8f5
qi2a39z7F+4879kSctNqCyNdv+hr+UbmifD8g9u4Hv0mH925LLhqlvTMiXw6x2c000Jj4riC4Rh/
kkxH465nyFJESEVwtkNZiHuXXBKNvJTE3PxmbEfPqOGsawPyxdbR/BoUWIRpx/c3003j+v6+PF80
OAelCFMIPq85Jk1+/eqfQ3mEfjrJReRe2bHlXlUTyQdB5VZxj+lXz28SncPAk/CGpvuUN/n+YpQh
BXJH08s95iiUN1qZzyJFKDaZuEtPI9Rqcfs3U0dEUIy8lwiMAjRWOCkOYYJ7geQXl8Q0bulcR8MG
C82HcSI/Al9fyq/tTWHIh935EM+qEVrX10y8SQZ3Y+nYnIvWwDQY16OnyujDCJLCNJchxI0JVqKp
azwMpu9q56pHuTIdH5oJJzSVhwKLtqlIoGMDxChoOBXAiA2fEWPiPih0++jHZ6LtbZ0Ebh+mttIX
5XVgBd91DC2A9RqHIFvNGQ6HCq0g8bQc/T/UBrMBQuTlJ8/19ze+G1uB03ASRyr2GqqXhqRzSpdB
bkObaeDTARd7HamJcX/l6OLWTPt9D4TKtRNiiL9XFe+Ipr4jDfB13atMjg3U8rclx4oASstu9C5c
nWKcQcasv6ESJpMjy4VyKLrJpyov7QqS6fwZCVYL6iGKpxTS2vwNjZHC1uQvpJmcqfA8k0bknaZ5
heAnopSNp164vdMSC+urq1+wl8uLnpAvVrFg1KAbbn3kG1cv5tHLcU3kfamqK7Y7D+tY8AkI7Fdt
cyYa1Gx6vEqpTaq/yzylmc9yrkXaPfuY0JIA9gVs3uw/hLJ6kt7AoqOr0YoTl1JweI4RQ2CzpUxu
ZNiAaFamSJUi2jk9nrFO59v7t4bTBEguNMN3TWIYyMJ7B0Fom5y1czwsTeiMm3nrAPk9Rp66VuEJ
oPEyC77soyaOoiwaeiOhSKSfomoL8top+cxWI+FxdzbYmM9p1QlI4UCTLIfXqTLrDnzmX/Mvcj8M
F2kUmwSTvKCBFc+/gp86keG9tdWljoFYIm5INErvQJbZr3V4VH4uR0y5EH2o6AAJ1JkaAhhkoAb1
OcL4neRszbJ0M3RZpTHPpiCprSBhB6hX/4MJABJNnLopjUiYjDBqen3ZvcusI+lmOpKUabTRCcKG
pDX+K/XLgILolSeHp6hKgfsVesB/zJCyZrT0n3/FmPswKNP3YkdI+9E3qhUw50NBkA9fvDKZ63sc
LOoo4K9goB89Ll0e4je1mZh7S5IiNBuAFfUYDY9Kuaswf2hKOHraEJCDV3MSC+SDP4a8gVuHJ9um
H+aBQAKInDeQ3ekNbJAuucUQkzv4Qhczq49Xq2DYgaN2YYGeaSR22AleTH3qgEFh8uI9lqiCBjBy
32eAh6kq93WWRYdqGi/E+gAHGz99Nzw5/naNLnOrS915WnB6Ja6L+V7gLlVCLr+ouBPkXgytCgk5
zGxbsjOrGzTQsJh1I8d8rRdvg3xfcxWOcJOvoJkvlG3PDilYocMQfDdr2nBO0qXZr5L876AuR+ZV
IPrtiaWetZ47GxJaN7nEYlFUz2p+7qEuP/93j3ji14F+yRoAMeH/9loGPNayXwX5gW9/AuCHu/Oa
ptKC4XIxhcvcJlNHeq/R8CA7o29gYSinAF5ao8H+KLkgUp1rhSjWFLdiyIdiIR2HSP4Zx/i/69Q4
j3BNIOFUVbZTu6TRlu0AXJgmmSIWHc8ZA++hfPj/dpiD+WZbcZFArZfM7UaJfLuFyQmtopWN7Ro8
OXJ0YUMol46W7NaH7m6+NMOdG4WdIM52aZWzNcVk/7DnO3rqTgJAzFxYGinp53QUqK6Lxj/47M6B
0ZZgTXtWvMRbggOaEOGeO705nJNLUpa95d5QNpB9G2Mhp9TfrE1m1r37SsksIH2Sd/8wrDG4VTjK
NC/7lc3paQUKSaV6z/1pfDUMlGUywb7UHcZTIbTJ35oJylZNkhut1aWhmGJjchm+hZ5MIp8ZfiuX
xLm7LetJ3HOn1KLTXnZ8T24LSMvRLnYmabj2ppslbPzbkm4lrRIKDjmmf9cafgwicKdfWZKZMVww
7LlDUx969R1iOxJiM1Tp1PI6mXmBVEjqczHmct8n0tJ2WyFp23t4Xw9y0cFMM/AIKXquViqFmlG6
nGbod607Ah6lTATG6Br6jsIzyIs37mRCm+4VuEYifaigDIJ16iVxDeiG0ZacevKRyo93qFVVON15
INYXQevynqlX/QrNfpAZicmabXzsFwqk9iVoTR7eFLwkQbd0MjSEuAMDWErgqxLj6OgkTqLAdzpL
vXCttam6cOmUE9Z1VFb4jEnLV1ywJKaIz0UaHWErmG6fY3nWnuYBQlcKjtlNcD/sfv/dQQiJ/YEl
LmD/wq7oaBAyOCjOQTc7qn3VJuTTwxLNCI7cUIYjB5fFk41lxtwlt8KTgo00dZCJ6YKolrgaZR7K
2F1anVFMgn9RdmkCoK/Yz/U2ouk0aAFY/7pDSXb+boun7nLMcFUejwdW3GqfrhqWp82OB2Ui/6SV
sw6DZk87sn0t9Kv3hXVoGxeAXmXvlwttgh6xjmzpdfUsdESEI/LlZcrS5uAM9+aDqGog1bgIOC1l
pXzjM0nKG6DA7TQFym+At2fe6YAGPVqCyBSyJUrZgL6nqU1wizYv0zT4d3R3DsWkYRpFRE7dVOg9
B3z9hiQ+ug7mMZfSxdWuON/3tuWIUtMdZF6DfpCs+ivSRhdgcaWd32WWXET6TsLdIjrvkK/CnyY8
swxSXhcRNr8sz6KUXh+Ahnyct5fUwqmczLcLyZau+wr0WMNoOgMAsVcOK+Q8ZAbNO4vzAGvCdrGT
DIdRjeL3RWjFEyGjGZZMMhFj7AZIspUM5HVZJ/RkVJ4cLhRVqbNVwDKS1dKgmxUltmLT19SCjgs/
OWq8p3+WfFAx5YlE9v2UPzQBpbXKgUxCdEJpCsIfZ3d6wCR4YA4rNHa2PjFR1SNxKFu0fKduZUTF
aHdNOtwLG+Y0rNv0Qyn33UPTlMSCMqmOXBs55UO/e12fgTEesEUjexk1+iDdAaq1Rp4NhhFlakPz
WzUSnmEVcnlr2sJ++5VJIcfWIRoptdoTGV+S9w0jc2+s8/t+CBsoyaAa3rt/M/CHrmpDtNULaijs
G8/tP2Nr2AlAKehSy+RxPGvC2MpxobAxzVrOSxQcwGePxoc7Ett4ptoV+xHI5VIntie5OG/Nb2hd
JBJLA1iiWRc/eGCTiHn0EHuIS305JsPwb5TCS2OKCoeaeVHfx32l3MK1gS55N78gM9DZwtgXWnom
ACswY4OksLtgj3CByw7g1FavTll+JNzFDIFND9trbxaKt0haJXRoU871w7iDyZRfoKIGQ9KqQTm+
CPcWaYUK9a1SLS5MPKkO9oFEidL7VsLxQwQWoq4l2j16vhEYFD4bIDOlv0ZrjVxLxgMO71c0nILF
rqhTkV844rRp/QFaDJutXLGz/UfBZ+L8eOwdn4ptq5+qYJWocEQpAqn6uEOrvS4B7R2aUMGPwqM/
UTtESmXzigZNHGEIuOgY8mzzEZNbWhWVtgu1iiUzZkKEopt6HeEe0w+8WuAU9sZE0PTHgy+0e+oS
98SFJViz5zY/2Kxy/2hjBDrihmIt+6Tgxm2dHsYg/SF3jOhhUdx1UmiA+Y1vhHXklIyNgnZN9z1J
V/34WF3ZcPSre/i7hayf0qARJwFPWP8VVwgxk5uEffLots3o4g1exUzE05PB+Ve9GSjuTxalNchW
7TDbGFNsl0UdUrlfoyNPGXze/xYazu/8UVfQ6OQsVlFp7ix3fcOR/eNQblEEFezzrIFTevwFq5mx
NmbowTHHmGICdMOZ1Up5bnRYzylyZ17GkGyi7FYf/lPhzhBqxPSk7iXS94kdTLKDeOXovfxDGm9A
k3WTi+oak+8HlJzTWHRKqMVZ901Bha6JTdd/C8KYPKuQBMCXhXqcatt5IKug+HxlPxSJ6QA9f8M2
WAjP8pvgtxYivSS5txpSd6A00784kWfkQfPtH2KguKWPGJ6eUvI7XqRd4aq/1nf+C0PXlcI9hbIt
fodbUm7NxoWVaIDnjPZ+jpKLMNTCNp0hCItJcbw4fqA0itiheyyMZ6VkeZk8IAhIPD4ozsg5t/MU
WMZ/AdDIUaBTRMmbQKsko3SiRRRRfxlq2SUqArWU5pplCA9lmY5GqXIW/MtthHzdjE7XHgBIT+rA
UuR7ybEvO8GjMuefbHBK2+OxSo2Za3G0Sq8aU0gRHggvv48tX6ZF3cQFYTKAh3k67FWPq+QE3F3q
JPPSt8eQjGrBLn34LEEZY4/vDG10ekgBlEZKSm7hluns9L+G2QwUEDuNXSTMStqjW7Fddr38InB/
6tKA7RKzc58WZnFlKY1/0WHS+JgpVUPaQ0szS0g3/YtUOnBe0H4y5TFmcGUICxz93R+xWcN7n//K
uWBMyx2TiMKkqgknq9ySJKZtyg7pyzuzT/AjIRVIbbXiOjq0OQDLBJOeY7y5KJVKKaKiSfl5zTY3
zv4nH6EfAuoYFu+yRrya+K7geXcZFi4uj1OGbJ5z8mvW3pJKb/cqqVmW7i5YbnswpCWxMGnVOSHi
Mt59ycJh2AwARpNwbr3FWCDEqL01U/PIydWkwwSXiZ3mEhzrmos46TCUJESbYqiTZEs5I2EmeTvk
XMuOeq1CgKhXol4yc5OO/QXnJIpf9zxOClD7IvUwysOg2DaXO7JjfmSPUEkJOqK4JhK5fp/bPAeQ
6kIgw5L7bBLY2zI6RPamKqEjl6Q84bIV3v6aoREYiac+SIOqlCJys+cUV7GtUSOEFCkU2MbjjAP/
QEHVvVVuFQDRmbm2RPPCmIFCya0r9kB17PaJxmMUfq2bn76v+4qXnxhbuDl4W3pJ0Fxyc4P6tRQH
0oQ8Ji5/x4tFMai1nHUjqrt/BvG5t7y12R2PWvXTlcEQ7pLoz/52G0zZ1AqU7qFqdQEtxxpsCWbZ
XpvJtwtWRElkbgL6k+7wMvm6Ow164DoSAZm1ABfRJvyTnUxY3nvDZ8HmcGFF88LCYVJ4Mk9NyXhO
IsUIEmepD1d/XXT6Kk5IHYfLEC3BC8NWIXFC2SFRpWiqNGTcSr0A8Enc7dE7FKBw2OjdtBAu2tDc
gVVuAju9nOIM7IDr+SYJXw13Km1/ikvHwBJ+dX7+B49El+zfzVIlq4N6BlL2HTI4WKrXkbTGz0AO
NC9Y7p35d3Wfuqtc0WoxJMmtd3UGtcdQw7muDwWkWof17wvLLKowbWFQng+ilWx4VVtbRN8y7ofE
q+wXxbqy9PvFg+g9evuXLp89S1ORKEdz0XPhnFAOmltBcs+AHUE2p7/LKUl7JxU0beb211wrrGe9
k3YI1PW8itSLrBAIKJQbbo0BEox0Da7gQBsmZdZ8v2UVnCvylW6tos0cr5ugxykv/VEdak7wd3t8
SC48yof4S41J8GwIHsAckPZ5ZizOMWH/p2HQxG8EeeykjvYXIxYO0m9ZmRfAGYmYLCcN/ZyNwHOT
58+/Jy+5jfJiI5bWqPs4ofPhw45/8n10r3csykBYfbdvwWz3CbLmmDv1QItOfvmhBx/UWQzsSWnS
1FOtWUJdK7CsPxwMkbMBLFe+l2f9DOvQnqk19yuLXOV+Orh74lNMX4YkWSEFSM8s/iUoKqyKLghd
B5660i7UmvnNIxjnNjfWt7U15iHu7bIlMIBwY35jf/ww4JL1vOiLnDfMERw4xWC8URIaVxX7a8d9
oflOxPvQRcZnpME6iEHI1dLgrGh+vi2uxCzWzQYNI8Zm1oCRgUBrPkul9dAGI4afiuuf/+NKVgZ3
sjnv0SVbnFKyUPmCsPVPYcLK1Y+HBiEFm15qMc8PyK4uA+j9wPWfYEnIKO/2zpSAL1sWOw1FuJKR
7s+FsSbfM5epraxrsHVcw5TPp7S6Cqp8O+Bf9s2ee/n5OOAznWtTt9OhUNg8uTYnWSOkBfJmfsGj
OM7FBsUYyYui9VGKwNgYt9IHd5nvDT//r4rXEjGXA1jnGg1STjjPQRpmszDhiPOHG1Z8Ql4+7EKa
ib4Ale+5MNdQM1ay0GDBQIb3PY1fuTGtyB73LlIz2UNrDg/phKu2+eipQsvxgVPN6pUa4ZyMIvJL
C3z9z05J3kboIGhvPlY8Ie2M/74iAspLo21D0K5lGZ8Feull285E2H96fwiNL6EapooxgwjgDNgs
t0nb+Eca901hqCpNMuC8cVaPG6Qy6Gmg7nHqviD+6EI6nF+2SIaxf8iIjkjAYQymrIgl3Mv57zxE
OWA8NJ2hZpN9437uChEEoeh5CoVrbGWDiQcBdHHIhjIlzlzMAE1EzPEl5ppyLdbXDpG5KAtAWvh9
i6yRqPFHcar0hoiQoa6jRXcvEHaqiBBZ4baEqUaJv669KZTVloZEkVzw4wC7p3jIDt/ThKz3ssWS
Sw5KarjnuOyd4tGqQKxD0+HP+OkYtRyL9sw06FKQ52riFBqGfYneHKsNldWVgzDpWSvwc4VKgVe7
JFMYa2Ea1NN3SOVix9pmJlkfNySCXDQIs99YnIn2si4CWb8CD2IA7YX12hch09KnysLRHqbrgqny
2zJ6uUTS9fTSZCvQFjhFNMZUUwZ0iQjAdLM9HIF+CAoBDAVci90zIagWldS+gm8r3TYXaGDtPCOD
DD/I8lXDXcS7GdYdgj8eIYacKfzBQ1jciChepVgger+Kq/o+yzjhCSrpDxZ4LhfBw8pLyaCoJCY9
2eMHyazIIBthdWgDZll0WK4jJ+9ZXgqEWyXp2QZLidv6zkMuZJskobvPrhvUltuXO0ZcXHXTzSz4
dgipkBGBcaAxivdIA29i7EkX0CmDaQIS+TlAjhusjiXTSw46ytUvuoEL4C6WLGUO0fZhQ3aywKRm
Tm0A61LUFlfbBgH/RFQFGE9VaQpb5JLhqskg8s8FcYdVyNaqbJICw1cTPDVXoGNpTUjgWhKhHPMv
EVT/B//7ifqQq8kswJ98E0FgVwXWp9laildbT8gibFfUUy7Up0QT/jqScrRrJX/d1VClbx5XGU1i
24dOP+k29xCMcWtt6IYzFm0kl8SQ3C56RvjO/5a/9Y+TrK09n2oq0UURVCaKna91os4T3vOT57ud
ttEZIEYQs8zWMpWX9m5z3j+sWJwCOn7G46jOhY1Q8x58owRKK403zzHgUlZK6bgt41zECcJZwAf8
+hTDsW4cDgRTMmLOVv4jDgfkNU19+tc1U096aK8nHgfCs6/8zle151RPZi2cOHvNXnHqSDKgTvLy
6nVIaWkxpr8I1Mfdw1fHsHa9M90rgjRRiZtJGMftUA0Fi3GwGK5cV38xoLRyEM+GYqdVfGgAEFS6
T6FmrRlSmFb+wiDLo70QcUm+15RS2wUl7dvwYMbebA60rgLc2hfsJ9FSTYtnh7CZPwVj1TIt26p3
X8iWICwHIgaT9x9iE8pvCxH7alhvq3vjK4GmvgJ9HUmRPxuNfB38GocI7B3z2r0RXTYvFVKga/eO
V5GadQwGh1bo3h9KmbwB7yhh4l5U024ujHb1/YY29ub/TVAJjf+o9J/QxEyyI+bHNt4DAfITshMy
iT3gjJ3K2EGFrhQvCw9DtU/YJAjgwq0nJH0VK2HbmQLg1bBmJQH1arcl5Eq2f6+hq6UOfhGj9gic
B/MLRshrstWd2AqIaU7is4kDe8hqOLGdvKAGl/sd6ppCtXEGTFwc3drEIOZTEOcciJ7CDV4QYxbX
Crl0fwF3cuVGwPPT1RqDE14Rc5MzCN0voTvkdlRPTkSNvhq/31O/jyPbbonT473/UsnMng8Z38C6
NkPP7A6qkrba4ypfaUcz5k9KzD7EYOzv0li1bT2CpKgwtk/hpfygN0vPaWdt85KymZ62FbyfELLJ
LDi3ZrokzErmhi2fxRoFBxxryO4jJam8Wl00nl6L3fs96nKVtToju0sfb5BvIYK5hIAqnHOJFaOI
RHk1iNGYJSN6Cf6UO/N4hQ2V0GumQO5z7O4DXncwpWfAK5ql8T6J+Qs+t/f91zeXeFK7ScxudoHZ
+sDSCgy3R8fmGPljL/Epn4n8Y4eXXxivH9jMv/iRf/3MCoLLy3i7EOoLdZlWysKLab5PAkLisSDW
vLCu4EPbNoXrMxXLljT/qcFPBbLRTE7G4JaY1dTlPPDpOz/sKNCqd90tyskm5YG0kXQNNDUd/7tV
7n8hIWmh9PUhoMaIFjsZUNJrqrQJ3Zad1xaSmDUxTFjpyfy/RTqth7JZaaovO+fAVId3D2twhw28
lnCOvJNa3s9AIgXstJ3JXINELP/l/IwF7eFoppsGnZwaaIzruuaJu4ckSSnUWGkbODS+1byE/usR
5dXl1WQmCPORGfpIUkGlFN99qhrqoKFl+H1lXJhjsyA1D/E2JU+/T5ZkuUdoJxxq1NPT9EBjfrV1
57rmJtLdnHzAkokK39GHmCjHB+UXOBT6HdaRVekU6Y898oCUsMkmVRIp/AmlYT+1dmUeoWyFkRPO
lppe7UiLaSkJOd1VvS1OUovtcRceFamJiIejDMHTapjQYHYvkevuuEG+iNNdciflFJeM0F9mBHgm
wJ/9vFgvqrfaNCRS9Q9YbCrbfR46SaUuE7zVlf2vNLu6baXlLBl5tdTcq4HSbrmKnSSJb1i/onRu
8XHIixpHoeqYoewi8IFmGac3NUc6HneQcmWwMC72k6a+mKx036KBDR8z/Wbu1Rvt83gQJKwipMAh
GxBgIcpxXEcNZKn6HqWC1ssIAWg1/kEbLHrizHH+qPX2Q9wMW75p15Xkr7cN1SNwbYNbC9kfVwJA
E5JE7GS3HasVfBvlxu3LcFUDxS0Ww9I/1g8TsLvv52JlEsUlj1FjLr26kWfeiCKYqJp0pOEbia50
Fyv5Qjiojy0XfPQMujTTrW23w93asTH30nZJ2AxF+fj/3obWZZyLpfRG/UOhf6gfKIQIAgd6tLld
Un1aDQIAUIh0t3kgHLQrDIItyGueDTy8jc8rXcqKO/O+KbM9coEtv4nb8CTtjqFxcsLT0pSPz6DE
Zo/z+CVXvRQWHmQ95lfmxTDYfPFQydvA9j/bUS9Y5Qh3doxXzxOWejBjxSOc5WE/XCDPiJtBJuOn
yshDakmhug8SWK/Jm57i1id8pqDHqR8oKyWOs3Fxw9e/eo8SljR3JZ3XYiyRQ3ufwiCJHvizOCoJ
Xit0PVKqRFmO2HIcIY7i1JvSbYh535i+2gh7HU9EAu7hMYYPm+x9nyzGzNNoe9VUCGqDa1KsLCWd
nB9es9jCvNjOLpguoQUxSVu3yWKJ7rR0Z5G8b8GXXk2qt7Umot3cEYHO/bRSichpOT06CKwvnxVy
xhTqWVWz+4NbYGuD786Cu6ChVst2Y6/KcVb93DdMHbC5THCEykW9kaCBBP8QjkI4DSLnmWyszJDl
6Zmc3q4JmwkOCTDa+hKNpMPNVxgjCOo2hn3jXBWAfqW5KHeUlXc/YkPr13S5Cp3YASERocxb+Jus
+aoWtLPSreWqGf0PCasNouTSJhg3gyV9Sf8dVvDm0nVlW3ZkmVtAW2h8aUXC97np54tSsP7qOwfz
vSShd+yDL2ujkPbFf2w6Bky70VnFO/mgYeiTtPLB5ZplhpgaBoawWStjM1XOHz2TWDjHN6owQfgt
+nNa9I5RJ6rGpyCzQAtXjaUwLiSKNJrBRDWIeA82X3UKaFuoIF8abXXIUkh/QOMJ58TLPGKtfds4
Osn3HTGB5Shx4fvUizM160lvzKj9w2imvF2z5UTYJPT81+QQFH2MhniDDKNLxeshkVql2VjwFfRb
34eRkeAp+P3F82tHKQ0uprk5+gPn32ul1ZtkUdz6l5f/xcgtwon7uurrSSbOFh2uqETJky5K0YbV
mxOWamsiaXmJg7zd9ssUOnZZ2j22oNX/M+OydoUMip0LXoNInZOQIr5fDQPO4bBEj4CURPiMhjV5
W83ZF6kWGJvHsuS38p4fAJUTYNPsXtR2b+s7PrKd3q+po9w/a7OwB/HtJIPBB99m7aNA4qRuWroW
4KBo4rwHMTbMzk9ohDSGvQbVS29jUaQUKAvRlE4kv8GOFRmD2NBQoECRaW1q4Riz8yWhBKh2F3pQ
xm7qhrMh8CUi7NBs5xmdG3jb6bIhwpEnR4VeRFnWdSRVNQxU8MhGUHFgJEOJeFUUkiX/ZbxtYAnI
hisW7rQ236UE5tsZ9fsF/I2mErxzR08daqN/jDHZfSAAVl8hVO+3RlldPCf2dP33WgJ86ZGSIxA+
tZIj83REBaUAcQvO5/ewlAcfX2oW2Ry/9GlYyFJfMLoV+R9joukXaLRyCUMExLkuTyKrkqbTc0dv
wdoZUxyruycRTgtlBbtbnLoLy3uD0WTh/dFV/2winHHLs8z+GtLTLvu4Pplm1pbUmUQhkqQUapUz
GnWY3TUOOJJ147Yxb5JrTBnr47qosP8srBrBJhTFOvf+VFKHpCzRP8G0NRIpJ0/meavAEfEuMZEm
b438D+Et4zGPyKiDAcMd6kNvVHt8E2Rw4eeSBbXqRqnERCwsGtlT3SYZbRUiCo0fLXwmWk6Hsd9n
zOFUledXyPBxpzOLOG3gqJ9sEad0OFVZO0sDbzJ0Lc75G9LZQywinVLZW+/jQBlw5TmEcSTWR/Nz
cuDSU/tXpZWITF21Cq5/reQJgP6YyFKyNeMeuXl5zjRCltkmLUZk/iFxKUQ/aMZ2YqjjZstd84RL
3Ef4zHRof0lew453dtbEJRiVc2dwyOk7rRJL3GSr+JcchM9lHQuUIsIrva2/PM2e9lf8ohQyzCkH
FKlvkbkLXP7/KASvY32Jzq3mJ+NC0sPiOPQhAB7T26+MSshJYAHavMQ2TM1Dj+owOll1Z3+TI+Kj
Au9GfarjR/fqwkxTBNtd71pAsb4abLH+S5r4pLD1AW0EEKkusI4M1JnXfKjmFBd04vI4DYNe0cci
oHrm1lxABQvlpJEMPYwzygBW6XHZTiwW7VedowydPsZ5ebO/0HSlM1L/W/9YRNn+CB0xLZMk9RPN
pFlAav21YkO+tQOFcloXpR/s4iFgT53QLm4wvuPh8iu9ZfxKn4hDcrVg3i5v1CqWMgkpjxpKA3/m
M8pmbZNPsEU3XPaiDi8LTIn88ihE6zzbTsbfMCJDaMtrdU6srg8WbSEgjzvf7g/8pw+qiBfr9xLR
TPWvex2bTckgXyApYEQ0le/D7L+aVfCk/RQJoazLPuVTq0oohr0IbvGP9YwL6rwXLum2iHL+jQ7Q
Uu/dgU6TWKgS+JTnrIYE4zM3S7F8NoOJQFhn7+yvuDBlsTCEOkvFF6a6MxOLmW1kDE8OrZ919uzB
QiHAl+e7BiR4QXyZ/5YIHIBHEK+KPJ7YzmWE5VUSuh7adIP6yyIVGVdYvKc7WYjKhCIrsJ0tViFY
nu16vGuF+9s2X8hhCOJZfIIvoh/BmPkOjF5kPJ1o19/uUPRRdZXV5XyjOJL7T72OmEdHfEhzbwjS
8aWmz9iwHIvBSDvTLWa6O4GpZ/DiG9NIgUUTSyhzFzElshBkjnAS0lF9r48fsDm+sK2P6gJjONGE
lL7Gd0FIyZB7XNH8awf75F/yroQRurNavTHYFkz48XHZpT/x3o19tx/PhYTPEQWT8yhhZXvta/Zt
MjsRZqMACiTSAX8vl3Cfru0bOEPDCBoCMWoYpoVuabqXQixsUbB5dJ92ywj7BC5+NJlG7jLRELfN
vQl3jEgYWCt/oAfe5sb6PI8d750ChefxLNo/6ha15LsTBYvvTIcTDlZ6hCNY53KAtSW1aLl8mnLP
pcooliFUoFTafu05q4ti0bEZmaMV0YGcwUeWvlIUpGlBxJwL8pAEefXdg/gCvbO2upW2qL3tc8SF
IYgenL3Li58KnBkitmqdmTPQYlJpIc0CQ9iiiA4EDgy/QnmABzikjpDUG9NgFn963j9SyPzUME4F
ZszMkONgB1+wgVwVGX1o9eE+ynGK1zfzkFFcYVn8yD42m0olwyR7sgAtx3c39Law4+TYYllkAYYU
sL8AL35AOY4Ox02mDjwtpw13gK7hbX6OFEb6YQj6WrjDmFFz2fSn82ApI40LsEgxa0zJt6QDsXkw
aykpbny7N5tlhLs5NoSBReeI2B5Lb0wiDa8xjsPkyk+llQxr/wkNT2giJIyf3+88daMS1/H3Jt+i
hzX2gpEM3JuTjftHisoBl+2aWL6G9SEqu7+MdhIDBSi9zLOZMq90t3a4ejuOT1SaFQjyrqGARTAf
fAkMp4gCCftTv8BCJFcofExTSyT1ul4fhKAhRnI/qCS4d728Or6YCFSUBmJcJ/rDP+OJD0IV09XI
efEIdaG4Z6jgAqLW2G4kTCgBtHnvx6iW7kT2TQNZhpBMayFyFdlcODDNM/ompNGk9IWMoDCd8U21
VHfoGzL2XvnHldqVCNNiT1ReS/uet77UDNefPLgCwu6zvN9gQgveURiqIKBuRpYSPTanh9ENjfRV
EmrSTAFlruS7MCDBazkFtGf/bF5kep/lCBe9YKo+Hw3WxNX5sO8RGX+Mhh84KOW1HJdpzcJsvbfg
Rlf0znE29B0/uBCqCzF59xcoart18yWVvU8L+X583avj5iGVEVrfNSPaZgtfMVf7DM7Nad8EyHtv
9QKkByaXYzFbGlh+IsUOPR3mmFgpsBUNRK0x7r3Rs6bpgcKgJA3Ri9O4epNA7IaE+pcgomLYrxgM
QHlTa0xgBekoSSQfCRPiv7JMxTRidIQ8IdIm+ljgaEU4dlF6daIDer98sBXfdEnRJM3VDrckv9wu
/TCT17yZE+2pkGTwEiLjzCVTl8CtW6Q1WYk7oxx6w/Eq9imak6LERt+68UtH8DB5A1dfpE0DxRSH
YDqzn0HjALFZCY2KWrrgXjxkf6IQ6hDZ7Pm3bjexaLAZVQVvQXISFCBv9qp3NmfnPP4W0yZDcX7K
wtmN4ltvz23TitqAS2x9cURY3SSR4Fu3jxviDQxJ5cr6DgaBamx/CuYBokrGNFPVx0AwihkW7DaD
H2KVDQYu2t/ksMWtaZzXfdDzIuWaiOZJX/9BZUDxNZPUoGLP4lNIvYWmOorcsL/iKA6NbqC0hXn7
0/2LrMGUQmtdtXMgzQHLAIvMzcZwK+cFoe+wAjk41ROyk9MR0s0dEvGpJk7i32EEWH2dvrLD5Ydh
xLgp45G1/Nek6J9B9JyTl88Nj12yrR6/uTxGeCxh8PIQyG2Am4XmIp0iviXf4bXc6Uk4CMW1BTKE
DXuWqsrEBLFjdVHO+HVeUJsdIa26mlW6OumOM275VvUCps0BoN6cWhsLsrrALnXYlwR9rSu4v/jT
24tGwwlcjskazFLQ2QrZ2afwJlERrlwj+7xT/AIBjYPldAe1+InkbEGo6izwgSbfQv3sA9+CjhLf
I81Hr1q8XckSveCISy9bgBa9nobCkuFY4Hs9lmMwjvyyxYi0kPd6g0Pb0vMwgccMzXUkmaRtXLvC
1EmRYGlLfcF/r/HhN65kxS0Fg8peSZQCrDz+K6VyZBVm9ju1bRMLKtiq9yP7+HRSugRBiMeIpZNg
qUO6Mz2gm0gYlcBgzpCts694QRUl7Fe61GxcrNrTPIlPrAceqWrzsLDDyoxGfXQsNZa2EvGZNczn
WyVuucbk5wekZY6C4674yg7i2W49SNSWeUra0nXCQh/nNeP8EC1tJJHmGk5fJI7D+Ate/DW1TKyK
2TMWLmgGbAYVBN+dPAEzuLv1E6rQogux9w2BOm3BLqWRR7sdAe6FCiNaXoCqYN0xPPmmtigdy/VV
3X6zGRrNtWiljvAE4+R+Y8V23P/vpjY9V+htBALbAtKxJW5sLrHwPqfqYWEr7KQL2rBPHflSGkXP
ROcRb2GdJB+fK+yoATHQ04o1UPK4BmgFtGYAZeuOmOkByw8HSKnyc86/JWd7yyNCZaxtc3Tw+PZJ
CyD0C5E3pgjEkrPrmuKeWTC6DJKhcbPNrx+AXflfoIf7WlNjEpB4FWTnGxkWMYYzK3y1BICmADRv
5+n4CrKOIkWlWWZNJCMQgU59rzMvl3LO6lMMGG7wmteeBpKCvvXkjyEW4cKDlrRot8X2ouPYWqAT
2mP5UzLs/kQ/M91H4x1Hxl1yPS/K0HjKqbzXKsIj83zpr679sIp8Roz3mnZOhTXYslPOg37DKZJd
BNy4dte0mIPeWLEzTI0TMMRZMtv6eIdU/ezQis+HVaAhgqB5XAuN9NIonyA3DI5JNu7KM8ZZo5wY
aOM7YtV7oAa41odhD9uzoBtkIy38wTbmwTYv8awxbqKW6ZM6xeLp/ST3lOulYkfr1zeibWoU2tYs
Ru1Rw2oEwjfqeK/SEC6BnXCrU3TSmdTZkVwzYbB65gyso3NqiOmcSCyS1qCY9ULE1SFEXZdN4vu/
AxguqUqxYb2vTiw3HnYN1kZcttNmHfbTWs28CnMYp6KxYDWkW0rzEJKXPG4+NYRv0Wbg2H/Q890z
XGfQYQCx1w6wpaO13frTqjPvYle7o2q2bDU/o6rM7t74jRmQno14qYf0C2BXRgDHPZkPrx5BUOKp
QgBDxb4j7fIr1cOnbzL0px9Te3/2k/ZNLa+a71k9q/978ESbYEospr96YyD+GB2ogWAe+wjGQ3wg
XC+9EQRcvG0GYxz6dgnXt5V7LpaEvKsehhJvNTVhCKyJ36kbU3ckaUxV6LBl6WAdDnyipZesMl/E
qlGr7c5z4gHuEV3daT1C7Y3ECAsOiyIjIg+7GkuXmlw4qFfyY+shlftxQJuitnpQtkZQZ9YXM8oc
VH05gwrZZc318zv7Ifg3SfYf9QvENZyp0fy99ElvlWZ7nRcVAMVVTn8rkwtBKhNXHQt+CII/CoTc
k4qIUpfvaGy3EcHMprz7yrtr++JdMtzm/cwW/ktHar+5UghHy/ooR4XEHP054kN3DsItvEjz9QKc
/yu2WxWllWy/uPrBuJ6d9kNOq19PkLov6jmM0sYPvuxkVze3bSbMIpojHOHiXSC/ogi1U4aktNB3
vRvRtD8v5Modhqk8wIhvRWeQyTIfQqQacjzQj4AfxoVw5zTNxjSbzQx46cRwJ6f1Zvc5Nxe1SFyh
04fM6j7keM7h1Yg/J1V+Ldh1GYPgpMZsZh7THukdfDSn3v3vvK1zb7hyDFU4ftcsRaU4KfCPcfgq
/8fxLdSkhLyigFzciZXJ9oFkbJLpAKMRml+lYOaUyD/eZZNUdmOE8dnmjgL4ln6ElSXGCX8bxOz2
KJaE4TnMR8Tq46Bf8+/3HFK8SmWCsXVQXBr1j6oaPsHPL8kflL35Y/Q1cm8QspY9j/H95kLSwuKe
jNv3PGP6LG37pi6DuWoKXj3EDHWFI0OijLH1L3ofzwFzj+zM0nt0fYI6+vjw7UoPQgIGOhm4Y0B7
qqAysX0qqcqOCn42VBSk42cd8CoeBQHuSok+5yYbBH19OO4DCkNsplow75Gj6EBeB2ztGwh/6RLY
kG0uTJnTXf3cYGrH4PsJ0PgB+IhPJ2GS9qVfd2q0CO73ZESMKCNO6nx8JICG6bpbowQEs9KNQsTi
Bv9ssg9yhAimdYjmLHmae4y0qogT7SrdaX9HWpj9GsV81poig9z1afDQcVBI4cfcQGhcPTQ+BX3B
mhM1xC8RinToYj4j70qXxXSIZFpunvbQVAczNZsi6jGSEEJ4zVZKNORCkA7uoZiCPI36u5wvgeid
JSEJYQirxQQvE9UDVCJ96RRxnNiHIwXkhyQ4l03DGzZBBWpzu8ZB9Sigyr6bAvxjacMhHhPqhNZM
0CXB6lxeRwJWbJtmjkkclynamqTUqS6mFvbHSo2uxOlK223ZDyqvXMoKD2WE/LrKZeV6DiVPGCh7
dDe9riNGn6uhVOhJpwefZ8E6aEPUTXKOgm/8TsD6lDGRXIOXJm6rydd2Ojdt8GI1NTBVCELfMZmt
xspRTPm4u6SS0U/VcWVqWgdfDpR5gRnNIwsimq/jqqmPq97AmSIhY1xz96nhUbfTXDD2U2DXxdB/
yOamWO3FECsfmZ4fguC42jtWmd+KsXg+O8+9YlUgq1ayBAKvkCtaN6BMNZn0kw4TLkTW/JDV7BcN
ZSqmBzZPQjoSGEdkcz6kyaRdu/aLWEzlDIHyw2kHKdTxM1S7mTufwnyQccCcPtDV4/6lPkKTIFf2
T+l5J6xHude+AWhUN4uqe6H3H20Kq5RCrwIJiqHjMlDiLVwHNIRQ9cOPIIo9tgKCbU3Fwg8k0Fay
JfL8iGURfWg0w2zQ8WqJTufznGZyxuC01LZlVmentElufXlDC7tWrINL+5K3NZY+Ga11O+LrbTk7
2r8ahc5J9CqsnSXcoeoR1i1AfYPtadbjUQwu8e5sQd1I98BJyuF0f/bmN0Fh7R0DDhOrjuUOTOwg
af6al9+y/o8qYA9UOZmqAf3ebqoIPN9boNqS3DRmoot6bpK38UQRUYNj8Ehi/kzY+rMCl5uUbyKa
w9UB4jZodPLm9qgh/PYKtCbu6WHdBHEWTfNGZu0Chwnip+NG4ez+5PpBO9JuMnMt2uGoBdMaVDf5
KIXLgTw81OTH5VqwaFwZiCgd+PHgsTpGpsaGhOnAzVds45ETYcwrTO056Azmk0QILtpJN+ovsSs8
Dnvuutgw3KsQDmqfD4vtPoXpxxDbhPLU+YMcNGheYlrcxgclp3V7wh63vnmEGGGI/86NhttmrYTP
HOJ/UANcfMDhHB/w1/czYbMLhN1EGhO3zmhe9y+/A5qmBSdBCz4uZvMa4a1JVp1Ia3/mVEcXA8zo
wDIE8CgvnSkZdxDck6Qy50NqCXNeZvH+wkFFEW9P0xT3gT32P0tNlhkZnHNVOi050tnIfrhsS0H3
STC8C8nSVTlBj/zc5bfpRE4z5RMsvl7/TzORfcEiz/tpKIRdqyMYDvIfA2ByBVTowDcoYVQQweMi
xlhap/cm5cukWZJI5qoN/rEBIEg8tHkMauJ17VvQimw3cPOCjE1WwyiboNEuoRQ5Z6GSrrfxWp0l
KRRdCr3WQcxRspZBl6N6+hmttZe9eoB8CQC/dfTm6+yHb9yE6pFC2Gask/UJbN7XfgfOc7O+pZZ5
Q1zuUfCcunR1mTKdJSW5tqAyGoq+iKzg+ojBtiJDPIH3jbted5FsRAykDxf+Ha4brDld3CvW/BIm
M8NmYxhDx42UnVrCuPNAkCuEwVKJr47RVdHFUvhgbDo63o8rW/feDKh6tUsNHynCHDnSLwvoufbn
GrTWxbvcb73XgX16YZvtLPnkP2hFjlfRGdL8H1DLWBW44/cIG5ZCWhQTpDqHth6MidtyvEyD+g2O
N/pT/LWkuOiyDQ5OUqn9QepGPtpOBaWpp3cZu86torAkkFLFxJoYi1HKnFWF5fRqE+wT4psfoQHR
CbkMEXl+wN+ye9U9V/17oZvHEyj6hdbtHVv58rrdLvwjlxwHzaI9gsVZ/8KJszMkniIQischZe5T
SMA1/8MtSogrDKBo9lDPALBCYKrqoAWQU4nLfGImpdPIkt5EcIp8IubZq5kRfTN+KQXynIyYWati
sqGeBClnqXVdc5SQX3DdDsWhbJUsQFvYDBSMXQu8ApD/DoDO/JW/YIZ32QemrDEoAdy3HXWxQkjx
cdUD6VOxwoJqjfzXF2810Xf2vE7FUbbvt49q7Ozau5U9KZ5rZ7C2C2tfIRn2yBk/v0+eAltAiq4x
eEu9DHYeYVW7dUUDMEI3JCDsssxCNANJJVihD1ihwzwwH3OCPShTn8qzpASHhbfqQT4cRpXX0ssy
rm1xP5SgMIVmVcpXwMxpQTPk0I/P64q15iPBaXZZgAd/dbROmpqoRGJsdqZNL/6dY8x08+UynXUF
AF8gyzhA9JFnR6Dy6rBUGzd5ZcDZw8j+y1dyF3oCP8WR6ue9C4D15TxFPUyqarx7xzrwsc9R0HYP
2Cm/n8ayy4wFC6ItExA1/qitndTWGGtOlo4B3N8Lr6jwjgSfNa7CZo5xYeGMZhw4ZAkk6JmI/8I7
E3IiMv7MVAt9MtsSe9RuHXvgQHzTsTVB6s6eiE+gt/2x7NdC7ocvDrlaMLAC3l+OPv+xI7kp4hKq
s9vEDYduFkMTvl0ttZIPaMhj5XsImOJmptf1LNszlqtcQoiIPJgC1b0DHAkP0i1xV59FA0zrxIka
STCDl+2XQL0e1u7X2fEbFwUdKgWa4yNKutuNdNW4lWFMv13XWh1Gj/kJio05guIlKw3GkzvydSlf
TFOHMLpkf919dZyjvEsP+T3ahx8lnOGKjKg/oMiM3uM4CWnKo7L2Mlh5R0PlOH6g5ueTHTXO5RGd
WcskKGWE931Zu+Wt7Xz3vUsYJQjiJiY6xLmXSsYSdUV5Gn22MtZu64rzcOrCFFPz1khtmo21ooET
EwpI6oCCqDGyrb4nEAWI92BWocqlUtnrJNeKpi4SzPYh2CDqUDZuW5znDhRL63u0WtqRrpwC+kQw
0NT4anq+1SDUPxmf3bgE01Ttr+0Y7BBzA4wXQmxZ/C4q+qiH/wq/6qm5DfOg7J2qnenECLVH2PMq
p4ozd7N0fEkt8qArC4UvBurrdQFyriIv/nxsVOBjuvlAs90gDVRn6HA8eqZhrtcrC8ufIHbBEqL9
pg+IiY/lGx6ggqu0AP+EtiY/ag56XBJmN9AJBQOBWnPspoQWEjITijp9444I16H82/x76/MwsU0V
4fn4nFIWy8TRh+O4uRu4/7FOpSoKol5UyaPlC0VrMOkpgDISIc/7v2LLgPfz4z8QUx0UfnJkRinr
DBj+BX3lL2/RKD/lMLz/od5KqaIa7UsiZxrj2uIUka+DLbwVqjFyGYI5/iR9U+rK/ZYgW9yQqBee
LsNfFFJ8pfEY05lTfhmM7jSImHslSilv+jXQFXis0SoSVbT0BWCcwZnzhp9GE/3mUte3fThK5CkF
b8UnFiO3Vjg+BF1CBo1XKTfn0iz91ICHf2tm6/Tv2YPddT4n6OxIJFwY9uyz7KfOQzgi2SNsJj6h
VdVSum3HG/VTXYtDyvmQGc2OyzUGQLKR9rbfNbFEm9mTVTXbQr0HYlh6aTffc9F0Qe9Rso0d0UtG
o/XCe2o9cis1nU0JuTMvO6j9CUXszONj76dE/TDuv91yh0c4AvLOy9gevdw5Y6TSXgWd67b3qWX8
4G1Sm++mjxHyvD/45ijlhGR5xWSlQJJq9yXLtJ24N0xIXd5fW2XtVF/dFk4wYDbDn97Mo88GLSEH
h92+82gvVm7GATByVjBwR9vzj3+GWUx9CvUeRfZ9pATL/4Q+UeWjFYg+eaS81T/sivI5GPnvcXos
mEGyIw5TlbhTiL1h9Fz4CTBm8Bfw3rXr3LEBhE/K7SSOv32gdKadDeXgfUTm6ClUrSL0mDBWNda/
PWLzITFpGaq1vaFvkarWS8UhS+JVMkxaRh+FtMyScls7yTV0d/j1O13ISFFfiPTxyi9gWeBVkcAe
Nih/jSTatwJcGPUQLD2eR/YWQ7U95WryJvQ+ri9g4hxj65jmdMHXa0RNM5dFioH2pw5sctinYzM1
ROKgvteq5cCt5wLDcvrAY0veD8omiDSor8pCp8PMUgJBsVed4NVJPAMEf0e8XoQ0twLrSALKTblR
7hvNg0cbpIuvn/ytlGJyj+3a5eHQ0QNxwiUXf7nqhMq/5kGp0LaM3y8Q+qgPN0PGk9VPjFuz3SxP
O3mRcJWyb9NtnwxTYykSC3hMwL7Diia6hYGqbabexieJXD1Oqr3yHIYdGz0MyxT+a/0wSbCythV/
ufc4mJjSKh9/uErYvt9LfJnZ1k8oHPJJp3KuZCvR/dw+tQNlVQSrdopbu35TVQzdcuVD7BYHc5LF
ml92qwDnXAoPNYsjoSQWru4KRQYKE2hxzc+dNm3fMMB5CMiXwDVKZ5/n6LtCKycMkbSpHObVTpsP
gzHmdWPLopGoxoHBzaoDgGSaPfrvnDuPWC1TeUjDrl/hAhwFgyoZJjfHPv9R6mV0wt8ttI/12IJV
q/8I9QUovqyl/8A6JtCbvbvPlxJJiuawgLH8UGhL2LLQrogJC7HgYX3ReWevZIuUIHHuF+at3pjJ
zF9kilHVQwqbloZ5BL5pD8T4mvPUqCgADBaI4UNJZJ2ITRKCTf55jdBZnEP6HP1TzJ24Dbkx0WF8
ZyTpybfA0g+pNABqwyuF24WnD4QOPWGhmAtWnlnivFM7mGOhjZk6Xi2qY5gFY/vkCouYhIwZP5XW
4ctQw37yXRypXgXKvd8TIwyFj4uigxd/kItlZ1+eK667QuIYABK2wW//dOpkOvYUitn/BzHXfW6s
SKs8qsOnIgyauLnTrCAOFK/SKt+dZZcfyrhEHIWwx+5fkltI6czL1LVanGAD6XttKgjdiU3dH7Gx
DktXWLkuA8BPKfncnZlFBAJQ1pfsiT74DTC9EuhVChqWjzVzIpz8HlyhpSPrnlfpnlKEpUvjiL0B
j57tXI5cxqi6cFE89iK1P90kR6UVmdgj4l/JuJ93vnZRWDqdSPJsFxNLulscwlp2h3AnLEUig3e1
ntexoJat0SN2dpVkWe1xn0gQ01sZ9OiYgDepbVW4aswV70kc1YXzYNcEIC3ZCTEzD5ukUNzymNJq
IKDrTmnLa7+mM54cVblzhokuKrWvlIwIpu6hPTqE0+wBRbi/IBpz4/S231ncVn0sEoWG/qkC37Nb
R1IERRfnVcwd87abjGL0emzrhkViUB7JAJqOQs6R81rOVXtB/sf7XBCDKm7k7z2yn+WkK7HD2Hd0
py6agFE+C2X3pk+xhmRcwU/4+Hj/H+qnkmtKunaRxnTCOqAyoBe8v65UNcnP1RHbZOm7IsJIqyj8
uBFDoin42zOn77MYcixaPgknD0dy48gX7wK7YWdzpRQNnE++DywsGQdYD029XOi6TaXQhj66x8cY
kufLbGtTHenfx93Yj/MyyM6CoPbXgM/qg2KJ4wO1jnQZu4ncDQLEB8EZ3vHNxfASU/qloOVciVea
oTzWt7nwR2B1kSCfSv0z6mIUKZWEudQbxE4Xug1vkuXM+XIR8d60Fol0KJDpLd3hwTomW7D+izSm
BG5WxPhQAdAignDYVW+Wxn4cEgKH/Hd9S5dr6CjZEtm0DsfQZDPU9MVnPGs9WpBX9FVzfCfVpbG/
yPTP9kD7EjuzFLurL8lRvADhnBdIC0m06eLBTOBZ+B0G8irT9I/bxjJ6ovLpt9dnvMDsWzIqpVjN
FOAOlhY3AOlSnE/FueaNP/0vrcpS2gHmqyUvaI/HFKo+RBvqnc4WYnCyBsFNKXa1Eu8XoXCq01wf
EdXPNFDJfuQWDJPxjBmIrZnpThs3RwYQYNV5FemzxquuMOfYoYhIsyPj0YRJJUYShmbsJe+O6LND
0eUxxGGRZJZxM8Inu1pkcMGjsm81P4tGu26b1N0X9TTV0eK7enqYoP/K2xPFVS21uqI44kJBkxcX
LwdqQ0VMm2Sdz9rkDCwKOIOUGld7MkRHSq11ymRnCHp/as4MuA9zinKAYoMtuifQdbAjXI6xxyrl
TzgN/DiQeRglc0B7IduZV3C18QRsvA/i7Ai7DoGPTnbJyEvxcMXd+g4UmCZha833bvdgNSOkTmz2
NGQYOP835LkjE0wuJqioI1ucXLELQEoTlyrniFVYPngh8D8f4ZH75tbYKFbsCJ6PWtYQFv+PzhJ/
ZFsYw0xNQrM3oRRVk9Fx15NEnIA+mMCU81Wq7mdy7XjDQ2PyAUHXYlWLO/tP/Fymfp9i/DAjowpY
VR+ZQ3Zv91yMeylgLf4le3rK/KCYFOWKxBEgDwstiX+RRGMfkZWtPS0r9LWkJEJWpUHv4ugTLk02
Uow3b42MbNcOoSNVB+H/wxAX+zKfEHZc97nkg1NzUSqgF8UKDFkQ2JvNfzmlTOKSnHwk+gCQY/OI
Vda3cb/K5dwtHu+24VAQ88BIgav8AoJ+9c/W4hnHF2BzxkoPV+UhXxS7jK95w9oDKMGF2zXIr4DK
LFXRJ2s6AYrQfYgUWRt/NJTmLOkHHE2RORgfmj6r0tTslWoMNuV6IcSI6zvEkHryoCisD2CoF7cy
xgx1iYBBiQf/2qWPf8RbHCfbo2nLJP+xz1bjR5o8szcgODavZjhLAEEICHR85v5yBAaaflQkrKyO
XjLTTi9M/T9jK2R+7Rxl75d56e4g8twUSIUsYwjB7Um09cZhmw4exKIRc7V2Ux4RMiAtNGau7SC8
iG9Q99BpwIH8IhvcQQ4Vv1ZsjFcJznuCkjwybyRb7+rm4GLA4Moby6kv191hnGCt/9hzuxeTkFNG
WbJW+ZkK8gV3OolxKJxRFjx68AqnutR68MVE7f2F5Wd4gFI9/LHREMkhHHuPSOYtKZMGnW5KO5xU
i1IaLzrugONe9v/nVJP3EXo5daU/hjxWS8EY3tfHWfX7bPfGXPMcpgY2gCqGW9sZqLBW4nE54bRH
5Gd8F/WOxH0NNzDINynbY9BIMRBH4VrzPmMH2bMphERD/DPiQpSVvR5d3XA5zJbeCRSuWNwitY3L
+VSPRLx9TXbH4LrJ8d3Bau5uw1btMz2OQhoxWG+wHjEO2DoNmoYaf4aDKIEuNwa3u1GcZYwl22A4
vq8PA+6cVgfPzJKaGhIYueyXEguqaY2WAmKgoMDuKI6lpvCrkPf4oqgY+ZAcPtAu3Qj3fRO5O2CY
LHE69nMI2vZhYrRMZHtsOiNStzKfwe1QSo9+P7xlPGMJ0v3vuc6be9hESc8cieqLfv8pTpucW3nv
+wMQGhli9aXWgyfBiZxz+LsfYIpSCF5yi3l8psxEb7msnuITy1X5iiEuwo7Cc4GQwWNpXsSdjMOI
Y4p7uenDQx2BiKpJf70YXwV3GoJt/zmnoWJlRIFztIp1RJp3wjP8h2De1juaiTSTSX/uNv9l7JFK
Z/oROLDU8zDmMkM3T9KKNRwSum3nDQx1DCVtOxO8vUixapLr7wLJ+P7x2OkqAVyaZvjovnsmPRjK
nrvDbGLhvIB4NQuVG16oaICfk/bC0pbFpHM4sH716uzqyU8dB3pJ4BbSJ6NyGtx7wMeqJmDBsXdW
tdqxMbm7lako20qEC04tFjrKZMBccLlOKXYQjUXaXwKJEmxnYHDYvtWgI/Ej+G3DhNlFg1zMzFlI
reM6asPXLGQN7NfLqpZ71KxEVR1nZ9nJQ3ZbT0E6K9B4iLCChlJChiW6W/vsSyVTZAy7O3pNAhBu
ByYeqzgSJGvxvNHmakuJtZW0pZ+PEVHm/40FTs/pyDxd+mrqOOawExE4oY8sPaD7yM8LbWRWidEz
7v+sSxQUr+ILJOwZvRW+4qMNFqVt+hklFjXOiRg2UiGKLeyYuMXlTTnb60U/HUomTi9xqHBAIawa
FWIgeNX+VIwJdMKpHWOL8g1Ekt5JOuDPVKcVDpEGb4aW1Zz8kqWFfdYVgwjXdXxF9crbilQN+A1x
K1uM9RRm2p59EgPMD5vQH5Rrj/njghWRlka84gyGtxNcI97IGxuT8ULrjTDlYSS2Cg8NM+A6yWQr
q8G2sH9A2NnT7W1FlHFLR5l53yaexOhPftt9JFJ8FDVKHZay8a9Y1SiV59+v4O9NhdoBu0xaDqz8
LES1EY75bNFMkvvjUrtcFzO+g1/p+BKOosVcBZfbpJkJZc6S0KnAJkGA/R8bxfwXA2H4u0B0JU6G
FWK3S7zrWEGRQYtSuE95SHekM0zK6CpKWX9jc2ARONWa0E80o/JM79zp2QmNQpmDOOmSDAXp0tFF
vEag227o6IG8h6c3BkyFkmlvZ6iIiJWu/Aj21wBwa9zlgHc4qJ8hF3Y3JiP1ZXbwWDJCnY/yJn5x
Sl45Qqwwk8aFfq39M2st8b/jK4bspAHbnwrMxdYFHw5krFQ+fx7hLPeTwuWUdk9+nZViAwdwsP7B
ZKpndX05cp1AmjcowZx7lFRDUrdk4ccBkIWq+O6mBeO+dCcAsJCLlEFE2WAeB+wJy9fkOqPgFFHr
nJ+CJZ2kXZ+1XVFrrxbtSSROHd0FpigLiU0Hpbqw2pjS1ilHgCmSaY/d7VQp2V/B8MDwZWrEdBrY
/+VTZhpE6Fy17lf3krEIDPiAZ1qKfWt/ObxjuuF9Q9zfOPOIuVavNrvP8G/ZIeqpi70P+IKgmaBU
85+n1bAiwKptQXA5xNvtmXTM6B4k/4DS0RU9AbBMnT6/h+aTCVVmpHslpkP134DI9ECy8H4lcEmI
XGgM3ZjUu7taTkdE3Lk4eZCMDP0PDBE40MT7IgKSFHIznTF+FbRC6wsSrxp2n7tRjA6sFv+t576B
p9tM+AXblHIL9YAD46GQp3JuVBLuew+TFg8dYCrL6wnQj/6Fkt6t1X9dmWGUQxyR2bUfsT9mrtBm
0S/4ENaFz1iorj4oFTMLCPWzGaaXWkz60iZqC3Wv+frjN5p1rw7kCyBJqT1xPdKlF89R4m/jtxlp
GoV4oRBxJyk3K2zM3k9EcFJVg6VepBjvjcHfemArFP+g2rLvM6AraNIb0x9q4nPQ9Vebh9XOszd5
cO4Gi6a1yDptZBMqvgO1q+rVhZ9X/fdIrojtGiLnsts6qkrDvXNH4vGLNE3ADVhsZRwV3TRm3+gF
GVt3jSur3fTMh+AmL3SIu0DdzSiNPYrfF7SSCxC9Y+MX31gMKnOiWk0rU4Gu4ZKwbmtbYuT+KUga
LnolrQ1fwOyLhZwPb4bEyTJDsNG+nDFqet5u297QeDSi3nbJvHhELkjTrtN+ldS8kSaj0HbEp199
vIZvYsb5BRWy/tZVzKFnNb3LgC/QGFqqBfAaIqSL8enH0IV0JXko54oNUXaplx/K7wg7VayB8M4z
mIj7y44yuxb37cH3IydRpuJDCQGKyY8PmoPJLAkaFYrjiRj1W4xrlR5WV6Ei8BoPg+sxVWjeR9ZG
iMRfGXwe068g7C+UAQBdyxgEwcFiLEq6+rBbz0eAdv51/Vf1aZCbD+C+wPXC254J+NAERa4D3hlT
oqXg5Lj3eJBvuJie3qWDIlgwBnroCEEw2PHhdjNv0h1FVido4SWdRI/09W4gjgd1M3/QJmqq38nQ
f3kWT/KNhFIqukgIcq8kwuDmGJZ3SkbA8z4mlE0ObcSS/NCUXWaNJ0DzW4Za4Uets/l5qkQltKNq
Yvs7T7OgDboRiLfG1d3+j31Sn4f5KG2Il7yi8/vrfir6rP4XP1PFc0PG6TLIK7sEP7wJux6WqXir
XHJuNXJfezYORTacvgem8aWUjI2yWtooCFOEcTAV2SMg8tJA985C+RQlsqTaVFvFCi/IjJCKzRTq
BanddFJsukrFm2YvXFJ5BxFj1lgsjR/KbD67PeJdpWrAj+7v6/xhBwHiCpGv0G0vwBk5QCDAto/9
/U4Tl9Ip5aeeDtMqwBGftn0mjxZBfIHHHfKoLG18+YCFoeNhwDzmVo/CX7iMLFfyLgkXQx7rtRh/
x9qbDnV/z+UWcLI/fksLpbNRiXajW4hk5LN6KQQeiEr7Os7Oj2siQqzP8d9FTCvdfRKt8SV9uUxm
cxMI+IzRvx2hog006sLnRn6XYqI4231bod6J0d0Zec4P/AsQH8QFFOYt7UtQg4TIVYZa9Nw5oHTy
SEcbN0VII+1+KpHq+wvR1ghS8wVhbA46xOjGWbHL0LxdTpUvESv1fiep4cn8fEV4I0I3DdkM+Kdz
/XQnopleX8bi8U+dD+PluaTJRKcdZWLcBPKAUs8Edb7qGdAJ9+/uvlzfWbe9ZGvvEft9vLqx736O
E3Ge8W4wsJzYQQ7EoQfQSkVSNncf7cswCEZaRVz8NX3uVv/RKgV16ahB4A3b0RbQXc9q4NLLcyxr
P85kvqSU1ssg7GG0LJFUJYjYqDlLFe1uth9gCo2vxPJUnvHlwxVxpSFlHvYA4pzzCMqcj5yDbchN
pU0Hm4jK70H7z//qmYxZt35DLid1phzY3Lu89k5IPTYR0G4OQfJyxm8olcsZ6/xuRglmERRxmraU
jrERpVACFg3eYo7w8z0zcg6FILg3RaHfDOKFrGTQRS+LLPNBNIfpH1a3IeXb5emywlmf4AjJ/XrV
JFBb0h4UtO8BuUaZNHVGbae6/f2Na8WimESD4hO/C1coHexc6XjqobgsEtMi8GV5Nu7N77awwHuj
lUAy/jnUBS/8vQmufSfD/30cwvcgxaegnKwTy4L346Ljqqc9lZdVD+1MHWPUu8vG9tjvxogd2UGn
reF9qKQurFcPeSG3sIVls7a9g0e8OX1NoJ+7AK1iDfRnMkz/D9sOSogYkm8ea+fqOpLcdP7WllAD
Gtj36VQHcoIenTghBUQ2NDQ6Jl7URsi65kcyMTjk6AOg0Lna9xwDTKcLj8/i7KoxB0NHoB6dYctj
xq7iN4MCv6cqYLOVt+Pp81GqIslBkFoHmbJA2BDjdn7H0YnkzMF5cw4fxLRSR63eTm1iaPPOZNx0
tjPgXKCXoa7x7kSTBnLr6akDxbqah6iOa3MyNoCqkPcTLvW6XAxkO+1h4MGJTUviReyYKsPhkcyP
DkH2SWT30u5tyVY+pYwmko7hUToLOG6inP4LSlMi2E/DChCX9eo1Rk6pFzTKW3PMHP4JLOboKIoJ
wD1yWJQElHiRyrAHaXzgxa3bewoKv5qlGoxNVOnj76wuvoBiQddYLSqCQvRxBFGVn2wO8679OApZ
sRQ49Q6KHHJzF7rK7iNISUVhXZsCSuJ8oKvLiM4CgruPX4r1YXqdqS9zXuTwfnwuCmpcVbxjw7em
eaVhbBah2yJEM1ynfATeU7vljFR0sWLRJY/jVduygCy06UHajbOmIQnOiR28lroFOZrw20u90kCL
dgqW2OD+SBhSEYVCvQ/HVPuHHKZ9pVtjbpYjvO58YbUUuTpSZCFSByEXY3voqjbKlPphk6vViB8P
2rWa1GIWHQkk6KXGfjZEUcwZ+1KheiAqmcrTQ2ANlXZ/3NEj1SEyRzdxuhvkZ0o6iH/KFLCp8VIB
6jZqUSYuyO+5rVadL2sqdr71MqiU2AoeASoHYt0GWRQYfQayP0zStNKrActmjbI4hmFAUukolhT7
u/wjZR/dtS0BBchESJYlQvZBPk/1hDXk55I1ZAqK2ZAcsV9LoQDqx3hihYyqG8DNXS4L/yw3BJss
fchcujsVl5vumwI+UhnjUnxzKYDjttdmylCGssr/BkWwjs6lNoKyY78NZyZyEOSQ7yxIA2O+YLhG
IN4ONW/VMNoTzumBcOcjxJGz/ICtBTHxLEA0s+m0uYjWjTl5eq8sBQX4ZiFy+DPq1YgjKwtUELj4
iI896Cp70JqeHRM0qWuOOEuJaTxlGHtd23phCpS1z039qFefp0qBHfXZxSfR3XxfiT8/qa7rVwck
zwCAICkzCNQjQRLZMdvOuuGwJwBj8RUYTjF4TyD/YO/uO+IycpmrF2iJlHqTtDhhZPCIBFMwrp45
9GRCe/nUJzuSpQtw7qacDnKv9EwNCw7BziBos/0VLxidxtYh9uyBjqVDhZBWskluwj5IWA8dRTzQ
XWvZE/upJnP07y5j+VzqdZQ6swqFJIjOHVosHPq+Tx8LhpBYO/wxTSQiYfNzL+J53CYpe3BKcyoB
Mecws0WLrcLGqxNsAZ8wsn+uJYbkjN0f4sZnDs+dn2VsDZ7IlebKOQ39yOwIxfZA/hzGsuDYmaRu
VNpdITW2LsQgB0m18cnZKV1S5I3F0pF6pizqihC0wwG1Lo8oHl2MXlPS/xgRaCgmbQJdLB01Zo50
169phnF8AKNTftgepoLG1XYOJSlfXKxGu8jq83qhsdfLWJzYamqELLDTeJYLTniwqvcyCBZYdaqr
wEAAWTRm2pFkUqJMsM8vlQgklQd4BE1CrM1JAUK14CcfRwYlzpneVdNOh6X4MiKX1FjkD/H7dplL
GSbyNnPyRVhTA6snSQgzn/JQK91b65QgKONFAXakM8/Fy8LLR2alXqmo3fNtWd57GHFJum3XsoTP
yxz/JZGftVmKGwcYh9hvDcdlj7XTnTJZSemVnVDpZPGuyh8SrZwwHeLCx55uhmBTTiO0+pEGm735
ACIXWrQ3szPoysCHjIuHhpk679yqiwqp0Ot+dGsYaBqcX1woz5uJ5o1fWUNU3bePL5o3MEcIzX3f
8g8Ll5QpZvHZ2sVEfW8CPflVudBtIYEmBGCW4adhDTEMdAZKe1Un4EVD6MDVNmqyfgyIrW0u9djp
xcv4I6kVQHWz7H0PxjWGhjtFX91uCVLf2m8RO7cSDqI7CorLdyGhQ4mhcK5qxsgdOXmYgJtvjSTt
smD8FLb2cAiaImDzIUjMj5Vh3eVZ7yUK9CMlsY6HKUC5N8e7ecmiP3JRrfEuEUqQ0YvdiK5Z5uPn
RrVv6RDrV0Kd7+NPPXNzu6yoq7nrTvEY3LyPvTvQgfX+Yc3tXl5ZGFCo/uUJdZFlRffhxs0X/xYd
Uj+jxpxK9+E6kXVTSj/KIO1rMVEfTWWu8y3qR8iI555sRWHRZz9RsjkA3NLphUwJYF9nzMH6SjTR
eGKOvaj8aPzQGQT43FIXevrm4V+OcX6RW9SViN7pQzVVZti7dooypt4/zRNHf96NdVgdPNEea5Y0
y53yHjzEcPE4DnY9wzki0v70RCSQp+FvZVYG2hddQwUf7EH93y9xNnsgIO0ZebngoedwxNpyOKoV
CqAPaL+KNUaYdv2ZY4szeudrYYvme6GQXvB1H3ooKTk/ixmi/E7rsddX4jM3oafzqvQ600/sPaV5
g4yFPw3Rr6rz5Dj9p/VXT7ylbr1tBmG3kmiT8h6r8XobLvfosh5/2hvl8lsjsNCk7DTmvmAZLOTp
zxupYCeM36qx4Q24NSU5+rX8TSI6agVDPISVbcXpCNPRanc90mW9JxVYjAGsiEN1ZJdCD5FC00YN
PRv3phG3/CJsAFRwARF7KDDS2LSW/+02mR/rxvordxjgjTk7lGVFeg4bzkX3Cf/8Jx2XbVRNRET2
08TYzbK9fNt7AqUf4EfKN1jwJEk8s+sUJ8RliIdpceBEBlU8IGXuov0IXDqOUtsUNF8pvR+kh8LU
s6RE5f5zI2QClTb9y+aLaeTWA8OCjDc+zG69i5rPefV2b6e1ScbJejjeysc4A6g2WRN2NGun0bc4
yiob3HOOUnYgzolsyUqctWE+ZGaWFt3gqMRDYAXBdGx2RlywAAVvxSinI3YLsY8WU0qFFBc+fJEJ
kDRmpv0fICJNhEjlpiGZA0u1tq/mImV5kj0/Hoc9870OKWCVjdI8cF3UmjVUgrdWXD9yfDKlz3rk
knQrDV0AXThKCYKAigsUiRdkhNW7yRtE7q3kXGQhCnhob1XHSD9xihkf2SmyfftvtE3kxsKvifiZ
QdvgRWH1rF0zJLixZajP2Cxa/SabY4Lh3WrNh5hYtRZlQJPVU3uXdJO8j+cwmyns0WFmuz3x192F
vbj89BcGG7xuaMAb7evavI+u5Zn5eL0BISLSVQT/pIE87pwJj+Ie+ZNudWOtAMs/RmEIo7+Bga7j
E0D7dNPfttynq8huwdLGQaRxPeCQ4yATtkE+xOBazhO8CPMK2sn69hnZ2E5Qi7jJ80+R1eLyJ5DM
OvxIxtxP+i0Q4TyuGOGwi7wkVdjQtWWfefLyd+9nll3I0CKru2l1OWArwbf0K5VOWEEJ+iM8AOhu
lnPKHwqw842xLt9jhHibenOID+k8/QrGo91bmJALCjoj93T7oamYjsj3hMYHSd4cgvGSsL1w5Mo+
jJjZBGPozQgfZyUatd8rfmQthCDxATrI3oOdm8vdnC+7c/+eIwyaL+kx+54eKSK0EtK9lgQDR5V9
6UalSBX2cnMZz0SOq1av3ULaRqmAdCVtzYVucdKulfWNt9ltJBWAlZBC7Z8ol2WGBjlO7lzXSFU5
mS7vKoP1wNaMlms1+MM3TG8rlUPwlJuu1IyW+3PWK8t7Hg2xVyCBdB3JQQDINws1i4NaZ9kHz0X1
6rgCrXqhHuDtT2bpifmGe+76CBce/KfqqIKlq0qakz58o/YGhP2nUFoTS7XarJvr4AJb67g6gqhr
rOVLRHvx6tyd4bBj9TOomS4tzBH6jwzxud1662ZjZxvZfwQS6Tzmc6BEAp+pzODqnRg8LLqMz/EP
9g12O7gTeYlJ4v83+y/c3absxr8mFRc71P2hm1zvJpGrLHxUElBmMV5ovwe/xkY9Sk25ZgkRMASU
aBaZra/LxfdwIgbEJqRC4sel7e7MiBwwtnZXPaRYzM6kkbvAKqQYVJiQHGc+V+pBhXYrWDG527f8
9wG9VKF8QL6Mhpoo0gxhnLo/0gQeH9xPvLDEeySJm+iGfRNmAs+ngTIxFEMbI6oBQPqY3ZWlqRJg
WLxs6/q6ZlD/TefGolx5vCjw8LawqW1tJiT/We2LyNKshA/xfHjtkoiNMVOQPCk8n6Xxe9T6Dr+L
/ujYBlC2iKAcZczDlm+nbfqjAhwswGURBIpR8DhOpVbLrRKNTkf3tdLpsBy8dVDt81Sy8w93CQE6
oKwwtvu2AAc/92RQqjPlq7BTdwuBUeIXo0d+VT/ZFiGDF8xKKjfz4//xFUi7Ypi/syyTZdoriCjF
jshdvKrRxZgvLXt0T4ZB5a+WMdUsbQR03HoyVSuTj0n+KtM6WiFNjvfxpQ2cBguM7JJIMysKmjie
U9Shsd5dix86kP1wfVT0rzsVNIlRPUrjQ3a8wH9JQf5FBiF+KtquI6os0KEhwRafhATzyMg/K8t1
L2Fd3C/2Agh3BeAjxjb8fusLrYu1y9k1wtR71P0dySmy8zCd8kL7v2umhDe8vafJokGD038X0nuM
KkkAdnhajUgB+oHgdVgy9ycFl6NLUMnZPmII8twBJeiVf7VxhiWLkZTh29faVD/acq9WIdaHbGoJ
WcxmHEelXNd6uLRLyktI4VDaOv7whg/hEcbkfr1BOD+XqhB2YSbC+fvU5+7W6RKssCUVYX4lc+QB
n4236TZYVJ2AKcIEFgomFOTFSLP3iV/9GGPjRtlKU05f2Nf3ghAnB2XwyLCkGI4c9d+y5lYvwI/N
XfCyXdCooUVYAOZAMMUhflMvpxo/Py1FRl+Mvyv3ZwxpiSKpHUmg1UhFInt8sajSLfm4puyleKU4
pxY1dyxrkhaCzXtKjsSBe/byS5sr4UUTeGMBpcT9sKs8F2qP7MpW9LTllpDnefH6szNuQZi3ZP9I
OuJ74+wXvweDMuNCRMrzKmxYGgg3vRiG7OXgnrQ4fIYbGiNwRtBGgNBRCHEHFVt44BJIgSbgQ3Du
IG8Dq5RhH6AWOqPSLzPZC+ajEqG0cKeREHVz2jq49KHPPWe306b14+WYQ1Qvanx6n1QtI9ObArUK
6OvbtK0tGESYCLbmhthyZNgDVX+UX0lr6GZD5/1ZhwDxQCH6vJSkiqP0dPKJO9iGLJ+T7PpmSjmz
Y06xqUtK9qiQ2NV65Vz7FJJZy8y4iAvV+8JCxRH6CLgVTusVGFQPSHk0IJHo5y5w/AB+Uky/VFCU
WeqTdf18j3ibuDE31ryOVdbd2uuFJhFCUidEgXGgYAb+LLXTHhaObKU0hCH3wC0DKsyEz0wAmydN
tBNUd5HTjnoFbCV7Ioy7X9HVNXk5Ls3nUZ7uB9WE6T5VfMwe0tX3B5OnBhY/IBgVROjxJlp6SERz
2KJwymMt7q7HEIn3slG+tcGSMCMisvMQgWZyC8B0eaDj1KUYH1LgV6mgJeISInCXW2SIehlrv2VP
7X4Y2KvtI650Dc2XPggTVyeKreGcjW195W4XsrkDM2z9DKyNCRpcfju3KPCRFLq/9m1IAkrhDcEX
W02RfC8hhC5s/Dds9NsKQvehXUKpAqmScBahlme6XEHXxhjPY3VJSGcHKDxaG+M/mv1Bo80tcpex
kU2IGPzoNjpi5liEcAz0NuxqkgIerJt/ozvpN7h0erFODqsbKsjQlkXKOZ7t2S1T/8gONK+wur7w
JbvCG6MhGsRuQ2gvM4VACzsH0PPUyGNoB1N5YcUHA9bMMz94D0d9D2ex4V8C2N736S6H1AwP5evk
xhXuJsR00qzsrVSNHWp6yMOL04YVVUcEuVViMmtmEMVE58TlBr2cqyy0yK7VLRolbUBcN7KqJxIW
FMxerVqT3JAH3/E9bjgNWzMaBwIV4OqSprAiKeZdz1sh2LL8UPdZ/zHFPmO7otaQdkmrPhXHAxY4
6IG4iKofSbywvJSUGxfIfEr0WBh9xKZxGEoqs8879pL8Se+LFANjSjNuk7vtMYiouDqqan1BCf0M
q9e0iv8S8JrvniFImBiNMqLAYsH1QBhnYibT6l3GadnIDcwvvHDM7750+RePNOEhUEUCNic6s581
3A0s2yFtkGDC0TTISHACM5Dyvxmqni4UeRfCljwq4H2vcxSoKdxesZgKqO8V3OMWMYAGNrEWd0QT
m24p3Sx/bnKbX0h6KCsVeJaGe5c5Sh2lJK9AVVy5GH4pnG10vT4u9qrkz56uERxUpdwUGLvGiaG9
l2lQAs8Mi/dwQhc5DvMesNs7JsqAkj6UZaSmYMZSOJhKeeYk50YGMwqkxGJOqLf8/vWc+qSFi22H
RWnqlhkMelpLKsR4o/t+M/DO6uyWr+/aJdAGCiqZyqLqTOJCm2pmycPsaeFTYDqZ4ptxNRsl3SIW
1qXq7BpeCm9S2Lxi/sr1MPbPqECy6nD6wUWkkt/Z/RBFTPgXK1Fdnwwl3MjlRBFoG0gB0JBYpYsY
S65Xz8AndivLrZB3XJDBQAWsNjl7R9HTzag3k1N2yPXu2kWUlqyPwS0Tuduq2IiK4NjEg7z2F7vb
2JFdAdSX/n/mN2JPm0ImRpqCD19Ehk9yvg+mCld20xe9WCDynR6Axgcsunfbl6FCV6a941xoQxIl
7kHeQ+OgqeGv4iotWJRCf+ipRn7xIhwqT1+TT6xnWviSNF0RwnfM/exxXBznwEwCVN9SqxrOVcdH
SwrPZiZt5C1CnPME11Czm1dEsu8lMIPF648li9sUAf8Aj5QXjnUjRUaFNm3826FWOacvG3Nzz7OL
8O/o3r+VjsV0OBPOspXGnQz7RcV4uFI5vvxBQ6t+UH6BlqQldQGHaeMiWe8PvpNOXJGIJ/h2ev57
zT5LZro+0LVGuK4gZ/jU0KbIdtz4AiTxPFpoPH9GHAu+jSHugd+PdO9fmUvGrLuGW/YEN7VigUY7
bD7J0HQfd3el3LgxeGsL3VpvC5g9SWdjmih9tglEjEQUEz25v9wXLoUBvCpAbWwHFcHbLLak1sA1
48iWRgDdPWKrTmTJJNbiYGb/YspVe+s+1O9Lxews10HT64qGaigk963cFPfc98wOz7Ff975tPqjg
4xX62Bba4rio+OXSf/K67sD3Aw6xFeZtaBELsMHa2APljO9fMwnnd5J2IdGQfTgabRfjnOZ4+HL0
KNhxmA/bnHcPPCzi/WUC+Ky25qw64hCJAga2acPkMSYI7Wo12E73UW+NGEmowBxzb9iW6Uh5V6SA
SK82zRsGtu4onlUx7a117OLyyTmuwmuBKk2thydrE1GOCS5Mz6fHtsHb1/hfUvUjZ8kSUqLq5KlD
KqDzg8PPUp2/3iI76cbb5y2DQWlzpeDBc3RPIikN9VcuSFjUt5eKt28FbVHAENy7wHjtRKxWvD9O
xYKbi8n9MGcTq+gNGbiQ3/xSf9uxc1awoDDBTznJ93iFu7lRzeWRi8Ug0Am664x/Ry6xyud69k2h
C13LHdhHU//HgfgI76gg0XIY+pY67GuawvFstzZv8QEVbihnD1edLSHLb6l5mg5vqldn/q1qk0j4
KV8pG5uRvXCWErNimPbYzq3RWG6xuotSs1GRsqT2l4kP3DclIOqXpUi/EUjdvdtmgPFM18hmJXCs
hwUwdVl6fKsPSiwWHUjLHJE24/+TJqmrBlVlCdhaZW2oVfDHu1GaTWZyqKcfzl9a5mT+qdysJn5Y
c6G02jZcPcW1+D8AYOp2N00vlE2PMfV2BlUT5X8TfVcGo+JxY47oaKRBei902sTfiVe/xG3uvHYv
LFAK2xvRqxVWnZf1y1AywFj1QWlqYV4bndqQueUnlU+b22ZjZqN3zmJb5v1ok3Y4cngiucSqsquF
9ZSpzHQlJNl8h/cQQ+K0qS+WX49Uu9h56fQJm/ZaLU8MpMRT0wBBoeFNDreQEFOIyUqTRjqQorib
9ekDUFJHRkNXu2Rug64h27KRZujwkB5j5jsCIi7BiP19jurk4WF/F4E/ZRD3fSIifI3oDA92JxmN
wB7xWbBHF47WtjoGk0zfREkc3N4eWRianEIaxKkPfOln7JJMC67EPTBobru9VwBC5e9jABbuKBYo
QNZaepNi03krMDs1045Oa9XEhA2OgZymSSBNzyVKiTseBw68Gsnbpi4E2dFABVeX/0RCqWBwmKyC
2YS6Dp3nBRx3IIQfyKl8kR/lKw8mnvY/QfnwxY5YQpKJDtOB/sPJpDLvk93dJ4vnMCcteDUyqUvl
IsVeBKb2e+KkM7DfAJo/WAxFJ8GLA5byUe9yUqKytODuraXzndMe+8y7ikCM55psib/KiLtQVeoU
pNjoXpPVVRHitVsjAEFMOLzYMhRdoagkizoDnpQn6OVHrxg52g9uCjdveiMHAV8ghh3jUxYFC+r5
axEg7tpeL08yob7OdhyoR1/30jD9WJBBrodljBkDMTvYufwzrHvgU2Bo7tdtTCU6JOMlUC+BOLEr
FKRZ1+pqz+5haWGw6OF8PoB4buHbx6H8vzuDC3MUm/LJfJpsNAGMkYVxrVO8MUti+c9gzqtarlnp
1zWu1s67QEiVFHhhQ8tzBNHrSSJDVk8+5U6RLoQ9IKjj5CAv1OSzQYlgGhlxglV8z6tKnsQPg+Tx
C3J/zuFK4RL7t9WXFVyMIz5las5FpEGzl42ms4PaWeIoL1JLaIJEvKIQwPsnlh4KdkeZKH9pGBxp
URCOhYydyDr2Hb4UZUZpbYfMj7mISyNsp2iD/uDTQc6kZ64ANp+7L0rWea6uUpImtxuNAwc1ECqu
EnZKb6LD7wGvu4Kg+PNQ2KmUqYwp0NHnYP3SK51Tm4NlxJxxS1mEJM8Vo3taHJ0FVpqOBYr0lANx
0FplC9+vEscYL6qN/7yrTrhZC4lyha2szsumrvU8fPmhqKSr24NW8Bp1pn3PKyyg0A75TAalzksG
bF9IfJA7CK9BAAACJi1U3IzR6H/xpw3sEXT8jXhTan47AxqBsIfD92eZi7TT2WoRyYnCEK13ZEFg
sCUCgB4bqI9Evjm9kDfzWkv/nRgAKF7wvIlBgXjEPNCBJ7h8vFJXeX+yRj3LTAjaGnX0F8NFIJQZ
deXd/TaY/pdEPW74EJRbNkbQ/dLyz6oHNTWXQJIx68cr/4o5ZNUa8OUIns+DfZiWapVfcMmDLgnF
ZizqyyTSFzZFqD/JuZAoAHNqJexwm2rzWullsexEyXti/TOUNGdl2oNKtnmcP8aiqN7gzxsxkMBS
IVmjjNid3l2Bum0qZD9UZ2ssToB2g0K7eDAOBZmnX1fP8eyy2MNWNNAjYAAUuMatYMl/aiZCrnsX
cir08AmQnxsVvDJG9DuiJYXoQvLyRXgZFVck2/qgrZ7KUvfkpSgkwrXE67iclW8tGdKsYuG4PPTB
20Lg2BDoBCB2ilr9wBIaiADwUnK8afqfbGentqwqp3E4NNkbj9/6W5lfloAjfyEt4m1UxusguW2P
gWy4ogsK/HDA+zNMHR7IBTNoQjTvRubLOtEeekQ1OB+i8HwQH7hcZs1/Tqn+yjSp5dxTF6mcOsTO
N0zAEZCXYHsxz/ftkVHE/k+61G5mVYGTLxRohwni/MuNZ9hHdNiCsH0/ruAHwmtaa/w4WUcIBmNz
AAr1dReDM7stjrSuFj6COthiwnCR5WN6Gm6wIBQwZyUrTz2kCdxdw2CgO0CwdSe5mys/Q3A3tmL8
IBWMq9u9wY7UXh9S4r+H8kusi1MW7lqPAV9pIOXtuGv68qx2ab+sqF5nY9nmPmzHdd+gelkEmamK
TTQq9/6Ine3sjxz1NRkNzrkDBq2lTN9OJum6mEPrh3Cvl1yNPMBru2P6QiWuQUnP0MMPuLvLSmhX
rCX9ynU+A359uZpYffEqETGp9e8ehSzK/AAgiPRRywuCKwlRE2Rj3EffzfCBrXek/cchIzEHTTK5
sndI+CMwEcnsdNuOfNmy+rW9F+gpueiVoEx19mcCCLVaplZDojZNfJ6hQtV1bKM9Y7hp/ugGJTbV
v8jfZ/sIyF8Bwdn8gopV7dYowRsJWGoVS3kYnFbVxbw0zNsQB386A5QL2fqIUsDJiNwymIuyQiUF
A16O36qExfel/vP7y5bJdEzFLJhVwUjimD/O65HzW8KfoWxkz7AJb9iwu/B/17ROpaVNL1Z6JAyN
FL3xWZEF5iQVi4sT6CRz2SghXm5vaHQiQxKPNfCNKrJtVuqsghPnPHv61Zk0K+DZOIO+2l9KeLP9
O8MhFfc5E6qcrloUTG5vNtcyBuPKJBBiwwVu1ppzlMcJlmLgJed5EiDbzuuyRyMrJpP8/C1pMP3W
AAOyjVSJ1an/pKJYwrhQiEwi/4xgJb2JgnVeTFvu1qpmhTchgT257FInbLC6jXCwzU+ZrPlJUJe8
/CAcDnZaildWSx/u3zcpd/th4GZElysL1Qz9GYerCNmTj83Y4sOoGZCLAz4gfkX4OEw0L9XJNAs7
howc859JeGh8zCvoDdd3/6qzF/OTFVwx95akXsgpoX9HxYQ6Iyegw/232yGkHRq1a645GXNcxG/j
h1Z7Q0NowhfHDRHzHuomY+lARc0Z0V+e/ptcja7MK+SNwI9m0Vevtq3E6Zae63QpUkQfjcO1uyXN
+2yrXmEGo3lgVl1ui4S3NK+vnNzOhdg70Uw2BBb69PZQERJr+5AdYPK2RveA6KS4OANHAeEvATe8
/voH54fSYAuhyxstSzxVEUSL3BbOQaUx5jjW4fYmZzKlPxI10M6PL+acvHxYmEKK4Zncdiu9Nd4e
dEUsCAqrTIf4Cr0UviNm5OO4yNemKtyBxiVJOE2fzl/xImBXV52jImZUl8mhjQPlz5QjvpTaA1LV
cqIxZ6ImrgMBCpB5g9/bTO9bPw4U/OJEvVMpEjBWlRPX6etyCNlB5DGHrGMBV4xdhIidwODUJxKZ
aEIZBZdzzbnWjZp6dZfaaiLu/ijzFBluOuvRpBfjkAMcUavqRrCHToKDU8zMiWAmXr3a09rjER5S
861RFhyWQ/xL2Z3CBlN51vuGgrp/7CUaaEX+A1vHYa+qnHgHbJ7Y8azVadAHjDEhKEE2+QIZ3fEc
QqVV8Fpck8nb5TonCRmkOkBQhBci3/Di5dIggQ39xR/SFm4R4QkgvtByJwSlTLxG4JcBKhQzI1q3
vIImo0g92fPPf3eAPLoXCpe4+UOR0ERilhvUt405z1S7c2e5unxjHidU4Xl0qRiTGxSj0DwUJHlY
UXfcINiHvStkAT3i7/xpsU7gBn47zoFC0bxgRik17jGvR1JPLgx20nk8+q5iSUnC8oyQnU3Thtbk
HpDivEqv/n2ikBykTMBnVoPFSX17c0xDcOB+qbXjaUMWI0SoVyIpsPJHGyL3nuaAXyQBA3vU5vsF
6e4Iqj6x+Xo5ng5Gpnnp/JRo6ZkNODcEaVxFdPFgJqgs45nuu7UjlqdXRYvL+AFYIIMkhTVihm3e
b7Wvc9sb4Bt9aaNTtL4WdbVncEepxz02iPQBGcw3V7o67kUGqUJ04ldojsrudXyelQVfu63lvLN4
R0ItpTb62NxeqRpctImNh6svTQYAFTiCtE8FKkbNTQPcNOU1SekUuMh33cfIet2gJ7HvxCZ12hew
W/VpreRc2fYP9i+jgVeOWUcexK0iYtaIIKidbYJYgdg41RB2u/bHYv+j86D3vCoXU8exHiO10eo2
JqSSFGNu5kqfDu4YxWSThl1mQSngkMz9q1c4MfZ1ydi7YRRnV2KY6t2xrwxVi5bnjxkK9qGrkDXL
q91Yt9wEg57KpQTejGUiK/tXY/Lf07ZnL/jzVpQx69khGdaxHo/JnAWTJ2Svx+66GpjiiZxmtKAW
lhj4+AGCF6/1Soaw1Nzhf0KrXkKbJKyXn0lqAMxYWddBrvTz8C5kaErYRvOMN9t+Ie98ktDSCse2
HbAdxxLN58DpMTzKWJwROWII8TshbECIh9L83ZS1iCx3kfycjMUeYOIBATtC7hQ9+x4VQK+4MBHE
+WUWx9UyeqpKzPzCHuHjvZxV0MSF8tPsM+k8a6ODhoO+Ysej9RtqDsiuKEpdOFyRzb2w95H2eLj7
/HzPq5DO+xj18rEByAKm+Mm4rE5QUCWx5luOqsqXT7/qANuMlmQfS3q0c+QgWMGudR2Z1M6W1tI4
5EiO6lMBd8wVL1JmfG0bb9lcSVgsupiXcL4YuUAfs20ZITnJw+jHS2ZpemGdim7MlRPi7pUhWMlO
m2KewNvYVqAoIazvvCbZqboYOmOD42kVlcSOg1wx2ocKAtQYjfDkx5DnwM3KGY0p22bAg80Kqp0b
FRp4ffWWyUhTOsh2d4Gk0YE8t63dk97X7q/EoWb7WKbRnAgwA490D+wk1P24dZ3gUVfcnUvFmsM/
Nse9SKFKX7apwM1kVxNObGY0vHRodTkaEzg6bJ1G6FspUB1X+GGP96bCvO+XFVsBj2pdMy0+luY4
E320Iy0p6QzIb7ERURcesrO8RLSF+YFEgkHosxpInpgS6nmRL2TP23DKNQ3NYcTLtWgOdnHA5ZGG
d56qCQRFD04sjNwUB04HtKZgXriPJZq9R/mJzLbJ8YIkb/71TSTpyk6A4v3Y6M9WU5QXMrTAeMcR
uaWN/rdeMIsndbn8ynF8oSztuHNMI3iTFF5sy88YBD4bVXVXBN4EER+qOXHosAptKSa0g7qci1Ww
8GViXkPV0D1mcUKOyBx/eilUKjKX0+4U3p5NUQOq4lIS85qlNKQgB4qPqkap91hwd5EZRBLZwK3N
rEBV8srjmsh8a2I7ns/dJIWsEiIDgFym+USFszEu+XnlI9tM30MIGN6ID8gH4mmdIsQiVzCm1vLR
Jkp1nY8xfj53aHA8o4zCbQTwYh2NiKVt9qoSqgh7HaexHwV/Orqzh5DtvvZoHSGIGTUy/BlY/+Kd
3eUIYOBoNyh/ZiQSlXSSFgLVz6ExfztSXpzD2Y9ytRuPfS3cCjy1TWsKetGIfIxf5p87nIgI2i/Z
0x22RQOE9QeJEmtsiJk+34hhw3pLJBzrY1Jr6y/O30TNUVunstSVO7YwzOHVnjTA2T0JjAslhryo
xWgaX4+8Poo6OiC0YyRAUxr1x6RDbaf2aVqbWjFtB9LFAw3hAKyK5JEpHT4AU+iEBsXjor6W18e4
/vKqeX46bMwhUQkhyMifGK+/SsSApOeY5VZVqgBKSiGVJV32TByHDY1bJoSWJfSkfz81pzQ4EXTj
iyjpPjRStgXlOUsRz6nDsAKE2lzUvtmci+9ufNeWSMCQkbYmvMTPaeb7jS9Cu9e76QfN6UpLBYB1
EgXopIk76JfwCvwku/fxpHdPMS8DtYxeTfJx5+lgHMjviFgcGshRCln2MBUuftDrkWoSLuYx4uqF
5iRTIU436MMVLnxWdQTLx6Tl3abjUri9rxB8JrVTtsbVE6pQoHj7a1xzZR78ZnFRfxa9khF9qgzG
k30VSduHGUL5fCQ9C0ezKyNH7T2VKdfRf+0U98kcdCxRqWoTKM8daudwLeMDuQCmNeHklU5dd4E0
eaOFXL01nTh2jFUAGh+gkUuuJTdviCC9yOnmNhSkfwuKOGFIAAC4zPdQ7lqRFjSxHVS/Ye3IYlOy
sKfEnVawISgdw+ZzCq/6kqxMAJcr1kguEXqW2VNURfYlIMnhcnar9ptwU702Q9AHpfINoZAOVlyc
FCmzkN071jVjd305dKCqlTLwJZKZIN4xs0w3yU3/nBvnEnld39kAk8hoIYw8xqW0MjpUx22KVVlH
BXqCggVnyaShEeo5XVLC7cu4+2BIbJnKuDi1FvUQt0PERnoO1zbWB4eUtVhHOnryqM0kTHOOStvd
j1uQbFOJtZdWQVt2nSEvia3vLJFSl0cW74Zi60JCRuj19RRpjhX08ZyCn2dDAEGnyyOipSMqwBb1
mB20QCOD202lVHG7BO/8jRGt/7CLgfzTX42meQa6FPH85AigetN2FoACbfb/ncEmHI9lj6xAl4uR
B5+qURCTA1Gj7wkWPkkhNH9wi1p01tWWOim4juimg+tEpIFGE9x8piiGejNOE1XsZPzIcsS6XOiZ
CgHIBYXs5vTCW+I3D/TzNy8F2RIcn/3gThCHyxOARzeaAWd2bzmWXhYI1GM2WY9eSrFXBo9T9DLU
pgyeit3wC91a848OH43DgbX/6LDT5BpjgCv3dy5IoKMJtHwwrFar32bm4PXlvP8tpjosTCxXcjvD
7XSZQMdw5st0gpNDdDuYavwe8D2jx9RZI0z2wqShl2KjLmto+kazC7Mit80EbpNo8XdAb1BrlpCI
wHfV2Sf6rTlqOEEy2sSp9yO5aFSfrCvGdV7LlhnPMazkM5Kj1f7FOMNLbKmmXm1DqlpyS4Z5wG9p
pwIh2HwXSri1XY/zTDX48A5pcE0q5MaznwO3lDrce/1foM3NidfZ7gZynXcbzQSw1ArZAoDzDxh9
PzAUlEHP0VNYVVgIbHfCDpv4NgU4bkFR14vRF3ZQgqo+I3f6XUPgkoURBE8Gy9YnQdvh+xqAHfDp
y1nCHN6ZDojtb4HWKc2KZ25IKtqaaMJsNNzrh2SuWtXde5V+ynVmjgBL34FJuxLXflFF71YcYmB8
ooSC2dennJbVYXnzV4gxW5aerPLzbPOk0FWg5s5XzC4VcfCH2+Yik+EY028hLYzit3tD48rTVv1U
JDlnyKuVnhQULaQrINwTexUWa1DTO6wMGx5knae1WNhLRVCvxnZlC86c6GhbuAQ/3iG8OHNco+cN
tykzWBkgbb88lgxfrWel5FC3+zK1wtuu5HAQPm2wVegZj4QHqDobIWAxQfY28tyPPAxkig2Dd4pX
GNZgIbymNOsY9zyWaWC+QGAUg7J2FnORWxzN+GA4tLKwylMO1cdMXynVoDBLqv1/XEb0wDr/SlbH
Q39t2kqzwpvg5QWEg+4rc6kn0z3220pkPwFtnphaHoWgRy+USABmYmPbVDqR0faKkYF4BJNNpS/k
iNdfuQ8CHIs8INDuizMuqWWD/ris9kCqOSmhz76gtDSNowwxA3ROl7GC0gIV43keMoWmUmT+tu6b
FPkkxRdX6q1RGNt+TnCF4zD7kTbk1FboynLdZS5034cvK5lXJYkEWj127z3eQtWhQoVljk6TAY8p
BNaWTNDAUH7drmvxKf0F8TQJt1wCYPUF8JMQGGLTwzrHnNhpRqYQMf5oF3MocCeBHxWD5rR8eOeY
u/kfmBtutSBY/0cc1g9HKIRxcCi8TB22XZxA25v9MSmr51YCcVnLrJpKEySg0m+ifaFpVTboUsqb
I6v8kWimjiNzMMln6u/9vBa229SRrzgHGzi1eGk1y4v8vhhaDuperG/xCCylfG+Sevt6xSC/+7fp
tofDg0sgYq+2vPnqxVzoFmPLu+ZB7XL+ZJiN73HOdwdolOvfY0zvI+Q0eYFps+2ipRJIfrNjVmp6
Iv+1gmZNDsW9gUTOUeo/mlRSFjc2Xlvbth7f20Q9NCGCEomBV5eiEOe1G93n97MFV5IUtzC/CDkx
dQs/qO13H72qiPuI0xj23uNazjC6quiIrKLdxN4gEVaSS+4pvQ+TmkvFzhQ8oVoaLo8f7btMrPTc
sb4scq0SyqQ4IoZrIdTL9SUThL7Q0Pd+PlO73msPbG5Qqq3BvPmIz00ugkYabukQzTvppuf17LM8
4/1fTPmOEDXpXesIVD2plkfJ5c+AQ3PECviQLe8A1Bvpx7aUcGgcsQC1/ie+V17cTBeU77ub8HAU
DW1idtGtUvbo9f+XOO5sDuzwwaBiYXt68g5/2fDy4cx1lcoqfu7jbviMrEQuljO5r46zViFCWiRb
T1Y9imRbk34lAo5Rp+o5Y77dbqj4DPUrMXEsVX9cjZ4CXJYfAIhTtSWUze8VLPMT2koqoxN+JL2o
KMBJCD5Y0suInWM+5cvsONMJAoGwTd+pOiTm1ctB0qWMzzKozdkGasmuueDcP529GtVLKhwpcQlS
92nd7Tk8Prt8fi/M27B2qs+pZUKCFDRxospjvEXe7/SBQqrkyusVLkLTRKgSFRl970lC6YYkuoVP
L7pbE3ZIOeTIxk8czuqKGdqo1IW2ZPnDFc07wTVn7tpuYCyxAmL/k3EJ6UPYLhyvyPeimJzxN3/v
lvQPx1N3nbSVknps/QO24OkVNhsbM7bBuY6SZt+oZPHwgS/KsZkDj5FxgqjbaI4QHv4ceClmLIl4
alo2c7xwGufw/pO5Wi2wfzUlSZQlYuGTUxxbtYkOE/2xBT0wVpL4yb3y9T/JmyNrUqGZ0hvK8LKL
Sd2/P7MNABgAddFaCfDhddXhamkiQDKUol6FtpIE91FZt8P9xXutLgZKj8R71MmveW/nGTNIuHAG
Mvds3+tFIKiE1nPV/M+C7RpImFKyaPgzxaH3zYmon+d9MBAjXFVg+fEezL7ycoN0C/u+rWesHC+U
hhvUa+8uS8zk17YSim1cF0nP04k4kFH1thygwOr+hJFCn1yDPR6/4TYX8kspAHiRVo0PcULD7fuo
H0fbETEwmRkHbJtPGo+hoiXtK908pyTbZDGi96yDsiKbKTuTHNTjVLNkdImao7GrkiFwiXXDr9t5
+wTEiMScmYjeYPajBW0kuvS9hsCjF+bKme2fbDhJ6Ctnmfqwur4+1DK0WqMW/lAeRh74Pnmcgzmz
hMCMvQGo2SsrmLV/hdbXV/3Mok7hXV80bzdETrhi7zoXr7DEfKMpgyoVXm7j4upg/vg7yRUMG4+B
7AZinfxDMGNtnABPapD9zg3wB3ZoStY0F9N3ksJw/fc6aBoUe7HclFUGOhzjHkMAMJypyt59ZTnH
NzM82JF0WhoFcjec1aohPnBaXQgOWyfH+XHdWD9jE2jXqo7EJj46cTzgZwoomzzZ7aDRV7jlQVfI
h9kpg1eAGYxumJKUIO3HubIJjproNsfswo5rfzzVAEMwO7/6iR0w2WeES2lrC15GyYnVsioziWHE
C8wjJs8KtJCUraPsGbQiSYE3l6scWLZW+eRdcAZztCmF7/hJ4etNGlP4lmSKVDSfcjwrKWMuaNFf
l7ysF0dwOnQF1qqMK/dPGZobniPmlK+HRKNT4jbpTeHZ/2N66vEHvEAp0byDj7gXMyowyvUKBYB1
NEoZLyOEgMj5jh6wQWIeRYHcyvVBvvYiP2byxn61FRmAGVvyW60U3jdtW7kr5uWWms7uKNvSLfEl
XC5fobizdbHqOWoCsV47fX6foq8D0kXEp2cvehlfPX+ZNhPl8d2DKypY9Z2gxaYQJ4XW0OgKUuht
j8cE9l4XgmGHhM/Xb/pJxJwU1v18lebzAN2pPSe8eFEXm88BIp+MENMLNhEFjYRytGdIqyQnNIm/
Lrz8XJBY/SjZ8BET0syMDqCXEWXsR4nzypM5zBFUcNtUqd9PsQeLrM671u25zaVcLvM49nphiljo
dhYdUQC36cu+Nabx3+2L6YjuOURwfMxRmkzY6N4Zwe3FXz9gyNfOlp4U7nwyPALow89H6plPQMVu
Kc1MyAFfkuKG2a/QtuhWdi10zoSh2EKZJ04JlWQEhzLdcyhcKaGpTnJKaQP2EY5oBMv/HDw6unga
2/Xoz+mjIpcXrxjCJA6D5vQSJnXqf5x7th8x3W2tGuX9cjMc/PTutbajSi5kcVzpBbDwcOOkE0kg
khkYlfj0ciLnPCywWu6a96FMSqnMIsiPpX4CbgtYRzfmMQhD2gfsQZ/IR8BHxHg5GHTEdCNptbwG
pHNi/rcIamRz3SH5U287xx1FpC6qWTYhiT3Co+cHO5LP2bBBFcfOMkfoKkMunvQqGHK4p5oNeQr9
l1hFKo5UPbWJPup5s1RZPLWSLF9SpHYP+gaNDqpmr9FlaQwzg1XWGUH1En40pXs8fkluR/V8gsLk
fAeCLIrwhRr9/KG1ULGV87NjwwWBNtcZStoxnNIeq0F95Y0qurJRZ7zrhFVJQgNbg7tvMK5kXhqW
5yuGsCn9K01ywFrR8cgE/YJ8O0E/XVrSdVPweTmbbxqaS2YQs5WwsiM+yG7hJbw6W+C5qYXOkLV7
/30ZYDA2G01rXqEJeF9APEW6msGMdON6rOfibUnulB085M0Ii3u9+kpX8PKaUUkdY1MDWKhFy19Y
Fe80SUUfbxWNeRtdBIG4L5ii6DOyhxE9i4UKGlkiX44nMBnau+I76jDR0K/b7eW3gEW8IE3cPeJf
XDcbPLEBSM5NWO1vBuyvMqBoKFtYfIMbxColmYsM3ZhYcaS18zZguzxbLcKDg+d0fMPrzdbwjwtp
18JQKRSPnSyGNkR9o3xrlIsb8egan4zIv87ZgDg9GYrLNL671wNFmaK2hG3UO2AYhqSD9CTA+7VO
HdP2M/x7UstFS1csotOoxpHK8l51miZyiRrr+KjvWtXnXnsJQdVO5hLdfwGasqA0xJIDNeMkfoHd
Vc9tnFN5oKy+csbCetk5gYkQsXK+18C41SKkY4EwHhEVTK4JYmpSzZX9Xoj8ULcfbWCep316RmSc
keWpA6TxaUO0SbKOm/34fgv704BviSlDbfEZXXPjfO9nad1zrPKMYZFZ7ESTX86NiIG9tKr8ipeY
wWxQeehPDG9xkGLEqSzYdEftcSsYCCTyCLYJVOqD7sIRkjT4KxJndg6IwWHX65ceR0tCi8aHva0q
vDlpKCNcA217ifXddq0IGrzb5x1+pRAlDwM7tUglODccXl+iMKzHUSumSajavfK3FDmkqdme7CB2
l3cymOv8iZF2xJkz70jer5A+SV3oMzbq1zYEbS+vHRPs5eXxewh7o8bZaO/CEgFeORDK8Gg7gp6f
JAJ/itA8MXHTZFcViBheyqjfxkvxqCpBMvM6fqAAJjWxER6uJgTPLP6e156SxkSUnQm3rXoAgNVs
yjyovMBY63CeY184jeJoSxD1krH/p6s5y9t4s4OKvHWXtBdX1dArA8P+2PVLCSqfokNvZkGE3kj8
r73SecymcMNcqPQUF2aOCLke9MbQuxNfikaMaD/5u4N/HSqmU3acWYjB0Qz1oUS4attVR9xEWYAF
dswVyXGZaN+zTRZh0dm66RDhVwnufakMU8GsGUKCr32FXuGJyevTdcQI9U6OJZoXL9RJEfPGgm1K
OqHNahUSuFWteBeH65/ZW0cAwt+znjjQ7jawi2X4Cbf7GAlCypVA1ONVfZz61c9Wq1nd6qlUe21e
uXDEpV7tTV44jXMtBqu+K1pcgHllo89LgRJiJSYiZP2QX9pDf/eVeCScuhaUeqZGyzvFMigjMyr6
31iDrd8dBr+zqavIUTa4ZNa7mr7lXTsAK+Z9rQ4DLYJlOlZg96fVXYD1gDegnBlylsDjO4S+ttX4
y84gO/7t6tpy2l++rltzidgQvBfGqV27kXP3uOtNm4OXzFNyoXBzL+xSVJ3ZPDg08Evcqi9G2DtK
KZc+a1LsiTpzUx94w7kgk6pISnWTDnqIDFVU/egbrovu8mVN6H0wlGXyLPCrvtGjSZEpkWJq372F
wtIa2DGbJaSIyGjK8NX7OsuUV/qOiR/v8bt8VupW9rQWFG4bgcOWwCAlfODdyyZBBS/V3hFkDhAu
iKFbXuLLdxlozUi+NQHs2vIaqnZkzWIeJ4X+2c7MRu2IXiTuNswofVPqeX5rcCGYzJ+GjtdhbatT
b/Cvu8mJalxQjDkw+IzD861X9cdTO2pLWWpnR+l+NB21wqtGkpjM9+2uyPKk/Qm5bIL0tU5s+TlB
pVxe/5eIIfBOWTaQFJUSVAYrQpyIUbQ5sLChpFjVV9mdkeYTg8HCLtFA8yEmF6qucSvQrFagdk09
ST5A2GCeZCGpLL4QDaO8uvf9fD7oT0U9T43FJkWBm1iiPGafcBDmlf+MdRMJzFmGw059z1/f+Cyy
Ndr0iMnZVqsU6ytDPQJa4+85rVhW6Mk2VCq2RZJhveXgLFyij9lPbuJoC8bralQdS6XqXDzr9vDE
x2jybfhS/aGqOzw2J4VYOh45oRjmhs5IRbemGsPL+Z0SkVtVSjgRkcbRlan3stzFYCjR54Pr08Io
SjWj2kL9lBF49ikIlQrQRPjTQZaeZ0UiCXPMnIlZFQej8E+ypK/IBLSlyGCiWGCYQctW8naRu/vo
CxTxr0fhB3VbZoli4zOotWl0s04LCeiMZoT1bNU/3alApX3ZSCPQcGhcSIlWBHxjpmTclX2vXS87
6DA1QljlCZuOWpehpfz/FQK2uqHT3pShcTaN/mzFtB78qG87zRuSYtOUWo/xNZWcxzj2miivZq93
JoxjajX+uf0SyLo81hds4iEvJHXCS5HYwE0Ixu0chQpyQIt1ae0MWpPxnJoBJko3NN3L63Y4RunU
PoG85uRruJfrisVXZMn6lsvDyCHRQRW4byAqqc8uHW6fa1dyimDwBGAKsWwk5hV8O7sOnt2+zfNe
Qc6Daq2jgR1WcnB2yDLBIsiQsRCDaIl3fau0uXUlbqz4ZZo0QSlsmszcDcCjejl9bpHJ/QtPcCXg
Dl3vMP2dGSd5FtV2kf5JEav1SoMu1JxDkbIUV3EUCPluS8hTgvlcAs+Aykp2xtqRdb39lAfbEbTK
LXuexwrTnVPEoHWldHY+TyQfKW338VGq87ZDvFI2uVd7Ks5GX4A1bZnXJtr8W+g35mGLofG4X0XJ
nkA5pqC/wd4Wwy1SaSFZqwGcN/JgIce/M1umW8jYJRcF+g1hngUGhxORebCkl6v5x+cxWG6qvqEQ
ogmlKaBx8MNxldis+7vEOmWqGZ2dWTxAszMID8zCfaZmj9cgs5NNr+R61faiVKreqfzElq2RxL9j
xtDOxCss1B1c8oEjxsT0WuDB8mZ80Ix3OTOyY0bBdmadEsc/pRF5BlNov8QZlMJ5zmhythBYd5Oz
3NB6rN5heY5X2BXbBGM1i+GB5BSOMECGogeSwk1/hlaWRWljqqG4i/pyHrrSzzivb7Vly9fHWj9L
+AV2KOoYGDWf+aDYaXOVnAXwJPoiAaHYfGatH+LdvIslO1n7IRJuicnb0tskU6LRlRjewFRD6C9e
bIJGhoc2AKRJBD5mw3C8wUTFupFasE59dqRUUCigoXDrRozcGxxHkypgQtZpXOF3nFIcZ10Re8zX
WjTKTcIAeWkYui7XTgfnzJK6aVZ/rXfr8ULXOEQ2D+ManU3GUJCHNIqJfTyapzAOlr65caddO7gu
VJX1Y1PMKB64B+2d7x2KMhyo8RWCRbirATT7wE8i1HFUeWBI+eVlIS+7N7qwEawjHT4m3f/6Tf8S
+3f+GAcIj4FeIVGDaBv4bi4RhK6sUCZmrdwudCWcxlipzDv/3V7FFD6S4xX/ciBtePnK6Z9bNFYo
w+1sKBh7kAANoIGw6siB00E36yteRX/zmv7rBAWkV+WsVgHb/zcbUp6U+SWwzk+OiiEK7crc5glC
pWS+C8lzCVotr1cEpmGsBaY1FT9JYOLPTBgXTwgI4/dQYBtoQxXleBO8LjPh4I2G6s+JE+8uJWxk
iZumz8CHHeKDIMX5KiIfrgFq6MJcBv4i7KJWB23COebcym541lrcrB8l+3AxRyalKbH/iYmWbRHw
gS+Kp3GbAgaxXpMIaBXj1K87tJmDVOgH1JoLVWydVloS6MM7WDVXb1pqx2c9jYWAnGTlaf6DgXo9
pByMQ5dJKSHWdXHr82PTcehzMzx9j5V57wDlP7m8oQeoJXfFASqBjog5hcc+G2ACvy7hRGrqdjvd
UbIXABz4RE9pcXrhFUxiUYBy4XFb8ZqKKunhk3HlvO82S5DUZ3NLImToAqEhWlR4GX7qy08pOcpZ
z/dgi8+r9QC9LZf/ejbOfDZKNU/3AsRBcdzSk37Ztv4MgZ6gNlhmlpt1EHVmbBurribRy2E82J60
lnRtYPKfN8I8a+sIVIvOxlsSwdRnOTeEftLBih8SGzk5LxpgVWtFmDIYOtE/Jtz5rl3oQXz8FL+o
GzHH4H2ytMdoxxwWt8DPk9dJ3JS1MLXdCFr+lNykUgJhfWci9l51ySN8BS9R0AeV4p3Uiep7KtBQ
KqrwuQcXjsVVoo+z/XDq2bvfzZ7s/aGQwYb5nk2bSHGZC6S5c58ZsMfK5BjZd0nfExYyDHKy6ll3
nyYVYd0eJHo4l0UCdJ4Oa+B/mPaELKOFmFZN9ZJIa3NYr++HwAqpT6PiwIVWLxHBYErikONX34bZ
/1oWZ2/WEfFG2Ii5j4TNsHov7XyqeDViBgaKIB+uYdo20Q+4oq1tndScDavP9wGKP36pL0fMUuGD
+vzEaXtZehOnO49UQB8AXpIAG6b26YxZgDw1Qmrrpha7CjUnRgDG8awDU1kxyLZV7dLcMmmUUSSo
0wRRx1+9zbomhGHuHV2HCSADDQ8XrrB6I47NMjWca65QtAKDCFfjaUpvwwI4TAQnVTuvcPeC8q2k
FsYYU9Dvcu1Tk36e3FKYCfB99mdPl2cIPnvrgJ0rafyKJiFobtMqs0tA7YSlSEQB+EBjSrctVMJJ
oJdANiCqKdunpED/MJxAp4PqqxFpZFLRvkmXU4g60DKFEkG16oNHgXQM6jT8Q0HS+NiPry1qsVjs
UDKA1uyO58WNyg6BBx1kHcM07UUAKyizlG1Wp9kdHja/4Ey+esLtpbCIrD4bIjGIKF3Bx0atmCHB
fWJFpw9B7zEUQQmfbDn1N+y+DD/QBiuBvm2r/KeIEQ1up58VFh+fmEThY4/EpYd2Sb2xeKb+oOsH
VCtnzXMhn6oGYQwXYztulj1r/YTsJ0btE5gd8ZnH/0JiwrH6zZNRibGjU6fKS5L1p+GMQi+0GpNs
JWBm1R3jOFQFO47wNUszLwXcPjh2cRVoO/iievwcKdO8OyjI3G9AD4DMMAtx/2KfzBKU3/QT8Iz4
aKwyToSYbjotEoMYZ32Ud+wc0MChUNs6NuCaM70okJZ+ot3NnsX1TzYwlssVmeulgdyx45B+spVZ
GxJgajfo3jvGQWODR59MmFz0ew05oQ9S+kmMUK1i3j/KQqwZdgrrYaB9bjGwxvfLrYK8GHjq4MIU
VvZiPkwRZSygsour2RGCD64Gh29eBj+kYVimOYvmnHYAwubtFovX8yiOTbFmw0ZI1O3zZjzJRefb
CQwGrMZtW/2NJGAaeksai1iFGVxsf755rPspUQOKdKWSw62D3uyUcqIDzYEuNcl/uFxko5ETxGPc
85vzvDc3rVvZNVw+WY9CExB2Z2nh9QuobaD+G6U1RDLAI2h3OBjh6CxcE2GrEp3AieI1l5oZl7yS
+rPnZ0rej4KOJ0mHsjtu7fmIpwZNRToYbVcAUXYEAR1fbMeXnrpof1kcOuGtHpblOV74O7YEPHiL
fOSvZ+7OTkGOQxVP2OLw2vDyvca6uQCb8KaBiPYy9zxncQSzuIQP3xrl7PUWurSHiahYQfx8cWyA
1DPiEbSF1Fp/oqbaCl33ErSRXtsDTT2Izk2IUKD4VhAZF/kuBuuAvtYUaXR3C1GVDHDDvfqLnupL
Cu3nJhZMXCxPc02msy3a14XV3a/cmP2/BjZaG59CSQvTN5VGpAVhxwl8Z5BLYYgeLbQ1eZmeZQN1
NxTS4M2xY+fWu5F9Bql/WCI0LAJLMo9XO7zpAWPtt3lHCxjka3wNqa2IpHHsXqwHIy+3Mb1N2wrY
lfz743HNXz6zqK8gtA0XOkizWSnO8X6bC0YwFLAHskONMBxVighVxrK5s3OMM2LNE/K5Rn0Z2hO4
QeG9TL7UEJ20Zdzccj6ZWr1LyD5D/1WM1AdsL0V1ZTrx0LITdzqtEwoRLBJ4yUogjOdiTEGqvKYx
RNHSQUIFwr890xA2qczIJnjXETPqi8cosHRLeEgPAHmiPIIZK3n56jV2X0AQvzYCtE/Ji8aZbDVm
cmHJHsloPE1vR2FwkPbdGQGlj8KYKoBWBh8raG/5/X9f1WkNnx0zvHAQXzLCn8zfc9zhYlrucLjz
hOzXfNPSStcG/8WwsD6c2XY8d/a4nvVmr1UZk86bgHEWPaLHSvK8JEBHj1cVoMchdRp2wq0jMuyv
rfCX2FGu7BQr8go98muLSJwdAA82e+i4yFA+n1BXVJqCryhzumr59faHPVr3x2Deda6i1HZgO1o3
sUiUgTvUiy0OqXLpVsy2hf7wnmY11nCBTeg+3IkYqYwbOkRNmbaUcxZXRuMgEwIA//dCT0/8DI9h
z2TQjJGS0sDNx9MdjcBfFqmUA7jdXbmXxX2dQM9SLU7g4tE1Zb3bhavS/cRvuAmJtHayd3II2+tU
gGYTU5Hx1DSysMdedk59xQUAaKJ4rQh8d1GG/t9iv90YLT1/HlOHNA+44vIsVD0PYcA5JkmX+ATs
emBvV3BvFA/NRRnsm1cD9hh5Uu2DYqoY811GAcrP5AOJvILGl/rrJ6V5ZeZ4gxOuS5+3H/yYVptI
m8FugosHQToNffPvpGWGASQBoCw+qz0i+VBDWyQ3RxX75I36eLJxpkDTpE4URgYhaNugp+aGH5xy
v2tUugcVKkrpZaHGS+NEItLJnmAsxSgeZya3XZGayb3BNv17BNI+7CHUI0xV3I1wacpL5dvD5LFq
z40eZ3BPekAOWdRi+yuV3nzZMaQQVwaBfccRsnhjAAblfdjaPPKVzdldMGSGOELnHnj8wz2ED/H/
kPg7sk5ulmwQO9gZ3k+uJ0BvXnurYpQfZB/eGDr4PbfIOeddahHXAq4zU+1NcvWYbbC/togag/b5
5aTMtugeB+CN+UtJNrC/XD3VnuAbO5xXQF6Arb474bkK3t6zY1N6t4lJcDzBTDu0qZCyFS6VnNM4
iYu0D7VwEmF4q+ziIPvYUIo7Gq3NVNg45cvdg+PY19P8Hjf3/JY+E4XRZ8EYSzTJyhN0SJjBugzz
19zMtR3/7ywsERSLYy+E2hpVsi4gmiwpwUvL/Qqq8HqNj2mgWB3XpVI9qrXHBG6stflFnymARIZi
yFXQagf4mFldnrEz0bIK3Jur5cJDejUAz1NObSM/nyxGaGFOwuAxQOLNB+yVpUR5JBz6y7b6XANg
KZFyX0Z3wscASRGNiGajNvezPL9g3xzGx/iort4FU8T9GknkGpYln+xD79A3FLe/Ph7mgrdD542r
NdQZHmHYB9IU0nhmxNhuWgYrGW2kf4lcRiKjrXJhdKBZqou8Un+DQMa5UlzUuurICS8C3VQuEP97
NlGkXCLfo/j9ZPKWT8WDL6pRwfyamdEQ+KWTxegEE6i++6qjXKQHcfOnP6MJEZPO4+icI65EePBz
Clbd4EPtBKGf2OykW9sPf18MoQ1rznNDhobVRYrdiGxr2H3DxTBzcW8Et2rQX/vYz+8iHkfSZndT
SJjLNydOXe8Q+fWvfekMOSKYEx2RGWsuXANhm48o1aNtipk8hTCoyti1Io382xpc4WGbq/S9zJdH
jLLd+BQcTwt9tqnJzmHa/9x2GXLQnOZF5SygGHxxu6826Dz5b1JLYEC3Kj73nS5gkbNGLCz4fFyN
4ANS1aGJY2BbCLGC2XgNundLLgGaHpxcGaVSP3h8JLoTtGC9Wk4Zq3F61nCCGXdz/CpRe91hkUEl
XET4/1nRF39MwcU7GcC5K9Mqa2vJfyOAFwldu/TxvIGBw0zvOD0b4iOIoZLqdmw3svxYW3xBksU2
YEJthAZuO8lKkjsqDDsOdlbyZDKqbgECEgOVPwXdD93jma7HFSAQCTLz66uxysMrX4uFGO7ew9zD
ehEj/rA6pL8ho430erNxgk9CHciGCVefSjkSbq0p56U8AKOARdwxMqIfXdx4M8NcFxQAV9ruxx1t
NZW1VciqIiJOtUeAtE2NNvi85wWHHeryIbd5JGnpo5QXQbrsCMDJe2uCfJ8SgxT/tvXC+8KHYSfk
aiVT/ww+AXxcgcUwVruGA4Fp4zud2YVTX1qVEnKdk3nMtCpP/qc1sBi4daTdTvP9hsiVMW1wqusM
9LlRW4c4gN2PvUimbMy3JXWxCE2rEwABXBXkTrBnruNz3zitpRlxxKAZU7iTYt/Pfa7MrURGLckh
f7KlUwK96GhWHF9LyltHPdFfRiMljcVpNDBcsZ/zUL+ozSisddwJiYat5ZAhy1CKuVrxWGM0iWwV
yei5tl0qWwcPM+UeMgv7MmQhUg6dRw+XoANC21BkQ8F3+Zolp4zzgNN2hGK0rwwApjSY2xwRxpwh
PJ528E96qhXLoAyOxXPNGk/cOCTsht37eylw0jV3OyF13KSPCMKHYTJPapTskmahk8vXO0FcrCmO
re6M2S22hdyblPy6lthW20vE6cijlfvCUZlfpxD51wvjq8H4qq4Tff4UzsX8QPIs09vvaptnPU4d
e2tVkGPqKDlMeydxXl7NQsoWQ+JxJ4s7H7i/VDwa/VcnlA632B8sP95PNhyuzY0xQ/m0VujMpiHj
HXs4aNjCkz+Fi1Y4n3toSKebc6ASxUrL5lbkhutGse75t/R1tXoFxOrCbSadAMg+GQGCekVahYPw
chEpJHfGeNBJtcGfQos1a89dDjmI9XIrxD14HxA5zHQlhp5wx2LW+PRYqEPI3XFO5d/otbIWX4hc
mvr2wwOUYyUmbxIsXLwdqfGDgYxgn3axDYU8dnOcP0d/tn964/a+mjwCKcT1ZYKiTBKjoG0rmsVv
4ohuL7vcyd4jZCYoUMtLU9D1aix67bhJEg5rhSkQ40RyNbedSxajWG6HYqNID2jOOLeUgwWNVvdv
42Zgy7ssP3MXoZrgnPqbNSbrin3cZpMVw+gOhlJjVb92wyWUoUiyZRtis01LdiULly+7XAGNWL4J
pEfQJui79IiP9cAd7n56H0KQ66xCWDWcphAoqhvU7v86q6dZf1JwrAawkD9LtHc40pl2GlbvAuow
JYkyBQlbvwKDHfz77Lh0mFuTJ2P8jkBCogffG9TS0V3D22jJelYyhAzx7ciEn+KyIY/WtKo2AlGr
6peSpW/sCuSiob1yiBzepoGcqCLGR4JQ3B9U4kjKc4RRVOw64pXGy4Cte2b7CMRS5GBUIAcDZbEr
xYObDegZQI7FlgyczLj0LXJAnF/1IUmV68LfnTrUjCVa197GtxO7qVlEjiUtaEom4gCx+oIG+etK
5cvGC+mzb3m8vDL/2ugDVCGxWjI6xoSqzR//NJYkTaA6wYSGZUbjGrPPU/uF0e17L5mGUU6OZjnM
048Mthx6Q+VWAa5lcFWq+hOFCc9ReQ9M632c2DLDujeUSqY4NL1oC5NHB+65ywcy2Tzs0HSvWSL0
fmCE2oyCEIVp/tDjnkSzKf7ir3OYOgpBkHtlTjcsiGwBy/kSwuWwoOM41p81c3MTZBEaCp2d6BDa
93UvRlsv7Uo4JB2k/jez7kFkIK26D8hB9p1BfsOGoGIPUQbbsmK28rZ6l7T6OkYw0nakN0SDa3DY
VuG0X7oGQ8tbh6JgRZmcgRb0I1kK4CvieS67JJGd7PYwYls0plbz5IXK3irLijxRDMQUB07zCe8j
pdvTQ64wxgVjffkba+ZEs8MK2ztPwGbqdVoQqf61uE3UgixiN4+k73yoSkBJQ7jms/recVZdN/f7
swvHWfyEqg0utY6XNk7TDu41ViZetGwJjjQFlNDyBC0S89y5uBuQCNoggsJx7/vxL6ZqkHQLeXGw
PhRCPFfqLmpOHcO6LOk5z8Kc9VflH3r2+Veac7CQRvcFkhKwvz8UJVOuMfgcj3L4G748YnZTUjo0
pMX9Hp8QqN9fxHWMJhs+iYPHEUghdHGRb4Z7Tkm+DO6uUylZMsN/6RhJ2ADhTEGOE4ptcv8WQolG
t7ihyGdvBWzxbHX2iIrQybCcTSKH+jSdcrFc1ableIDjWqwwKLZEJsoL7/uudQSTy0xggPHW0vbg
1ndjFnyfmYM0nWgWUXXFVM943v1FHzmyaBNn9jRWvEavNfnzct6uJa0oYZycFxhAR87OlKw/KoPV
+io9rCLn4L2SI8DtZQeARD5Ad8xoBxSBwjTLZWYvioouTWLZjBgGm+9TyBWEswi1WyXJIPzhNdvt
FZxi3gIbmb+qyltpXsbHMwmrDOeP+V459gDNqYYrGzwYEsUQUZuzAtN5+Wv+0lwh/YMdw3ZDJTFa
NsQudW2v7theeNFiOnLlP6mJIs1AGMOMazZfHR7K33LoLN+2CQ33Ga6mBNvRHyavYInUYB50oYBy
wsvHYx0bO3aaJJtBOvV8QtDhX/Qp1JXBDOBK8GBm7vRu4x+5c9OTHiqPPD68bxKQoNBDR+3OQQob
juSQoCiaZGD5QqJdL3FeCwc4bVZVv/2CfEw/FWe4OmGbwn1OfYkYhkJYmtmz1MXRS5EaszNcNXP0
wnbw7Q+7uvcLTjcc+mXAJYyWTUtb0hrUUQzS1OZRr87OAKQK1q0gTkE2I8tD0Szlt1YfOVPZs0lW
X4mQeattY8IW5cW/wfbOhVTSWFE/XPLkDx7ZP4TVbjniYlHl3eBsq6hSuBK9ANoXmbTPAhy7rX/r
NyzWO6H3I4zy/t9TqA/C9waRq4RqsnmIN9jvzRdkFcYW4BGj4I3ZGw1wp+dctsLJbloSvERrSfaY
xwJSQZTkKA1qG7GE2SjQwZzPkhPKvLrk4/V1E40UaSkqVlJUeQnLBXGRsR+/Hou0nQvHQOEZYO2X
jBGspkgomkeqfdpqsJVWWlaGjrpeqv1dtaFBh+JqfZ0zljEyxZXL/1B6WO2H/p213L8v0UXd7CYW
oaXheyBXiThTs5XpvxDC5sm8iyIzYvQfLmsYwoG0YOCKldwfjcsTIiFy/F1vV8WrMweObSNlnUZh
Ok1zHOoz0d6qVheVhv+J3MFicvvMvYWDF0NKQ0ZDJtCn/61PkA11I4bzXfUeRj1EKfXCChsMLBWA
g2287yg3Q/HPvmh0xImvmgewMieuss2FcoETtY/gKqjrJWjAY3x/EdbyEbU9FbXi/QN77lz+ko6y
1dmR7SXinXe7whtRxvhiqfSdUMrXyBTjY7TVsS7P/0Ib7uXcnHla2Jd4XvdvNSvAgSX8kXBogNqp
oo67soDhdINkVqTjSkgdCOFxe9/85Z1b1Nt2gHSjmnzh+L/Rs0B2sFY+5ib4c+SGsFdPEXz9B3oE
ZscboP+tccORo5YZ6WG5+oJ6/a5BohTcdmxiYAx3Bkydi0bzMWWaKX8uZe3rDtIs4FmAHmVHukT3
hJ+Nvj1aHUI5EC47XxQ1kjMBTbTBX6juTW7+ScoSELaWlrFd+G+LJdHMwO2mAHZeyppdTXnbTYiF
7zuffjlCIOiM4Tu4YLTq3uoulFbm8VyZa0eWrGp+DzJfK81vOpaCElno4IZuAnmG51h7mAF2P/nt
Zr43kzgGMikZ8FUe2r6TJT5XjeG5MogD21UiY1AF4L6mex9b7DeK9NxQTHIiX82Ys3JHWag3UXg5
QfRsXeAMpHC1BQIgYKuEGg90za5Gk7qi9MkjXcTDH1Vf+//2xguNdzV8ZZqHdkEYm2WdeCQgGIEL
tUpZjQIBQDKFNjktscQVU9bpcKTVJgcWpJB1qNLpYpDoC73UlDidUmk6v7FLJEWaPq0gkFkCENHR
lsDQJ27kXyruZ5ooCFEOFrOoUFCTNdM85xhaTn1ljEf+djFGTbOfV1vwqlJ0+euSdLWaIdTW4hj8
/tE/0yMrsyb3PZuFXOmyJxrplWMrzccO9dfQP0x0vlhfhp8ekNQIn5vbdLFbmAUIrT6bvEw4JsWx
aWAnN/QapkzPbiEM55vh2K0no1KLcuxW3xH2kviCIxiekVS4I8eYVgPIoPpKxQypmoAmWg5BsI70
FOrv4hhF8z2qaGnI6pw3tAWC9EeXIviswU3FVF52VUS3Ot5Ut1oH9QEPCjx1W/oCli9H8ewfP8bE
BYGsrIQMOKhxKWFffaDEE3tZfBEs7z7nB1cDZtq+ujHO8mY5T22LdUI/ZriH7SjPoe9/duNvNibo
Ae3ep2bGPRflPx8UOquElyBBe8fYWFxehrxjY7YkaHzBPBzq9frwgvxuxa4cEtedb38MD2jRuKiI
CU7iWNa0DzHNJPPT1paZ2vAommG7on5kFDl8XOnzTTKJcFGXA+Vhqxv0P8YUBKMHtlPD4gmIdkXU
QW4Hhd4A5pWgLkMrJDE5WXtb8a56OjaloOkGtzeA0Gl80KS0IblmUzQmR8+LfnFLl+RPUxcltNpn
xF7+JM2waVKZM3/KhejH3X/LmgQQD1aD/brlP6D+8d3TH93Dryyb+ZpRO03kaRnoQOAWTzKvpiZi
ggVOM7ruf6nIGg6NkLDt1JOoSyxEbPKUMX/PAyyQ1teCUIJIDNXWXsPDtguNYkaxYdJ04CiMPnR7
lbibGS89ETB/+JtFqYwaUZFFWzvp9B7vCVzUGMS5xtsSxzQimFzR49cviPNh+woMod9iwea33Dji
HngYeEhAnkguyjVLRWovHXO3AAQ0IHZsHWwbqlWkMCVlwLda4AOXjaAGuAwPLHUZJ+/Owd0w3uXr
p2g0hPEPOH0fABWxXl3XGDQhwPTr/rjeiEsFqwewt8I5V6JNDnamuGFzfTlRigGpqdrJ5KdzOE2T
dkuwMohE6xZeA+D06En2RbF9scGPEK97FJklW1VUZHsNx9ZcGGwknRFU+FLpJOJUJtQDQWxIxfpW
JaCEX04ajxz/iZJEF9QB5/t4fVRL3cfPEo3A+SP5Gfq/t2N90hJ9qu+6QFjYd8U9tlcwJgNcYvau
Ohiy9W7SRc9r8l5n3lyx1++OoSBkyft6Hh+8rGJb7iZAl+3TTG+jLHXOwKuLiH6adwM70ohFhkIL
xuCEW7YawZtUKny2aQuCFzpC0jo47CLn+t954KpVhagqKdmCuQDSnvzePhQqzTedxB/cegOAR+1I
6yOB3vb9BMCoFUZksioJOc4peN0cLpL1yiHKousr4deIXt6MADaYn+2hNBuzI5a2AR/UWK8bH65i
BhqWELY36HZ9/aMPmNNt12DBVydfeFxaAjPeOTxktr1pUwJ5uRPyfzwUpj9bxK16Roca5f/PquyO
035xlo2hf5BNCteddL6+lmqc1HfW56t+BUssIoYqxMkd0mZujN3NvM5sqFKfCWxoFcHxVcP57CQT
A7f41ACnddUxeT1uEWtC83ZMbOlWSNmaicSkM+vlEaTgjUd1J7TFd2dYHG6tAyibUTxvvkjT4gdh
xRh3JyaRPbbM6pxdQMadlIr0KrF+t2nSY+q1d4y86zdk51TgU9pFDknrR0RGb8UBqbehIHKBxOZk
OpK6EWq0bWqU9O4ss7xRwlxnWQtRlytPHhjB1mSYfSknPvxSdTAD1FeB696xnZivzHGtgokgXwNQ
xoEUBcyyGF/jxlmOoJTuHkYy1Zjnx5wtFwnvWssBMK1TjxniYHPYQd/K3dN3VzXI4M/RjjZhxWrn
URDM36Pgzmq51S2M/DGKiFsoGck5p/Y+T1v8lpy8ocd6JXh/09YwBC/7LASMmP56rHsZvwYfZYGV
f7XtBwFN0zkRmlolqwYF3skks1m5hPBsYVmhkW0C3yXJrZ+KrnMf1h9dIFMDnmlky0QqG6vyZl8o
q8AMMsKz1vL59Ir2g9eZp78HsyRr4/m3yp0uspitN7YFjfDlRVoAk6nVfe6BSDwSvir5MfrECHIh
g5ir2tx978qSJ+jqRFRSj8RqLmVdEMOM9lFQNjyb5Wwgr3/lS4TYjM+JkwssYbZL6ylOIXy5IJTM
QLNEuG0fnvZdeBhDs49v6ShMBt8iHOZ0V2kdF9nXhk4d5KbMvzFrstDBpDrqFqSO+Ltar3iQweDP
RTi8o8OfUGIDPTDte5HWTexpFYBVJEiz323QaSoCrqNFcecUWcGpbRMgH4Xm8vYLWP4DUu+ShKbp
rkiXjD9AaC4fOMZuy+Zt997z/EV6HvKfNMVLgTvS9sX8Yd8UAueSG8KuVNsEVpJAaqYaAJhGgU86
9VHK/QORjr0yQEgCEVSwq+dAr39h6wj/2rO2yILaDX+ibutn6WE+j87aMG/h52pd+jsqGm2ASnFI
xED/jbz/RtcXjuPBQjCOqp52/1dmeHtjeGUgzrEod3f+iGaNK1iu7vfqwGP/h09MfbEPVDV9NLji
FpGIGpbLOrDzPbq/yx0KmWJX6LrLkR9CqVqnY1wc12mF+1mozsbTM91GI3W0zM7G/5qmRhJg3U5/
LATn7VgndXqsy4eBK1mjM74mbZF2iU8HxeySzrkmdSU/6okhGidr/w8aFlYIGpleYv4WZFmSt62+
ob1gt07LIocfWpAZu5q9hyxNUivDMMm6Don99NpCxgLCnjrvUEwhBN78SGbgD0NQU4W2nQyaUFhP
DUwfnOZpRRE28sIcRly3WaaUyFgVfTrfdNWkvuvwqOrd1WkkkeoDC6hTpQ7b3ZPhNUL2gXxX7GX/
5joP5R7clSpgSWEkhK0xt5lfgDiu6McMkuPW2eM3UaUnI3GrsOhhYOe4Kkpnjfczhhdq9Kp9I+Y+
fXx6TZwGbUak1eAwxUsRlO2RhjSs7Dzgye+EY0Y4VARXGANNodbigcYnLNUk7G9H02GbsxWdLS5p
rD8YpoT2HhYU2Ck+T5CGv+GHu5cMmhfn+x8bZFz+hUkiQWhvxF6zTbLdGp04ZvogokO5ZdWjagep
LUPgrk8sCc8hRydwGX4i1Md50cCL78a9XgUwkuG3XIefXhznPBu0S/9+PzqssZa9BuMAf4qlLF+1
prXpYaIpQkGUw9vWm7FKo+F/Qme0z8JRVgLKnjbmUATnTWx6T85ZPPm19ArnpaFNMDG6nLQe2rdQ
oMl4t3mhXe1pRXLo8UKAOoNoH9wrZ27OR0OgOCJMVYJlBl3bRbIoN9j/CYtoZ6wkmlXjxez2026A
c87DJwhGi8gtG6+WsIbW6P+UmI5uGrY++HKKMs4dsU3PHrAJSfFyXMeWF07hGoPzebXTIBS0e1TD
0C7B09IktfFFNceEJ4IxZ6iT1jhpVVDmWFonEHxxih46MxTYwi3JDYq9GyjV943oqLmBUc+tTGUM
L86aQJEp4dLX0/837cqRzd4s2nY6dz87VD5ZfI4ZBJSWjjL3ZfBxV646aK3COtXr56i0EMvqvT2F
f3cDmskvbFB3DTFcuVCIoI+0vZZbK8/sFTPbctq87vqdUezNaqqkIXBIv1YikIWE1AxCFdlgXi7o
DmLKJ+11uuu5Clab19Tg82lRD0hFocAjx7jWShANkdt22Rd1Q5D0Ha02l5037lVjc6wMKKL0ftZq
grJVNig9rV4KVKBAk7qvL3p1UjEidZyeNiofBX+9okSzKNODEvCnNvJ7PLP6F8Z2h1pVfrYF7D01
waU1Rmum/P1FeMWHXqfRRn3eoRrUkz38eFnLiXIQdCoMMv5wxxj55YQd4q2fNo5XnR8hA39L6gAU
KsH3lzlDz9RPztKfYqI173mEjezdlE/HdwmagLNldKyU7+eVJeXKE+RPI45hCLiVYxWrVGvCgjWA
C02QmHDO/D3jq2OP8gI3oTC/X5MzI08aWsdkt9dVJUTJEb+5b9ZWM0K4BTRF6dWWTpbUecJobHN3
2XnuktuR/tUlEGLZgg8HgdrhHCYnzsaW4F8utbb/VO6zr5DRG9NYcRSBkYeavzxxnBMNY+sagHYx
k5SWQ6hktm6cecjx/82bYVslbOwLStVPE8/mAUbA+Z8tI/x5KyWBycr0MOy3h3x18TtlrfAHCdR8
7Un1ZlkkvKtNXW16R7loQpc/tyyjJ6cqp0+n9F20/ZJ+Nj7f7WLZlbpOktmmGBWl8WVmlFGG1P/F
o8HQsfvNFY6gzgp385pl7Co6Vf6HNTQKctcWoAAirMHGgUCqYwE3jyRdU1rm8u0T90OhrvwdOBr7
7kp4FqXbKbajMz8qY6fvACbc0Nvw4iL2NMF247Wkb10AVpwt4AWbciQiGdSI3V6JpPOdwjRbV0o5
xxFJBwaFXptDILW6Qo8RB4OMTjqpXf22Ffw3vZb7cq+m5OqkTcWEovOAV2jWeCc9aXek9WiVvNV6
S3FlG2+aaFpL6H7oj0JF0d9rifki0daVou7SDXX8I1pbfP5vRkNqlfj1pnPHD2E1TYh3yeylgF+g
Hvu5EY/8X5yR3E+Wvj2Ie8zrhvU47+cuR9h1/2CIdjElK870LcX7dEmh6RO7dN2837GWjHP6b+YI
nGxkYOAMlYQEwpLsYgiEW0zgVujMm6RYbgtwymbD3PlMBuI10TyEo00l7V4PLthqndUPqA4sb2nD
I1zTgzWPlTktUcxbWGEPf6AHMO4+S9B7P1R8WJoWt2e7OSg3Jta03IyYWcRoCJtBMLCGdrLTwNRu
u6eWyAsHExG6Dry22cl6bbJ/7+MSUHqeRynU7UdM5SquutsFGafrsvAoBSPeB3gdNAFTio2BUh/h
r3PwFHGpRFcRXFSXG4Z8D1e+Lm2XyjUCmS1UMpeEVhygLlqvKfIHW2Lu1CLZltkjJccUOY4mDf7r
98bfIWZF+KguwNy7Xkqku1qqJ0eq9wYtP5jxwq03vXVi0Nod2r5Ju7Jba+mqV7eYRACr9x+BtG7T
vYjhJM6qZ9ZVZ0qxl2YWWV95r5HyApoJ/4lsnFZ3ImlMwmdRidbWeMAIMAkQhPiyTjxkidRY/7Do
tKA66cx/9wAXNvqgFz+XFxRTd8j5mLCXYE5xWAchRV9Kz/yYUR9iEhbV0h/tZM9AnE3qFmW/Ow2/
gNvqzJNqQdXSdhO3GqVMTuosk/tes8tkLnnOitLB0kOp3EJYN2GfxMv6JFdUfx0KHc9CNPT0Q4ei
MFnYfhArqpuvlplgioQAYlJHeJVpNn5Rh4yJUE0oauHb1AwoipP1UORuE+mOoK5o38LvCwBML/D2
vtw7Y91EDFLIkSoMI+IEOj252zH1Grx7ZOKmbuiqvVUPIlDQhso2mVuRbRYTffAqrVaqxuoWMoU9
f5WFVoVFrQIs+NIlzKUtNJcZ6jpHIMIMYUQAJ782DgUmHuNLuZ1nnw/iITaXhV3cvivI+lh88li3
th1tyIQvnqEks+nlh81X0rbriu0WC/jKIP67NW+lmzPQykwYzNhb8jJz8fKJszKwOu7NIiVQKagl
9Pq+iroZTAttP2WthXfDzZSSHEGeGWNANz5yG3X9PCx+5ywPfqeOKddYHoHCdcqVqUD1+AJ4PKZI
qlZ/E4x5aWbagYnlxJv/AUabY3x3yepk2VhEAnERm+uGy+lrr6RH5OWhriG9mquFRwNFdUk3u8s4
S6m0bt/6qlxxQZRu4+hhcwRitlimJzd4VCbH/aKNvoF/wT6OkvamurFfOEWYLb4LsUGE6JW8lNcv
PbhS/f1Y2QmQ2iMAnVcGhc9bMBdNND10lhrhMM/h5O10Ow/Jw2kadQueCLRL/6pcNhcR3x1eLSo2
h1KI6aTyTrkqbe7pVvm8dnQ9VR2hCtgxKQ8ihOqxJxi+xtx0Z6oYgAltTmT8SYcuhqxbX2vQ6wz/
8C+AaCK42DmuB9fT6GbZAgLtbYCmeubhIJjey5hjipFYt+aY9AORmXCNUKqZoh/R22wnq7La8V2d
5UnBx+7x+mCcF8oTLYj8cAoPJz7pch/Exond0966ZLx81N/MwxzrJ1iQ2xj8t+qQgVwmegtlCZ45
zYf3U2pY1wel/sYaDKspyFNRAmkWbN6kmp1WtGy4xvtIvvXZcx6Sty9IK472mMy6ZTKDTbLgCjYc
M5XAR4PBIMyFta29GcM3e/NYlklVBOCebl+eFTn1PUJGkgfc6r3BuvPdwqfzsHsB9TxGCYVhOZXZ
CKi6kv4IbC37AVaydq45ErNd0+kn48WvVt6QXWPD83uWEyqnuW1krzY6xFmZ3tjSc9cLmylod0lI
Y9pzx0xpccKbCQlxoRgW600n74LEehKAdBzTjk+zXlDrri1giqesYx9q+p4QwKEJN7Nae1K7aCYC
sZBCf9lZ+vn+/cLxAAhbCWv5UGIor95bL20OO7chgrBmwIGinyFf3sLaM67R2ZA+C9yCLQC1CYQ/
rg8DHHc4JZUcYaDoaebgwK/cm02zmHSAtSnSfQIgcCbYkvPFP7eO45ZOgR/DHLzMA9yEKflP7b0J
JdS0wwCKQmjxESfH7/W6cz0sRU02geTBqp3hgLsP+e1s0E6tBuDam7SNUlIfp77B9bRNdTRDG5fv
Zh1GZTzTJoKpC+BgHT8ubQLK/bXSWv1j674MRSBXnmu8G8Mug2ZitMJ8pwmxhmGOh1vWXIBQoffU
u6W7/sHxijVl1dIUQq1Tk1IlGZaac4dxKUFwWBNRSNkPdiGADc/pUERiF5i/OuVHiRAbUPu6VK2k
eFSdd+A+3UOTCo/2Ywten8/fBuWdSfvsJSpXBd64Kyh8iEkaJj3QTx5EsZW8N/2hhlnaSku0nTT6
KVM2yKJektQeL43s0QbIXJKxX5Zm0VMT9WBureGvLvjU6vLz/PBY3NAuec2A/Zw/Gx3qWFbm8Ex3
nE8PRfNNFKnpTCEGi/Rz9lYPQKviIPjaqIs570fLYKmKeXUTn60mnNsD2HJzZgWkwOFBjR0BeZeS
uRvfsVbB2+ziZfw+GZ6YuoE8f7ej0+jjb2kIpw2L3ypU0RkSJW6N4qyU4XSZS/4nek56nXUyUPl9
W6uehATz/7A6Ue9wcVOfs4uhVWLVzlv6IxNBuccEKokcdUB/puchMopg/HpSHFfe5kXp/rxrafoU
TtJgHjNP3BpHSk3WFBuY9e5qYbA5fhH0aszhOg/Ph/IJz0xj8jMTt/Sc0JqXYysS+Z42nYqKtqH/
o9GehX1jcPV1mTsh6+oa6CbGBpkKgY7FaBh40x/Q4LEKlaWEzMw3lQFTHPgVQxLnm3GhM9W194se
AQe4Mpo0GULEqLVjYHHgzGUgn4MJZmk23NVxe393VCYzp2LtzhoMghPMRrCmMjcl+g7mNbhpEGkn
owk76leA+EltY2qfYlAWH/hrc6+FpW04tCicNHLEZwvB6yEmTUDZNWl/JA3a68O6hN2UNIMm3Qsz
MOjHZlf60+lX/LrqujTxdRKUy1m5kG9MdPVa7zpPHHZmlitO+TR+8Lu8c+cJbNQp1rFAXHjs03Gn
6+6qvHoH8v/4mvz866xA5Y4Ai5uvPSA0o7P4KkU7FqiJr9nciJO9JfhZo+hnWnb10Gl+GR5MuviL
nW6WQ/wfCYMqIL9lzkiDSPLA7GzOL5q60zjbbqNMzkmu1JhKwlm3uDqOVf8FmGeoQlVFLwzPuGfx
uINhvboQWuintzUTuOfArtjYsflDAQdWtXIzA67xu3RE3ryPgAP37B3rPCcShQvmyMbLdVwYr27D
h9Fdmsb25HbEZBBN7ufjV41VUDz4h+cKmK89mUf/1u97uG/7cp9ayiBppBohEQaz+J3br7/UZkFC
upkpH/wpB2ObZaGf/ZTqgT+A1+f9wKB4oR11KLwq1g/+XQ3Y3Xce7hmIZkViGVRCltNizVQHa5BM
zGevkk7Kr6sqAbsvylU06LxLQ0snpZ12zMS6Ls0mCy+QOXY0STYoMwfMrEiMMBJnI9rND8aKGFlm
WaPoIvasQCFCVkpl7uGIGmEgAwYk70EaT9hoes/qDe8Inp8gaaBUsa3+qtA0BZ2BTFUx4CzEqmH1
D942diPu8aSu29eai6v589eGI+XzaAN1pTVxO1VDtvW0+tV7XMsJbFtDIa86VZ0dDEc9ar/2tmRd
2SrMlKtsZo4QVqgxoodnmTfZ7NVPRvoh04YS98BaY0ps4wEomld1T3S2+69x9kqMdAbPJnyFzUO8
UFURXD9pgq9zkIyg7vRs3vzZPcg8IMVukArimXSSefTxKVQo77X10DvpPPnn5/SeT0aoM1uc8eZA
8V8fdistxXT4qGrrFdo6TX76oWJknh3nCqi16dFGyM9Oh9i0R1qvYwheet+guGN+P+obz5LAWk5a
bY/ceePlXK8HeZfjiYfCZ++yWQmFa4M0zcUTLna5clIiPTqw3L3DHcIeaqjfNsatwKRkJjZIht6+
7Y+B+Iy/A7qAkgYX2w0olb/n0iHtpWJge6w+GwBZd/1foT46MZEMaK3iv2DRyOCuPjNj4nzZMhyD
Y9VoAL3TsulhxVbTiunuD6Q2bOfi8Qqqzeb9j1O2+I/Qx0ZvHF8jPkaFq2ZPZR7R0MjW2beb2/MZ
ZDHqEJoRDFSwIFAaAVv/bfxafTK8YolRrOwuEC62ghBFtz1aYEYNdvwYNhWl2/59Q0qq/E3pHPqA
cZxCKvJZSXynL5xz5TdWyR+pkhz5jYCCaQV8PQgsi8M9OvaXpF2vVyIEpQPlWjpV7cOVvxzRNmKn
HIVj4l9uShUiwZ0FX03g8/+gxLLYuNv6QoPvIgRYAqTCzWXtnbWs/i1cmFfLE9ua0CLPBxz1xjzt
C6T4I2HBKyy2O5vvaFAmJfJPCLacRHy1VhBW5WKVudtOVF5X+VIQ5p+yCXArB/toOeyQq8Am8WKp
+ui5ekZHrnkpLw92ixXsiZgBIF9sB1TMitHOterzwbaY94uVCGBwg818TuwFW38yvwtIM0d/vFXp
W+buFvHNP7GM4YJJ3cn5zxd0ZCPTihaolGqmW0y0L2c0gd2wcB3Sgutm1xojqzMh1/n2diQTQ8m5
UFTRu3tY1TpW3+gmi8XmPLttPbMLOu3O6dmJAipUt3ps6yxxKv3BIxQFPQxUXiJh5gl+3Urbe4Cc
nPqVDXwo2kSDnNuZBHdDdb9rbyPKW5OScoIhJIN2pFBTN5aDU+tSzE8yJuwiOV/scM8LOfROSXj1
8C4XI4SDv1fIejvi5q+TK+QtzdjZ7I5ENMzvfXoKsC5nqwDsDjdnt9Wk/uXQzznShOzClFUWYbZY
ni750qBfliQ1J55/1bNsaHCqLqdAOgcQSD4kGcq689XJcXgg/DZInsGmveqeFdwUSjrkZUl5glz+
baM1OZgmFu27U0D4dKpbyJipr2DH+KUTH+APi/qeZxCO6ZAK2Nnto+UgOwfdsv1L4rQBKIvJ34ai
n5R9x+fY6vex1iV3YO6+oNZ/IcND05Ta2JAAfXFt4BlGFGMJFgGmbUJc2Wql6yoP3B3vRxCF73Mc
kILRuKmfShJK2H2z0vu1XnDfwfjyKgB92tjrJ5xbotgY8quz9aRvWz4bJCcu25yoJnMEOJOBBcCk
3TfnaqCvfHvvvO/LRowWN2pZrxtcQHGtO9d5UU4F7qIP6cBjw7TfZlokUsaRdHOWUkLCVvmZUFsv
4g/r8Lz7ZOKRPzin+bvcSuQ6FW+KlkJ6dUiP313QmUnlTfq5xTPDUEYx3libPkRa48Hx0ah4koK1
/4PsGBVY7CU1GNJmNEKePilQhoqIV7+fBRjP2ryMrCjWkuMhLI5jciP4qtnrXp5ts8picLWIBNQV
KTaxkewLlACaZ3/OyJRwPAUrDeWOS8nX7zO+H5k6NUbSORVV57wH4hoMbuT74GDOSL6ZSbf0UPSN
lo9SEu3ZeBIRUxxkYjzfrpKLSa7tiiNsAcz4wFXMLgENC3o3Rt/2qw4gzuxD7OYgZoUWnw+vfEKg
JTQXOsJmay1I5HUE9ViPw4QyY5lz87W5+K7yROY+aKDRyBnsxP95yNOHZG5iDbXnvD5wxT6Dn4/b
HINhK9XSC2Qi+zkU0+HIPGve8kjbJDGaVE0KeZHfZ22X2x4e8i2l/wDlvhujw1qI4UNTogrNR89c
z+gU4ljcsiPQO0+RSSLf/XUx0Bg3O0ZKxnLvbKTe4HcBNldUFDG97t1GBA8ZPBDQFqRwAMZak+Ge
9S+oQXp/wlcT1Mhz+GiopB8yOjhe9aO7hHPAmuPye13u93Kp0NAsS2x0GVOMLNUQIF9MohsNZQT1
Xxl81eQCwsifU6vJZY2XXN/L6VZ4IOGfS4HFdhQBiNV/8PsDXg9ApjMu/wy3B7hO/400gsV3i0dn
npmyAViMWND4rI12g9G+Nw7CS9x26bR58PHgoujT1g2QiWKS4G1jZF3/9rDBVxROyC8qzF9VjBG4
KUmTLQdr9Yil34GxkQnxVtGwzMzu9FNFPBYcWXdc5mHAUzTE5n09uQwL7+6oujO6iis4pFncsz+A
KrVDVtQxiR5FykoKk2lxxAUpjx8KG9wuHq7nZEbjXbNh49Vs3HWqsO9pj+hVvJrfTQ53fBHtloiF
93x4/nUOmEua3xi1VjKxvZWTp8MNfh5QII25vsOjury0QenOp9eLJyg5yy7EW/rbR1Hdd5EwbvTs
auL67syjZEH7wrjnqOM00j48YM0gryw4bZnUYJVqE7iV68zWvC0EICukZLRt7/wDAm6KDQZYVALt
gyf0RLInlTmcIqLGt8UroJbyNQxa6tIVw/3rjbT2ApvA2cZR+K4FIMcKfIVyp4BJkgNu3unFp+yJ
TLROUE4XK8uk2VpqqFK3JYGcJUXGuYVGU139yE1en3cVXyUKIJilof6BtratKvxMlh9q7f5Ff2Ue
bcubNq4TE/cCxT7UHmAezN2FDpsopjephcklnO7tlxzOSQpu4jPVXlA7NxEevbc2a3KGH/8au3AY
oVaMVQetwntAPW0nBBDMlalBxuDC2ERliJ1/qm2ABK1NKVt0K1G/9CbUwxHQI/ml4keihH97yFSR
FcctMpwut6PqkIfSir9t2ZhwBK1qqwuoNHhGG7b+1rUBlNS/ZyamlgjoL1EVX25NKwKVKrRRCyZF
xLzUIeSwOOS8LjtUMIQhV5Ad/oywan5iAnbiCRYhKsZc7yIJb3eejoz6eYoxomeY25WDlI2o9cBJ
7lwJ6/UOgY9Og7QSkLLTOCeM0qHlUxnZDi/mtfHEmlGPv/tRRPNu1ZyCtOuxjTRwGFUo1ad4M3eR
w7LvHD/ptmNF7++++lSgNtdx3Iu2nujIEA+rjPLGZlPP/TsiKJdBR6EWwbuLEoBPR/PD3moQnLG4
qfY6Wpz1ZYAaLmytflTJrJ4AvSNzETyRxuhLVXfLeVCVx37MmoY8bSJ9MixfkHOi+suFle4JJiIg
eA/Bs3+UW6o8Fv7MutALJvJcRYk8bZRx3eEBqfKaZimkNkp8OGoXYnMLRezbOCXW2h5bBfUZ16Es
Mrno65+Gx2EQtIrHhDY5C9zDOeNEOgkQyrPvUkJC0xeCZErZNvwUapEufip0HqZz03/CReKpPIm/
E8NCwjG2Ui808LIVIPybPfWMWUWk55BnGu6s3prnax+/NQVugEwMj7g6rZXzbcarab0optvUSRjw
wwQzMOkyMlICSn3/yp0+kHvQH52Qg9vRzvGVNwCTLFQHReGrfVRPhyRwvRhOeCvaDnr7YRWc+vaB
efafgxPHZ8lfJEDGWIr+95fMkfOK13NQjgA8bKr26zQhhHLn25pWfEkD1RnAOkTGp7FxjlEV7k6P
5wiCK75DqEeaRcF4AZEkPYIDK//fpd/eJP5pMTwTa+qcZZJRhX6EtGTTgHxSY36ioODMGfkl5X2+
fFlF7MTwHwyhizcfvW6s9Q6qAohfPn509Q6s8Ibgq1Ft+nrizW2i0Gyrdr/vPZjOHS6zHI0kZ4vN
4qDurM4Jbf2V+jkVcOBs0/ExaHnXK5aUs50V30Z0lMwlYWFbFL/zIxKUUAYwt+VL/8IEZXgkdWw+
jYdsFa4lWzgkrisKVPr700CHNh18VS5MOtGXRjKXAN3JXyiVDxjInF8YOxe+w8eAyCc9NWLQ3foh
f25KNnyeS6Z6zMLxvOTTSU07cnIJdmz9WKDXcpA4X8FjmgBehkoglFIwSV2d84s4Y5eu4tu9IRsI
Y5O8mUv+l0zagtaORyD2qdQ1NDlvkoAmrNhYTzhsruMpmofJ2Cgb5kVBrtJ4+DvePU7kJoqhFBv7
YKRoAYnYnK++7Pv+YYLzD/2QGWOxb5g/7Yd5lbF+QeozlFLkD0jyCjdSF3bK4zZ5cAP8hkuAMt/5
5UVFC6xVZlXzX3ElMHnbLN5q1/i8iwnrGS7N3PIcBcDaPKSez+6GrPBKaaRg1PL9hPWaVior4fuX
opBT0wzcJumUSMbAOPE2MJzUuIayxSZEO7Ti4Sm0rdtkql3q9VM1cdHCDe2Fl9lOx9I8dNUUb47K
H+VIGyhw/feqQudGy0pspBR7Mm8LnsoP1No21o+Jh3/j0XGPlc2AOB0pclKGIRdZl8eanDlLzwtT
c41wKtK37YfV9fwLkGLeuuAd57QkqD9HtoaEYR0r43g4Myl4iDUzPNVyYnkLyGjJGoDTHwZe5rm/
ojNS8zqunXQwSRTs08m6KqWdqggUgPPnsF9tSqd6/fyh7twqoRJhDPIfsekJD3R72XGxNm/j7qsd
iqUXfim1nkyPtkWRl+OaIqzbbvYxp0px1HXg9tfNFNp38GaZi3Pb+8taDVHEekfhuqe4JG2OMxpa
KuGLLBV3uQTEMmQFRh9Kc+YlZWXrAwA526nRlKs4KYYcFVx67/cwbC0GuKah6UU0wxjoBgsKf3zp
cyCI6oqYTBZGId+E5t7URcEDfbF/Y5CAXspnTLB1tyOELZv+idKj89ThEi3Kl9U6ScweT1suAVsE
WklEESo50WgyRjJRnZU0wM1y0IsoU52Gbmgd/4dHF7yRkKY0jBkeoq3LGt+k+SiMpgGg9VS2gkbr
zoe4KXGeP89ygtQyggIbrnhtirJ++leBzMHComgz2z+iqRM1NmJYQgUFlfLpaW9M5winpNH8EofN
Xyn0IEfDybq0eF6z5LF09SfuRb6g3SAYi4fbUhfMB2SP35KLfSfwSDvCxZt2wmsqbNQyqjkWWvKj
bXA1CTAfFp7cAZawV0MbqPG53aCXNbL36eqr4j/pK4vAlDlMvrwT1koNOyn6WoSGs5oqglVjnrhc
MIHB9TDQs4KnZoNCtHcbYkBQJ+YGJTBfYsUcmWJFFQZJEi+oU09yjGO8ioDuS5qG+EbxUVNzY/GL
Lv25wbqe7KxgXjtW+p7ZNeqoeeldZ0sjzFwc9TPZJipDUygaTdsM4hjU7ORcFy4ya/K2Zcz8sDEN
5vPWxwyFQ7WdC2ybzbWLoPlcmGeLLsd4g197Dx6C361R7g36nTv0BCw3IYEbfBAzJS4riadldhYO
d6dDN0tqf13Azk5k8NVsOpO7Dwhn2xKC9JhL1M3051uY+WaKJWIxetRXlcAgVN2S00aXJoRGS+ru
mSzwtGL8fBPSV33LjsiqxjnymPMigwOnIliS8O77M+u/vTjZj7qh9fVLCOW1zyhNEC0x/sME4/vG
Lt9Jq3KFUUJSndplENiY5Hvssv9GT3O2XDoikr59bK+TtHVz7Sk+F7fk/TqKLYhxmRreaK0iGgeJ
5eyaXLcVEkX3BFR7wlh9qIJytN/h8HI99y+QwjiGw7/wSpss2SaK04CA4GjL0I/BiBO8IjCqU2Rh
boHZiaOby5nSAJJ8bAFVgr0FzYRg5ZclUyMFiw7quO4l6FmAPgTApMve+5JbQhIVte9tv2g7FxWH
X3JTuI8rwcdP8CuJqSwdfFYq3/dOF72isaGkFW1nLESlFQ6fivUG0LpaTsJDisd20O41+34nH9a4
7Wpo4Ns/Ig8wHIM6NCSWRtQm9Kq4Lgxes5aDNtdBqGnE0tTn30m+hfEDUYxCTC3OEdkUV4PGMqr8
2GQmHqZ/QPzAyfHpo+WYj8/NYp/hoyq5D+9zYQ+7yJLjlEafXEMqQxYJ3NqdFYwUgOB6SIfnFaG7
2IA24SA/LV9TFgsHvuA1FjvafgbCBrT2+gFpvGFjtEznIOo6AyIJ076dSzMHNyECbc8jfntmDKDe
vRUbKALoB8M2EMxlWKn+32wp+gqNQqfciRSKNxi92UqLkGxoT3i/BTMl8Oxkx6ORo+XN+8L8+36h
238XJsulo0U1MfJc9a81yFumpnck1ON0LtLzROzCNHc4xWqupLIYnmXlZD6YooVVlIHB/wn/f/TE
w2Y3NORVM55d1yVgz8gEpyttGJ/+hgfJWx+/Vaz18eWqFlBtc7bqI/o8dYNCKhRA4yp6C+gmMQAp
E7enoGEADbo7kErt33Kt9cPj9C6Ad5s8P1KAtoRo/h6etQmTdJwLh4BtSS4oUH+5DAWV0MRWaHil
XHezKy2e+WgYKTUUCaHmdH7gYOwO4mkUXiN9ZRlufJqcp3mNUZS6hisur0493r924zh9dm4yNzKb
ipjZTDKlsCKNezeFD0wOXMkFbXqIN/3KYXlGBBTSgZUSluG+sskvAjooFUxFCxFow6j5yqKSThip
G31w3rPSfkZlhMCQgUNB933PX3sVh4vFQzRQJD+GfG1cQMKDF/VP40IYtihM0JslCX0uqonTUgjc
OQAx6Rs0qtOg/vSfX48K2GCM1qwIW8guWP824nDoNNasWHIUDTGUJhgriQdzYNbAL+HSzTxEJzSy
j2CO+0kkPcORaHZRASpvschKemN7vkZHNKED0okizy9LsNOaam3GaayqjX0Ij4wwR50Y+cGfdbzC
egqwanNDytiV/fMwhd6xZ46JQy5vZdiHRklFirX3eigrJ1pDHQOlbegbxgoG1xgSlGl3nMsw2NmW
Hbuhw8qaT4n2M3MhB6DgNxbDSpVMHeMwa6mU96WvuQGNZMoz0oG0QHSpfBSQf6+h40xm+SpAYuCW
kEmFF6P6GvoH0zV4+Ykx++QggCRt7AsFrYOffZew/XVGgcLq9sLgL6y30nwZfc3Gi7SH4fQnLXh0
/+Inuf4mMcw1FMSKMyTKrlfQfHpDXPhc+hEveHWDiDsD/G2L47kvp6RKEWA606l8EeL2QsErBnpm
kkSClXntxoQ9NkIZQLNH24SYqm1UjeCLAQ5TA+/aq1euVWS8JOitR39FYMeCITNUX09UUMnSdCzU
Jp8xr3p+R8C9Wy4pz7BuTvoEDheu3uQalDb4SEiUXBiR5QF3EBQJNvBlcEor3I0x6c1wLjyF+klW
I0SzQjJWrmBsSM07IO4aETWB9a8v2V2Nb+XQ0LqP864Gf+qU7xx1NRnsLCY4tkNt7fIBMtq/pr+U
1ysTQO5LMkyDJWyjRAfd3jzpgujvyn2xLJ9dqNj9mOa5xG7ryDGmGZ2WARhB/NlIpGdNJwZ8l7MI
ZOJBf9RMQb4PbOz71jc1ZLxCaOlc6PEqBZVTJxek2zqTQQi/Cuyhfa7XHW0rDot20QUII5tIjCst
waD9RIUOA0WMGRo+Kqoq8aYPaDbPpU/3vSX1EdfglYeHbiEJggZrCjF2vpO6s8m0Hm02Mgrgv+da
PCyXJtaAQfUdRZgihvNtBvWW0YFT8bL6n8ii/eHp9vAX/ltcEcS10lt48XinJrsUXb3DUE/UDI6Z
UgNj8ZMLV4BLIQ6keKcrmC0EQwWbXqnFdQk/Uf8Ej9Kp74vdQBKUhNzXE5duOqpdoZMS0kT1u4Vc
S0u+LHoyW4MZIlDIgwtfPPlijQ6nbI0glc1VSf6nOYC50xK5g3Wzw1a/9mjLfm3ZxP9xGRDIh+x+
1oKnZY8fG+n2CnzT4No+zqu3N/pr0/60Yu1Ws7CXs/Q7lL2NaMBA7IbMdN7DtsWk2WboZAEGSPAz
68tWOIlQi8ZUhp8pAS0I5YvDa4OSokwMWm20Or2lsB1e74u+O0BZtgXozCimlyhFxCHWWhySWjb4
Q0ATQprnYNfb/KA/rgc03dId/GUz6t0lTWbgOde7POHlZK+i+nOguBjt3E7hNiYiK09EBWaKMIDU
eVYRRFZF6w7Cqhiv919LgBo2NC1d2aM469uKoCSUxc/zcjGF2gwuH2hKZXrJXVDF7KRn0HAYn6cK
4E8x0aKH8zSQm1NJ205OWxyY+1s1fdClKa0rxz+zNWKccIqa0AXRDtrEKiKE5MyOqhcyTw2/1VEU
gs9cXEjmPv7CnV2UqC0E5jZa02bBuso0aE48STCu2oigz2+cTg/0rUbQ8OhKD2lBDEb58c01CFRu
D/6+fjL5RCFEJyzJunnAv08XOG3qJFM2SUJ/rgfXV++50Jb5igb6TH+wj15Zn5AaQRrgM0Dty78p
jHTvHMa0+gvtpMb/k60Rex3cv2IKv4uwxt76+L3l53iapOl0qWAzsZcl/HZaTQW24qDMvKJnilmU
CDvkUJ4LWnqe7v9Nh/Qtwh5udGrPoRyTIQUWWKEESlCAtgpLu/cWkIg1h5Zty1hKDrAc8Bf+I/AU
ZqtRf4cXYWrf8QISsAQgaCbD0+KNrmn7RRijwXUVm2spOZcUAyZAiNGQZoCIdJzLi4Yx1kMAX9+j
9yW0ZhKpxVONOm93Maoint34sqNgxoxZbMWwvchLIdmyEfx4JiZ8zbcY9MzbarSw3fYzHyNbzFJB
Yu/EEV9STfVvE+ploIZRiIMCtF0T6l77c4GDJSSchj73ARvffKNDFf4dLe7twBTOskdJdgJCUBfJ
og7FmrnfvQBU6vs7iujoQ+lF/TSJWmUCqq+6NsRDaEbuMNl6zWn7C1iY7aYQJX1gUtY+pYzmzmzf
DHQbhJ16QjSkNDuWMvyFfOiCU4ygYe+MnuixKTomL5BtmZCO03fdKcodNvrU6HdRaPl2pPCavfWF
VVO4vux4M4q+p0NzhVzjEGsSUm4zi946FIKri6layPq5MjN0XA3NWQRThdKu9aubkqm1DOp5jL8e
WMZgzmNulfbBq2O0hgVCD6d4LvaqOjo+GfWWpm1pylwniKV0sHHEJzvkZrLMZYw4Gs3SevgXgpRM
q01FDE9ZeOap09vMW+g38XjL+cYK1L/a1rDhbCqWEnnPu2m2rkwskNjjJ2sVN8WN8JRVD6RYtp5D
BxXMnmFavcEE3g90X98gtu9cYofUNzS2Xh/gqKHvlYQvZ7E1F9ho++oWSOJQmNw2clZ2dpWYpXa5
thlJhT31WwxfnIkvJZvm/oakIsXV+ZjHullazMWCr0nLTudLDcArmVfoxSBoFBmHMHk/24B6Fhbt
1rnhMVtZrhsUWwI0ZKFF5UZEECs79k3zSc4W6ckY8CnikaNa1tMAPQ+JpsLOfxYx0lM+XtYa05Zw
8+WSc+cb+EF9HhuYAsPQtf6h0ZnjarTsExXBVbl39m+cBblipC9ATgs0ztzUj4RiEorJaQGGPLyC
R1UaWclPpAIbk6TxKmF8/fR+dlZKsFBrzyjlt9WofBLYnkob4Oh0U3Ev1F+myaDbyyYPgZXvP5Zl
3G4YF+wcQ8FLTlLMG8V9GeuMOco7lmYvPWqgyjv6mZJsLn7anWDFl64SFcgv+IX1KcA9g9MFLgiD
9BkpNPzBc/0gKe315WnVDrTri5nxnkUXDtqOuCtw4BEFZPwiCQ9pwfnVWOYIZUBF1rOgyrMedljY
NTcPiqmmE1BV8U2yljQ9nEwuHa/+5CUV/83y+XtBXztQVzJX85TrlNfBpqYAvVf5RlrUDIaFO7dS
jRapLH90aoR3k0v8HobKWli6tNqIcHLdqz6cxEzOWJG8we84bl/B70kIqu7EsrFLOU+eNfpgyHLd
Phq477z0RqPfjB0rpxZnaky2YL0YVMTW/zQV1vXE03XiSQzg4LVsXx9NCRZeISPqfYn1FWf+EGUu
Yar5EOlqFj2dQClnUq4N1yf50M0TGzDhWXxkwu0N5pFpMjJRly0SDZCtA13VeCHiMOqKtqWa7wy4
n6ubBOXv2n2iotQ9f0416qWtP4F7Njcejo15KMwVdhXyOvOaf5pjqir2HSxDwdxuanFA5hTmcqIr
HZoPITYwlajmHs5qI1sbnwPpjSNdfrcXYOzqAq+9gUGCo+S0hSjwQO6f8UvNT7/0eZCGceV3BLrt
qfWUDFT33tv0ITVi4Z8ShCC5z1wZAxf1QsjlJK38Jbnwaz12zxo6IWDf8mKBrFm4uyEFNGopK23G
Aq3AtH2xnoQdLZdol52Ds+x67V93UpvyQWlrdEF3ksEedS4yuq7sMZgyRw6LAwsA4WW2sp8joxSA
vb2Y4jctaP2QJ1au4g8BWDWf5WGfKtvbz8OGLlEEfd4vD2AabofpWLjAFP0qJefCOCeGCb4LyikT
3AJaHHyGnEDbnPlHijOYNeFAcdnVKtQuMMPCOPfMNNcY3HijPW4sVIaFW3FH99pWyL1bRsswdBu1
aalosXtje77XV+18WqFc1QnpLByyZD9Rv+ujyQVWevd2Td4s/psx8TJFzg4pTzfuX2ecGUqeyqk5
sZzPrUpjrFf34aSQ7nj1NrcAQq/5Fb1qcaIEm8gH+vQC6J9ix73ZL193A1t/ZAXQ0FMcIrLNuquq
jPcpszwwAM8UWNRCd8Q9xmxagndHtW9+AJsQDt4LCYZdA3vKWSXc/nWmVjR7MhTEvZhbbye1H+ZV
0cOzBQvJo/xDSZ+vSq2F3rvu4ahE/E3Y4SOE0Ujf9tz6vJCixcYzWqw4L6DOeLr8E5/2M0LX7ga7
+Xe7SQLBEy/G104JDn7gjTDnvRjI81r1lTwaLeMCIshd/cpjG8avbrS26QS7NEFTrjC8PXeU+kDK
SIp5TkrHr9KtntC+IPO+9OGqauZTnctIkhjpjUJTSRSWPG4ybMpheVRoyg4cyYtmL1LRDHciiRMf
dqYYrJTaOtz0aiP6NSLn5ABPf1TEnPWyolTesrvx+CQqBKoOyfiXeUxnYxsJVzGyF9tdPJ/8EpQx
97EkjUi5GU9z96BvkAWIpyTzGdocujnRlgJozt2IVO9W2Cz8QBDpbMlOvsseKURJpqdD9vtFFSzO
z742a22qeYppeM6qjSmwDoOJyX+u6DNjYJCu0kw9n0U+cmxhZRlNb206Dn8b6pP33t6Eh5oTGc1v
+kSn1yuQ9akGcyG6jPzYC8wFmwMgTea4cy0B7UUBSvHW5zcNxgGmYi0kxgxG2GVZPdxq0asXSKo8
kA+BP2YDVmraN5O5uV5b/7wVv17h0V37m4J/4LaBLHmapfSeDIBq4Ev00LEbEyYC9buXWuCm1+Ko
FW0hsr7CZnk8eC1Dw/DZ4s+aoqDRfr5z5dPsX4Jsto6Ereh+uHTs+yMS/rcEvBT4IsKXu5irSDzh
vhTKN7dnyukX8OV2yEtywkHOHOfc/AdW/Xk6mhuCVeCYMFgKfoEP+UlzlvdSefWP8GkK018Ro+ah
9iKEimZ2L9YULhJVEa6BdNSdCjxPo4JBbjFDfRiX21EqY1ueDMR9gzZSNdusR9c05CfRIzQOT/OR
D2PyOme3CxtQvMXSsR3jSif7Ryu1kUMHn55wCvv2ibOSvuhNrvV287LKxiUZiDlNSg6brAoIVlTp
oOiJI0Ty1RadfZXTpVG1QtmHMQwqTG8Z2yYxV1muTLpjVQTpXX1KSqUlJx/zO9mw5sphfWBiGELL
wTLb0sNcCkHoBPLl79Z2Du8ZMK7nta5u6IuB5gppRTSyLyxkbMq2a/96B7I0roHyV7OzgS8jD2rz
v0PpwH2FPGqv9tO5HNwjUBJlQcUasgxKFbAkkJNPu3OGEAcF3oo9BhSSAl6cPL09YjONQEdpmm+4
ly1Yd+sp4Ukr8EraXZVthbgFhvRGhUw8Cb9cIAvO7T8CDvfyciKsg73ZXR4ulbg+cOyrjV4RE985
0zXu8kKBsiJiI4QCfXwR0YfM+MWpq27cXUIllRYzhY/LtbRY1RSDMec7GunJXk0yM1o+t8eZWoJj
cvrAppSXKFETzEt3vtqtrlfC09lQBn6vy7BrsxpqDtgTDOenR5E8bhxmmjAD0gbd7oM/honWaxkR
7+hr80nfWm1S9493TsRvuDBWu3xKOPzR9VmhLBLgdyOme3OtY66PI/7NWPb/kW6xchbyaFnekKl4
ctwXZRvJtJNl16M8UgC8uwiQt39vbncm8bx7XX6o4w/rHdxZGhjktZRydh/vFw+aC0Tdt7JwHKh2
SRSAgqaeMJzRvUh7OuuZZDnbyxSgZ5z/JyrIs1QJHv/DERu1L6jwKR5xq+Rdl7FdJib6sV2/r4Dw
zhWd8jTICD/9Ix8yjDniJ1UQFH0WnKUnU5eCMQMZuXqdKZoRSBoKkiASiAdm6/AZxgg/GRk0tNUY
67mRcqKnwv8vtKEEig2IkZAX26OCMI2a0TkUxdMqOsbMloztQ7t4CDaePXz7SolOnC4M84pKeSGj
QgvooVBYil00qpIjxgLaYk6l1e+Knwqg91wEqWfd3oqnb6aBB9g7Sp9RPdDAQkm5PN8cCsSJ4u/B
0YTQOCC/iT649dIGJnldR9fb4nYZEdNuF8iM9LOeFjOxmKCK768+gxv493x8b3NE7aPzZeOVR/6J
d63q56SHoFSyCWkhjAx7pARBUGf1PHO/nIV5oYFFTalv9lI+VZ1VytOpJ+iX/HAJP0Dmwjoi7EX4
dEvCfz1/zH+lyrb2Abli7kgS0186+IXuBAZtFZv8KvvMN69mRFKeyaZ44x3rT9hJYsAHTjdnBSZH
3vgCzPzo/V7p48OBJ7hem3tAvuknV8WBlgkTSTM7bjbcJpwmhj6oCE9Nd8TKSbDgakAXBwEyCObM
qtyUbSfG/WiTLrZHeiKz4PXb7Zl1g9umoK+yPJFfRIVW8QoLNvmSQTp5vDpoT8Mdkw1RxSXoO/pA
h0HOBhUwrqx26VkZLm0YwlMjp7BPiv+c3jOkoSjhJiPql/x8fTCd9WSlNcc/XfKKuir9u+pO8woj
nqJmOBYw05u1aGH1sDhXo1Wny85+gFX4onRPE1RpFpsHNYtWYfdLIdAtKbfz22YgZhB5tA3sRQTX
nWfTEJYLE5YZAOBF5Tw8wTeLb/7sgmyHX2EBOM6ZtDxUXPJSjQ96omiiZ/CIYv+SAUueYHYDEnIO
48TbTQzEndntWa6dn4fJcbbrEKLx0ghUdildoyclxhj3HKgOEhJskHdFlo98rIPz6iNdHSZE1Fde
ht144uDBe1aZWBJP0/f7JXjwnngGJE8NETN29lYlXIKc/4Yizn8bYcmj7taGqeWIPFvSlPgWrjrZ
8lzpnnRVajbRNwbqq1NdsD8XHvw1RiSnsflrG2vE0BxOFNiPQvR1u7a4ttav6Cggo2ip9DJvol+g
Qmi5cZx6dhtsmF/VwvJuJWJVyHUtHM7CD/8R7np9+Ty6fZSgBBCi8EIYdh07OI47MAXjnlbk1oGP
7TwuSEO5trC9BiUSzebeKn4wi2MTGGXZAk0ITd/tBHOo5arvkx8Y6bHvvaE3pS0zyDuQK0bi52U4
066vHmYuCMWc9zb4xi2Hv4YxzvrlxgMehKpkD67LPr9emrszrQ2IZlrhkamGAkOF13ipTTrPx2S+
9APK80fIidJEG56SEWuoNEYq9r0uq8YPTaCRrJONXUz/9WGYxsWCa5Blh5hXWtSaMJJ6rir2cSsX
YN7jtMIfmFgE+vffZ2UG11y4KvccufCiLZxsSpPLMOlD5syxEXTR+Dk6gSANitLIqZbt7qCC+HUp
SRuLsRuh6SK1D02RPQm/HgwYWDzqpS3LAwTYB54rRoBbNi8WubW1/T4kgialEn8lXItq1VCyapVa
a9+HBzuzFKEHcgxMV3slHWfy4gsqHrJH3fNnhIZbQfSLrVPtw7+1WZcBFKGi+vQN6rgXVil/lO+K
EFYUAGZUnqk/ga6xwcTM4gQieA/b/yCpEmPXbWs2RpjSvvLvltO0Rfyw8be4Wft9wJ85hZ09fDtY
2Ezcqec6jCA20t2q1hpw8rRen6ndc+gAYCQf0pbm3b+hrGI2u8HiuFuvecRDylCJrc6piMnVursK
0uFIUe9CIaFO0udYyPUeel0u7yz1Txlt/JeBgylk0TQHnKn17XH5nDsv/2L6pqb9gC2qTjcHaknf
0GIaH9bJImuoufUB3SbFYlG9Wqo2u20FDt4Xr07kn4FmlmqPcStNEp/wImzRsQ0jLEi8ZvFNYLvb
DNq5B1j9IETasJRl76CfPk2vh5pF+J5HCe1P6+Tz23kozr0HCfwQ+F73y8gl3ZLTGlPbYpcEXvc7
0KWv19O1iCbcEFir4KBzia4M7biHcQ5V2I01MqbV5iV32FrO6d1nuxwjfJem3fJ3R5RZAstBtRt7
3h6XfcDoGQNFy+AB3J/iL/uOpEhyfmUaFdi7h5pBnjrwzWR7QHAFGYXecXyzAneM8ewa/IlUcnCF
tRZUTqnZjzVlNy/CeBiVfqdgTzNiER5VCO8oyYQyH2OsI6caMl60kvpc110yGbVJWieEqr37LkCL
MfADlILNySWDqivxQXyn2PL1r2td4nTX2q8cUWb/ARVJ9TOvH0CVbUBywuXjHV81uOJSnNunIbI5
8hC+mah5OVww2EauVh9lNHs4VKq6ydfLtBCrGUIqyONcw4ojFZRRM6q9B5TANhMTa28Bo1Vhb+S4
YOJuo9+s0Rk0pOHlThRWL8Gm3GplDQ3bI1WPlLCYkPqzC/GbtYqXwe9HqKqRJVNYg9nKTgM36S8Q
WCxlP8M8+K2OskKnVLbd661eWL/zk/zA0sfmF4n2xSD7zSG0+g1ub8e4CHXUUDLfyf86Us4VtRP7
V097mH1igyMTsJRP/M1j4VAFQQKrDby2+AYX0sIg+fPtHaFTvChuzPo8pQqnI3s4Jw4VV+Yrjks6
JAj5K7Ne50weQGUV8xEzukKHx8KQsNQ6wPcO5Z8+K8MQmaTIkwb9zqO1wpF/6+EfluXc6d+5CUy8
fUqctYuQe1dDak4dAKxPkQTfOO6dIgps5oLujvEOzHY+ivkXoND5REQ6yKc/NKikFBzAgiquC1Rw
HI3s7p16k4v1wov5ncNSdEYqEOmpPfXznGQF+5xviTdp4WnAqYl1pMrsOX06+34xIFSAGY7W7AaB
lw0sLVbzK2d6tnzsyTLsMm3fnfaQQ3+IUkxjZvJYa2oa2WYfXihKOXmAS8AnOFO3X0n7i+QL1IYO
NjQMo9iG9Qr6knm9v10mqTZnyStPV/AWlCKeWp+aYYcE3j2lQ7TZTrvioGkKvb1fL0dowC2C6YHS
m7M8OYBg2x1ggJyMvUoOwgs4QpUBUur3I/Fv0OQvNHhaEODfl88/+YTHZ/Nvg2JD1hywfFZKU6/9
vJ99K6MhhPeV33L8DMlH8b8Vp0y5nnJFxhHHxM7HujYEMmoZ+hKtOtKVn0V28r+FDqs2XiThl82g
xrlyhbuEQThaoNeQFK+QQy/qQPT83XSX4UevocCglnvzhfSSzkjKFWxVTApncNruZgIuC1sXsQ4a
9CQ0mEeiRxfrgt1tnRTYKIKkDHIu7cE66lLW2uV7Nc8ynx4l6LpcSkeEsPz0pnK7CKBKklI+6e4w
8AXY/kFqEibDyos9bN0FwQywAV4toaczqnczCz0zspCoa3xHvdhyUUuSNsOyxIQ0PeLeYShUTK3W
zdMBYKdz4uc6KfrEvzFN5ZMNDv3PU9T2Q9+sUUbY8GkpBLK3T2c9km8w+TbrTTdew9I3hhZ0L1Ta
/nHG8U56LZcJpv7JmXTyCL42aJ5b8j/YHtUQ0K9lskZrTK0lPSBVbifhM27f3ryVy32kssaKEAaI
sVVD4JlOEBF9TEg3CGsg5DGmQNO25au8s0EE6a76b27lQ08SjYrPbUUgyBpIxRkRttPuIZbOQrmW
KjQ4mdeq9/9FUl9ubLBxUunyg+H1pHCrUtDWzK7ZXfOOoki/ezzvmTIbGEF5XDhMPiuEsaHIP9f5
PgVYGX9SX0wDshNNcurY7d5H76HyGNMLZENTsBvmTbG2Jna5+uSGRj1j63inuvuZKV8gA2DQfu3c
6ysuH2isi9AWwrgUoQsD2TUVM7O2Ad20o/7L1VrjIWSm16ndWq9Tp8PAcGUVGQZTaxinXfgD0QLr
jRBeot28bXV387Tj5x9Ox1lr8ZTHCnNQbw5sQ1frpzrmFz3mYEoTev8vxHbzK2Q60HIaRDG6+rqk
iDUgvb7jUj9U538mFcgqVC/e1INApTKGFt43oqTbDpBAiKC05Yxevw2sbBjY7jS3IEnGSrHccLN5
A8hnTGxugz3MPcfcg95sTXONBxaXgAT4cOYM3uC4kuSKOBtjeUcwYz6mYk3T8ms0L2rp+XPbSLaX
JR4aFmIGxse7IK5hQJTrMasCQ81qCa2wB/AcLvvtHQ56IFgJ1YucaI1D2cQcmrDT6D8XlfGc5luT
40BO5eFQ/PzyWog8dTMPP3ZLagAhjC/qfqf54Ugcj71uaIWriEKhOdG8a+ByagKByH/xAjSptTd5
/o/lSXsCr3zO8PcYznpwOz5vPcxgCsXQG5MNcgoX3BtPD0WYcPRowMul7jE9KyZisrMuqE60twhr
0mIFO2QpFbUao59nwiCegTeeSCy5+SkD3umi6ECdUIrJKNMUzaiPK5FHXZpTAGTrG5dYzpKP9Vzw
E8PtSogl125dbanF3MIc/iMbaEY5wSvt8YLVYb3e34YsNu8yzgPlveXMHU/kIAquLHO2aF1nF5Ky
7dd6qrEqnH8WWvtaRNgr9AZcTwkwIS29QvCv//MpPsPbucRtd93tfvy1De95XAdUolQuZSKKNQGH
+m3U7jGlGMMSgC3PiXXW4hOd99scTHPY44zMxxf/dYOozp0UGE7LdOV+0+chOJUw0e1zxCdFLgaS
ncNWl9HfscC/Juu7mYLLRD4JPjO559i+vYQvTZQ1W3TVDB9x89BRVuAF9HN4sLuRGRwPzxQlrcxQ
bOJk4DO48xGC8DHWfekt8MQcgzPGnQJb93deVeYGx9ngS5yh4CQHUwYg98WAAqEks1/5iYr7ISKI
dGU0HSBii3N8k9YWMxQQDTSSsrrUtN+sGt/up0dA5ORHiMEq3Hsw93x1qkuk0bSEHB441vN/eXDS
8/vTudx7qb4dx64IB9COzKqqG8bgocxsy/JNfbENTw2wekMEPayFlhMBYIJbveY9AvRks36wXBpB
bcW1Z0OOQPIAScWr9dSy6wGWBdIdMpNsDb5NOsORNO906mjb8TCT2VjmPlYInKsjBjq8Y87+mUSA
ZscngIVK4idPj+VRvzVK8Mb6S6cjkOIemNhibfsOuN9qYiHVA0/SV91mMulk+eijvxwVdrhuw8SR
6slxbyneNnBdhgm+yDOCUApDP0NQWa67RmQbdixC51F7k32Vit1Z+Kl1SKVc8CTTcV+++Azjubyk
LZk2Ab7kTCQ/zlsIlGk82+TwLFdIyPO1hdlvW/WmoBVs40j0koFhFol1SaZ7R6iW+VhdOTcrXcY/
rozFd9EXp0HrAhfEdQtlqOXLhRXe2RgYnb5XvyaMe7JMn/EBNeS3tOauWnxL0HLEgROS0DP/AFLg
vQhsKZCRpFkQdxqprrUhbxVIRrPbqFnJcP/MxYllb2MuAcMta2PnhdgEF8ZzNyJ0FDuCZrB/4LjH
+PU1IMRz+mzWioyHLMU+T0UnQaQJnsxttngxvVYibr9lcgTXlujgZeuj+So6ZR5sgvMq+N1sxuiL
J4HOW23dBmL2j7C7yi7ZuYVhGFPl0hTrL87VpYAG7vdrogSE3WTiStnyZ55n6ak/OOs+mz64U7fm
VYFl6nDH+y+kxxQ5wgfpp9Yi+VCX7i0+apxF/dTD4PshgSnVKSogEau3GnXG6a9WqcDAmXOzB3YQ
Koz5LN0ybd6tyyW3xJniqvO/h2stqajtTyERd54/B5N7Ll0kHcnNR/v37DLvCSJEuLsP3LiQ6n5t
VCBw17nf3ivSAZI+ZK+9Os4GlBn8AXmXK7TtQEGmaZZgSIMO2tHIXC7vGs+VBhYH7olPTvNpQHHU
t1SdM1/gaQJEyxP4d1JO6oAHtAtZSuOytPV5ZmIRrcr7K8cp1WOog0sS+Ozxqc01pb+2G6/NlyhS
HW+STi4qDUpXLxR9KpdAU4x/rTeSVuA8lBbFBDh5/VS2uhrTaGnV2Ytjg7TzetpgcXdUEVJoauxh
94EC+MnYBvIZMi4DPwNhXBVgkEF1sLKfp40zuytDyhtWrOmqr9MBTOV+biVGsagxdmoVW7jfWY4M
7VuZLXivwn3xsaX1bBpG55TpTNgy7cP+g8AYV1/utOTSUkS2N+hcdlo8DGoQolk6QYwFV3PE5jlq
AX6WchymefCMckw5v1qAmED6lTbbqtIVQVoxjRphnxgfy4pYfFkjDfXX068X/bPn7iiGNwdeHldP
NJE6VS7z8xpR/S34qu6wPqVcqFlPskXI5DVY/PTBcVWmmd4dzXzev47AsjvjVFaaT6dKUvKbqq5n
KTRzCJnwXVD9lXMnlWkGyOAglc+VrIVpi/U/gz8sOcPxrybdLM/mzqgjBss70Kg4Xu/mGiLBjaPA
4kPoEnPFyLq8HGKxXGUH2DJMSTJv+MnaLuQE06UnIRU8o6XGKMm8mJbssfPEPeX+a2sIq3dwGWoM
GoQlIsjJlW2/jy1vQ8zfKCTgyTnWAmmyfELnZNA/aBiMfnwJ6Sr+UzjuGQimR2aB/MmN2Hj0yHkE
/iQI4gcV1Ns2XJ2QSAcpPksV8YGOe2Jl2X9aU8+xK27BgnbVCC555h+8TXH4okoNIAQOa421IC1y
gEShqn7dwR5K2ODXDrkxEwfIA2eJNA3HlkObmF5O9Wucj59Ben36kG3TEIogdmLk0zlFsOdsRcEy
INq4G9+ErAfFK0xeY6UEHx4/G7qHZbiCfN7HgsC76zP46gCNQbgKx0WskU3MIcTf7vjar7fmqbLC
kengT/BvWEpBqvlhJQkC9+wV7xwkMkkm9DGLVcPWHrE14aQp5W8k4JB0j7dR+LhtDYo9Gva02EYm
YQh7BxDmMh2d45Y531iv1lq0k2gVAsXO2S/JIc4+LGo3Z4V7sbEceyo+GLMwcJD3WEzJ2cKI+tCf
tqTONBBco7/EoS1i2R+lYIr31m3HgQnf4kaAhnWMgBG3Qn905M7np7Ae5+WEhk6XkEIY2b59Fmxn
1P+d4vPsgCMfzUng75lsSy9cOpE3QF8S4kFz8eIa88r4/CgXETA8HpB8TIiTgaJhrsnUAPvr+P22
al2BUd/tBMEwX1wq5ioLDs6q9aRAzrahjy50cDgIMbpMWOJYsz6p1KnVwgPVz/13i9lMID4f0BfG
4H24u4YVbNbcjTk9Z4xfuOL5ZpSjlDGvCbZi/nbX1973dWPc/J7/kQXPehlef5fch8bQfBCitU2M
3hZTgCjpIZHCOmhEJS+N0steksqCMPGexNuFPAt3jX1R+SK/W8vYSd7Wd2b4zmiBfs95KZVwtvVQ
XugeK4gTDO8fnwOvDPySL0R0h1XMpVrau/g+lM4M/iEFVoKI72f5IR5zTnfOo1+2KCxdkJh4GDWU
oIo30RnrlqnxVNwtzZL7VVhp/JNroW4LZzXDGRtxSFOxEctp+de8TqTQ6yDPhZAc0/yWzBYAvqVs
zkRzdmtEFMuBpHnMk9F4bw+1n3P4bh54MStmFnZRukeZaj+89LCR5Ci5NrP6nWID52JNEDnmTBmv
xYZEiOGizvKMbG9Lz3rIJxtz8RPVjdXUT0G86LkTH+l2ukTQyduRQjdLWueQkUMMThjP3/NsOpzN
TkqB0PAF7Xt5TnCjgiRItPctxOFqd174wS3kkO1ws8yDplXQDe7iZeSefqOyNriVcHR6zKFGdmC6
SPKhkN9t1Zbjp8WbDI/a32eFiuER+d+5jIajEPoX3B+DENsXPCik6OMdiz6HzP6JSgt+b5iSUYpF
dNkAFCGvxS3KWnAbD6wGwIYNnBNI3mdhm1kmTJKVYJJJruKG91OfOg2//Ut9EtiLDq8D2sIfrzgs
5L2JCYYNZ6Kx68b08FAStHHxxCSV4V+eWmdvZAM+9O6DHI6Wu7GTENKeX9QxrwkrVVuIjEzNwaJu
ZKFopW0TZwep60tW8aE8iom8JoLcjXPobQZzcFjS4aJjBVx3mAlgAjIsHJeVPaakl9oWR9aJ+owI
WwFYbajbbI6uMRz5To/sJjuKnOE2DFSnXbRiC76/MwJSvOC9d2JaK6sUmmlKB8GGEqRI+0fVI1Fi
AwzrhPSorGFTy49fW2oYydtDWHnI84VG8Ir3+4l682Q0AxXBdcNJKrehJJVwgZauO7yiZi0iGg85
PruUc97qhoY6P2zP3bE6GOoD59qku61w7NPqv0FWatqQn8Ui60/0h3yRCRQwnUhSA5WgdbEW2e6S
y/9MZca75aKnJcifqTyK1KvbGz1D+VnUl2SUkigmH+fdnGVDl64Tdqnu2nF6SpK/pmbAUTXClX4K
J+LTVQ3xoxGK63Kxova40/jiGkGdFkPWOPP/rZoRg7ylp/DJuKOMaPzyGu6fMWt/69CGQ4O5iarp
PnQMLhVj/nk+04THUSF2MgtNb02X4o3LeNdV6+0aP2Oj+B/Xkf4tXsZA71NF6KzeEcKZ+IBAJ5yH
M6L8bslofiAG+KrInKW5JDa82r99Nvw+cljY5DXFHB77BLtZpg4LidJcRtjvMWS0/BZEcfgsI1I9
DLxqVMZHrK2ihmRRBPtXIcJjnROybF7VtFceHiqMMbtzl4H8J8aqu7cWZpttopCbCxLutRtLIvAM
7guRUROkp6NFH50U+kkh4yLMLzXnCnwfXdN6mAyKbuZFXwf9PmQqb2vLu03rnjDch7q1ShgZIQG2
KsjI50cICKq5KWm+fOVHl3HZFOpLXpE+tYuh3R+CA4wBSXd9PZAnLBjW2Vq25s7U9f56tA6KBR6J
6YIMELWNapNU1BztEWYUIPYc8XxHrDeq6WJxcRlxR/TttaA3vnFu4tkj5rI1j3aPSbxw0hj4pkev
nfzrZj4O75rWXUDZCqvbA8lJHmZOtYbfpytac1BEAnIse5CTEQY3bzkw7GtWc1R3r6WJL26Uehz3
awhA0OujMMdTR+5lM/ZQQw/SV/Z/nRtgHBfTMsR/qXXKovKrB9kH7E8d+q3XCyiEPaPI9Boe2g10
J5ld9+9ujcACrH5UHpUZ8dTHJ4fwdp0JVSPNY8SNdW9h4trDr0QPsTj9IinM7+eoPw8AqqzeHD2S
xOKtUkWIAedNH5Ehy50OLfRwtx9Iid/31ROsGZebnBe8qH5J7mJfZxUBAmpKI54Rng+kxSnjE06Q
13VWy1Gm1ReI388atmtz6q0E4SoBAfEVtNmpaERr1izxvji5O1fvo/L549X4L4BUaQzQrxhWCbJ/
YZqYC+rmO73q0MjAKEVMayu85N/R9ZH7AAy5bJGEvtB/Ud8BrsD/yDHO6I3WKwCVyNzzhA24uRbV
ZoAD1ZK8KlhwcCDiwQYGdsV6S05Bt/UlVIDdO2X4ynLQ0RojGOb7Su3OlqOm60FBjDHloUsoLO2h
2Gu2//X7aTtxXm6btxXg4WcEOzgUrLWU36OCG/lVbYR4Y37Ez11fkfg0vNEMFo3TwBYJXxG4u/QY
78LOalWwvitjBPZ/bIpBI7iDNqdtUUgrmUrvMFqxt/ouh2mI49jnJxWkqf2f9O76LipTUocUCVbQ
QVf+Ntz/BDj8tEXgVdR95VlD7fXEt7A2cxYZbUUREpjkYSP5burQDzYVA9z/Moskly+Tmc5wqYYh
jN+kJLc262+pqpRdX44LLKPQYPucioHN8t1T8ivA8WVp8iBgDUJmiEZjCUfLzKUA7h3nVrlY4lgv
Kp5cxaJKCcnwKfORGSC+QfWDowHePxoktx5AM8f0JaOSUG84VKXv+Z+J2CZd98HCNCQjC4WLWd3Z
gLHBkp+yP/BI5i4MpQxFdm67OJewFLqksFAz3HsWgeBf9TqX3eCicX7kH3fih9KzEHOxSzZbEstu
PdudFbvUuGPTTj4oUCfXoRMN1n1whkRUKvWLdTU7sd/Sh1AAUagsWQtn5XAI6f9e854Ucr/X2sLK
A+lp8Xcda6Trf1cjeOZuNsYCGBGKrwWvLfg0t7N6/jXDV5V409yr6vVkNXo+2TuNTkLCmh7hNdjp
/Lj+CyHr54rKRyJ9PfX6yvT/WDPDw24OpkXiUvBCnPl/P+UJlO3YVe4nuMlluc5xKU0vmAHRgVM1
rMaX4URqkQin9SGuwjggKr+ZjndghOtAj1DnLn29eGAKsksgx6qVcXemoJeUfn2cZFhQ/oOhDb3N
xnG/CAsu1RmU+IbLHe34bEzo+xnfUduqWNhXpIQ8QEq6OzOkHp9oWU8kS8m4oNm6fKW4HORzxHeT
VsiV+uMrxpyD7ZQEKfNZyeZca465frt3KeHOD9Czf7DEJORCQ+4JrwgykbPGziI/IhKqMzpCXYVo
7k1zqnuQMpRTCwaS4O4iFBWGbc4ShlqO055/CT1EVACGcgOqyyUoGxJam1J6WCtbbm05on3MzFtO
7YiO4whmJuFlo+754g+XU5v4OaLfnA3ZwPCAuRS0Hdhrv2Gr7uTbEnlg7pJXaznFCa6zb6JUX0vo
+jFU9huIXqnBqlw6m3Lg5mxoS1FXcWTIbQfeMdmwKYyPE+vR0xrjfz8w+UwyACTpdyoLWXJKFwNi
4iSWXCTOkI3/YkNqr0rmOezJNBI+gvoiw7EKEIBjN0RxikGPtYJXDp0SzJ86YA/zRwoQjxyXzzbE
q0gvuC4Nmz+6H/622AMX/S+63VWU73i5LIxEgEVrS1pbpZ1rsaFYhPwvuEM80/ygWsFcw6oTPx/9
IS69FKJj+bHZN2DpFFE1PF32kGnSrl7Z1jO5854pYCmP0nrBb8X9cDRfemC2mzQMPmpTiDeXV20y
qeR+O6cU0fPh2bOxqyxXUe2MlhuKABsnq7dbslr+AFslLNmx6XPIJUmcFJ0I03n9gudrBg7hpSPP
ynkejwCevbGjhH9LLPFTKtZE+zI4bb4+b1MhKscZ1p0zvbkoKyMG9a35OClMjVnbt2mAtTlfeF0/
1dy/F2kRUa6wAT+/oJ0BFcbmgxTrNG1VRtuCkCd4r3WNU8HcbsZAXywfiGEpCjeFmkSk/0TZbO+W
xY+FZlYcVMJYYH3xsVLJuZ0ptBYVwijmg+bvbLiXNiwhZYmo711nOyS+Nh2tfoGnCqjn44LVgjLr
TyAjVeMWSEc7r0V/TU9ve5bJAj2mzBga4vvgdLSxYL2fjbN5Tigjx4oPodXKfOzohgQO4SFTE9ig
Nrl3IkdaUpT/Hp+9JitabeP0WwxskZL4nBVpE9sZrfjoh+UQtMSPKeEUj31qjiLqgCMDiBOMW02g
w8WtKjriPFcWf2FfwrX/GoMje96sFZrvld9tUZYpVevgRzEpMnZT5d6CmyiCqMgoO7rJpofAskod
Qze2UPBlCrNFGSHuWYHsbtirOEHP+mzDXzfKGuqYTEAY8aM20hMEumTqJz9OudDr5Muwtb9hWqOg
izwvPnTNEdb+3g5X98hrPexbl4VpHcrrXjbqj7FQt73v+wXvdUTWGdjiyK02wOzmMPi6rSUPC5ZI
SlHnQ2ogghoVEEh1/1HZvbMFMP9rYwUklgBR6z/fR6ADF1u3OmZjxH7v08kO8E3paxssUDwelynK
GwZWX9c7gMe6BS5sOtqEAYkv2ZAPiweTk86sQB87lJs+dCSh49xCQzp7rnyLuR+7pmSdWt+iJ86P
PmUPb48iVykN1o3IihuZRaUUS0pVq1Ap0nWjc7iixvfVRwj+/QlLCB2RQuBsH8Oi3enbM6AtzDdM
fBX08wSIvRzTAA6wQq8ixmfgPLI9gGAXvmemXRyNk8/RuB0LEDVmd8RDsstM8JI5Q5r8ZYE3HoPK
Hrn99ms/0+toPIZ/6kbYFMfuNVJW1fkb/IIP47p9T1a4E2PjHGjsvQ0nUHrY7p8faYsNZZCbChiG
YSbp7A8J7GAGAlRFkWKQyRaDqgWdVTudmrLe2h4pUlbngstMLe1IRjq4tDI2qvtCowE2uw8cSr7f
H+HR/dZQzJRQEjpTrcFGw8M9eDhpOSiL99wC4LOqhJFMRR40R9Xl5LfgSVcU8/dvjwkzfmgT9M2S
28upnobncGy3u3GGSsb/s2MnCyHTWf00rbTu3ZKJl1af+PPrPIHdEMf1+cg6EY16wfwI0OIrHX2d
HuhOkkdrgjQiYhaW+Z4RN7+56qmirv3tPkkXTq84DTXeseEhGH7Rt0h+IXnHR5ARAlQUg+BGcfEg
7j9G6RPex2Mdss6V+xIDF/YiFKksu3mBS4Pt71YAflyQeSNUp23PXNqJWmQB0h4zrOpvNCah5pAw
aFVL9L+iACxaLyGUspA6+1Snp39XmCfP2p6E24kX3GrCtSKvDuiWGG6t7TJzKWHQpaxJ2Oxu5TVB
Fm/YBXdlMpTDIdkkpU6wPTPqTST14iXoMeYZFmlV0R9nwDof6o0dt92gvs0vLI0Fi74+e2TcSiUI
ishkVOY7XnCIYau2nRtbBLUsbPrs1LdKaRmAxj3pZj5CeAmsU7nFC6Ou4Ge/SyCc0fFhe4N/obr8
mSpd5qzgFqqWXNpUJyDiqLb+pF1Hj5unRGDNv7yhYiuf7HRNlu1NiTrXtoVumyj8Xit5g7crFHUl
EQT5hLo/W4ELAP5hX/iJavg23kX8zFLPzreM6M8GkzdQvNNWAh1raUhZ0FHLcL7jhl74bkcIb3oB
QGVJU0rPsyCPtG/jr30yQbQ+BHF2CIeT2LsdZJP6QWkwwRmWukVuinUp3yUp6+LtLfV/Yc0ofHUs
IT5jEDhyETAzM9J3TWmQR/NdmZ9xbIEnYSfccX3rd580EsSNzt2Igr61zN4L50W5mmTIm2ds8kgo
97B0IqFvOy1fROhUd7czRVQrUJif9YZV/yeSfji4p1pSQ27+gJ4ngzbtRjIOWNkDgBziqh5swjfh
nOxks1/fMzJOY3l8usuBzOweM+YP5llqEuE4NDAHNiiVP2ZHNbwIAqfLGwrzfY9uX6Zi3wIqpsLk
Hx5uTnAM1+9q7LXUjJJRjYROrsKSHYostMzm70+YqnH3QSkgdVDCOkyMctXsL7V3iJiArQb8a7fQ
dfUdxdBoXkiFcs6xlPIMlzbT+b4LcXAMY0OS3E4r0QQIHB9Fobf9h5vh7mGjw8pU5FWoS6t2H9Oc
qive3/TJ77XzLLFw56xEVCSi0J4D348AVDqgWrhPoHccv/42MJu9tlZumbzvBNhnVcBxWk2u3oTe
jsUkkjFPAfOB6WNpKfvnX5AZJGzrRQTl8zeFQOnr9B3NqKNRA743i+jOto0H/xaIEGYQJaXz+Z48
TV7nh/YuCyVjsUj+b69NnAnLAMFoDZnB+IuGPvkuT7/CItwnFKouAIIMoUUawCPgBkyGm3ON1TIS
sgm/58kyxw77NdNCZd6L3D1mXaBbT7HXRBdXVZsH0KrpXgAWt4wA1SDsO5OK9+eGprU46WnneXQy
3dr/zhqR3UdZRle/2GYGeBbG2mQFjkB2uZK8dHbe/m4vKHHP91bJWoxLQjxJXVM9/i3JQbMEFWDI
w1vGSAgQaWGGKYhHbL7e09wM4udKJFQlOPiiKgyEEk9gzoBHrvdGtAB/SrRwwDbqnUfw8Ad1U+W7
81IdJaDbyumPxsyYzFxTCScVGFvVqRIHzGfDXcRTWDB3/fbSE12sqJ70+jWV2y6WdbiyqdKq8MCD
M5iGGPM5KGWWhnvQNs7mLgLR3r5XVSJMeX2FOUdsMruryVSrYr2/AphqFctjPr9k2LxIoByoFrbH
gwgJW02/D6j1SXweZFRl7ehJ0PrOLFcSFAPEOJlC2kw3Qdast+JC0vOmfcvGeFc9a2L7YsnD0yMZ
OPwSKeVnpRyPS4uqETFIJKB9NvU6Cnv3N2/n1A+AFwTaVRu3EC4vwaN1uJdwSYM9/Mo670Qicd8M
5fInF4llmzBcFTaXyospvFAFK7cPkyGf8Hg5O8rIgKCHRBxIlWWE1BoWmPNQAVdlfzumn9pKRrUz
X8ohmkq4gObgYZVZ6dPx3Lk/Z+Z2kX1m0GA28hVCDb/9xwrAskmOZBuj8vjEt8Hu17Orv6pkbbvx
MXXlCFR9TZjJZPMMp6RWbT3PtyHF/e1KXeMU6j5+UHB+Yb/sao0r9hsjDY+zhLrHyVgAblU3tCSE
sIH6nmnVtiYJ0rTUf1rfWhFQRv/OKrfdCPit2dR0JGi+QNaFJUkWG1ETpeNZJVEjAyV+d1Ov0C7a
YUndNwvQDGxsrEQU1LCs7Ypt/MakN39eC7FlFJUjFJmrYtgRZG4Cmt42NGpBXc+U6IrMw4LoRAHZ
ZwVBHfUsAXvdb5gc3EmjdxZ9IZgdj6Ksv+udN70/oJcKuD9csPR5uLFPMlz2/kL8zRUdETQw4IqD
im2p/6CjgUV+pJsiCkPczSdMea4rluD0r0mixkMNjJuF1dWd9nwKIBhIwOK34gZPcgVWNf0JNQQW
N1vCrC8ojfMlj2kqTLcYCtpNmv916FfhRZp78iB7g+mWIuaBFo3iAUVO4KirrtE/0YDvgJ6cURjU
yal4VRgIU/r1tKgCRQVe/ybn7McJkOVm9a0ylOtwEUjTrwZVHJygQR7b/1F4UziUlEdsLw2D0HW0
GPuunIhIdUruz7E2oQYBkWxgrC588QRIekqSvZ+BYdpwY2X2zdnLZTtWqih3uZnvJkDDlKFGVRWD
yW0SqG0xyGJcRgyzHX7enda/mPdaPNXLULuRlWj20zuy/k31GUliTde7yEIs4aB+sA+BSNbLjLyo
DGostteHL4aqnUnqZgb59x9z882GwLUZ9CVc+SHDVGwiMvfdp8uBCsZqIBNtp5G2v+QH7HZbHrtu
4jAxdBCfPUApHnAGfCXxAbjfgeZCYHH7zkwHuXeouBaC0SfzFnFIl9QZh8vl+x5cCP3kRcwVkSSn
VSYe81HpiiE9+kn6Nu5Ts5oYjEUiGbUQX5hBEfqhdp+qpXgvdrB+s+7+twnFc5HWoK7zVnrzMQeJ
XybydMBtHqaaMi7CTE3y+5pTV1F67JsiCz0eMiNWvnYKt6SqdmGYbjgv6VH4+e98w+Qzu+UW5t5q
bHFafFxcEZJyqHa/c2dGcjRqpgVMMaak3IKiO++7Ck2ZwzdO6iuXfh0C8ogZ0gw0t0JFLB8nOhjE
+4Mp9w54sxqFYMNLRTOezQUykHWiYWKPLKdU62h8D0ssd1s9aLYA1fmHVzuxrG9L1A3elEotXMm1
lCe/BoXjUqQZnMtY6drBYGGUEBlm2UEU4HO3GUwYmYmFSc5fxMTXbS1V57UjEVDzEbTewt6pQnQL
1BFwbJDDD1x//mJDNfUWutWoxE60cI+5rYbjh49X+VEPwB1e0xxlx32hZQOug27N0cyOiz0vHXfM
SVAU2X3HqhvtSs0G1oc9lfELsBC6eEpoX8NLV+1Dd4zKe5UiMLlS7eZKgavLkiFlfAPgUkr+gWin
8NbrlpLeAXabWNzYyFPgW+FchZbRtMbD/mqrMv8I/RkZKNv4J0cG1H9awk+Ejya+/hGerREJV9W0
iWtiePYkCiPk2rP3KmRgHV5F14iopnUJgi3dIkRupejU7zzCYgYVeQmEA02T+/wH0dQwRin+dmow
NJg3SBUNEwZoWXtOEVqLPLAdaKvD+wArOkTS2GEbPSpXWAnkQE3PvPDgzmrWGzqewVwWBy83V0Qi
S7/dnTNgdp8WpxvCVpJTps5eb/5sFWhcQacG7ZVwCvukRssoDQPbalUPtrqeFMLZZI3RmhvMC3mL
V39IN0dwFLhlttT8zw4wPs/6De9x+YTIRcAWT/Pqnes09Y7VzVK4FTKkcJmIn+g6hU+C7Njzj/DE
V2vWCP+rretk2diNFqMg1xCdnnIxMo2DUrxo0BijsIHUSAids/WyPDtCou9yfdDeEyNdMo/lkepG
qNi842QqO8dIpKfwNSsfYhCbJ+Ey2X7FMh1LV+rXELfH2N9mYJgvk22tQbRUbZlKugo6F1NxHD0Q
9rE3Xl9DVjofD1p7Y4PH2x5rn6C+aL10xTmQZhuhwnAHmdVRHEsK2pkNunaM2hVY/uH9ECzWBFQ0
n8CjopO87IwzIJPyi9qSHrm/b0xbqJXx2s0PLgN0sKVxRraTN6YN6SqjzHcyw+Ly/0Rswg7qhLx/
mjGaD0+Iv/RTtejeplhAcheh9AbIyonBtvxsaeX+MqKmvAxgn0AskYEWWukdE54IzkId2UrmGL2J
wIRVFZEv68B/q+lrwaO6hpwHvxNCY1zzaT3zvap5MRy5QpkO8P3mAcsHNoENbC2XfsR6KMPACTrX
zkRBqeW3SyG1Y9c8HYiZPDiFOusyKjTDLzFHi7gb7Nwb7do3zVD2xzbaCMJzwlMvJPduVbKT34D5
FCI/QTGNYpqWvxfKUBAAfB5uiLcC3whaSoGh8H9lD71kJxKc9jfy7J82MgU0GqRK7VQUm+EYXJpq
D41dtcztJDeU9c4l7ezobb/wTbwdW1eC1Ba+KXcVEJ08w7gFOP8MW94IMNuhO/SkG9gxK2ni7jz/
JkZkeeCgvnR7MLeE/Sz9B+rRwmH8j4egmgCLZ1Qe7wIFEF2SwvOJDK8T1Az/8M3MTud03vvVc6zi
GRMgMX8d8EP5eOCafms7zBw5Ojr8PE8i3UO8odNTrSUhGtI9S3JdX0YhhvxyqIkUM6t0lLRwPl9d
EL93Yzi88S9cMLyJo3edmG4xtHlbJ9dxamJ6q3g1b4egQxrh6Mpfnd0gJCFieIJttEFj4qJOSCwz
+zxnqdaWUcqI2kBcp3X6IQLRlH8iyhy9hOrI2VoiblwamalXbDYRbL0eBDNDMcQ2ovRvCFgMpMYx
jX3CxTrkvxOLSv1jwAqwTQV600LD5fx3+Bu2cszBgNk3ezuJc7BwdXnLMO2yi4K26sQc1zyOvWHD
v6ukOebnvvz2lH12ZccHBEn/O1bB21x47bjpdVyrRNn1BrRyp93oD12P7Rpm/8fz6fExub/YTBz4
SMAq2VdzKMJadQgHtS0bCx8IxyADTI2JtizchkEv/TP3PU5xrZPa/d6L4Ky6D8UTWACmtAhi2UXR
i2yWzrscv8fltuRqC06WXHm3nFTPl+n0ulfM2DuSKOlpA0QVgIYllywgARr4+I0ei5wDCjQY3Jbw
ghk50ILlVI5x0JDEgy9kNJ3oL+DPBKXZkfzG+pJ5ODjD2yEUs06uyKoDXTx0NEW59tcmg6w1r4EF
v8zuL1LyjYF1sMK6B39FVUScv93Fw9crbDSXrGXoJb5KAuif4i4m3g2YVtKHk9er2GpjsgMyuqP8
0dlSn0a2w/+eoDH0BHl344WXPqAqystyby+5dnZU9Q2TSNqStBx/yNetFlMUKxJi5MVCfZJc2gX0
xXZiI+Yo069YvTmLOUqBNWE64DPkYW/AYkv9EMNFp0Hjw/Npn2DtccMG0Mv3N0nPA0GxrEllHohR
xtRBcj5xzrYloYVSyr7P6l2NfrK/m+tlJ+fyaxQpWMYGvyBIMYTCG9DkOpQRzVNahRy6F7RRY8Np
TAxC6AtR8AxT6YOWIzs3ODCwkzncX4OzowmBN/Xi6MPcV2K4eQh91dmDrT37Gmb7TfZJWTpOpksr
uDOZlH4ytTRExaOt1dOqvXsd9zTT+JXv9lqvJl6/jmfITHKH9ZKcdQOaX8NKVra5i/K1fzHvyVPa
WlDRhRLrfTYRbAXwOJJJKwdQkVN52OaQf/TBa8bEhvcbwK6JkJ8wbQF+GbIAy6gbdTyvGh5xFupf
N3Z2PsJh2tM0MB4Qy+D7D+WpMh+BuMKWIX8Qjj8vw02Y+vywcl6yC8xv4DIYBx5az5sJ4kPCynzu
rfmYCGABCTuxyiERv5u4lXlQMVFQoltwZasLyiSaoI8xJsAOFHKAsCZ0hD1xFEjZu7RZYMFLgkqh
+YDw7tHE0CqgD9I0ghupTOTrpJg50RVAf2SvFVCmWJVKbg5eHp06SONMI82+dVuca9GnaHrtOvlx
BH1TPmDz1cs+/0wotMsQNyB7fpX0+X+65jV/Y5CJg7nhdR0i6gys8LHlaMp2phROeCWONA5TH+rL
Jq5qJQSEg80dPCb0HvQ5sw6k4ZvXU7KWcC2ZW9AY1JGV1RSqS0CVlsTjWa3D8cKbQ+5a3mC/3ru/
njBu0mLTJrskdkSeGNuiICeg6RYtZzOGn7DmAbpJ6mBGXGbtu7BZX0acQCoQo9sfAqsWes8876/i
EVmxHJwaIAYu6f0BbSRoeDk9fKXs1AXsqlau/DKvU92Q8JSBWdeXk55/O9Tx/Uto1RySIGUlZRAZ
yBHUFnjbF8uCq9worE22q27R6XvP4PMGMESAsysQufSlYC+8tFTjomFOi3E4OMcKB/wh/WB4jf/+
gOaRYl4vhP1bNrQjfAaMPXlJmuO95a8X7E2zhHcH67OB9Qkm7OQraAxtrx6I2ysIXZqhjTiCvRod
EjOHN1OkZHvdvVQ9m+Ked2ehlg1eHhAm7DAlgrrevjUrS6Bj3sOJDFUG5XQkBPs+CJVgOssy9w2L
sOjGDJXroQ/vsG/pdjR8j6PuFbCOKUMF1DQ1DldN2pUyZCI781GCQEo+Y3aGtxfXPbTbuj3cjUZA
Lr9wt+Mi4YXPUTMc9fMHnhs/rEE7FfS8uguzzqRDPtlNqBLfCoc2huPAK3RSY59FVpm7u5QyP2J2
UMSCZCQ7yXpEWY8yNrRXs94EAJMCUcbzq1n2eIs7rIS/k4TyGOMUh7Rvuvnmd2CvR7h/P9H0ZRm7
fmLD2ctLZZ6BiU1LfAyzqeV99dJWFWkkKeAF6zJIV89V7kyryCfsw60BWJ5HKKic0z7j3E18meFT
57pJy+om3+DZac4qGwiB0UhdBHbJGuPq+yFiQ1M7Mj1Ojm8kLB8mWKLtrYUNn5Hp/CAJ5hHz0RqG
IGYbs7TqxsD70BLumbcwu6qHPyddocpsEpj4WhAH7elNBQcnZ5EU/ziJSW0kTnArSRmXSKUW2wp5
YxTUG0vX3g2Pgtqhciz1nGnLmuvxLS9Mbzc9bOCnw0l0Cu1G9v8ufU85Nu2zDflp6PIvVQAmdKwt
mOO1WqWHncq7b+i0mUjErNdfopGaXd51q+gCv1hrSfIMqN46Rrdv7rpWF9qB+lSZXUvyzTsG0P5w
LCilg8qacfeW6yQxy4zCcSzeFcBpuPWZMkLyvls/Vlm+yw0MdMtfNM0lCCSvMlNXjeaOyy/2zquy
CuvDQ4GYQHBBiHkOHrx7nIS6v1tu2hDHFxmQah95R7prqvPRGcbuOl6by3SfTDRNmU7rNVuqIo24
tGvPe4xg1qxeWS2SHGCmU3+EtGYairm0J5t68gD6sATuo0Re/TeW8owY8BWkoUJnoSqNG+klr0pN
59GhNOysN0Lq8E2XgMqSy2vasEjNN/V/+JGPeRkZutRGx50F/OeAoWgrd2QMU5MswqebW7bDIEU3
4b0jrua7KfKxYJQO4dPlbXbwGNfTuZNjHKf2tSIsei6zMfbr9y8Y5vueYIJGMVb2QnSKUfP0SI7q
VMbSZNbZi+7lMhLGNnrAr+EUyJJPXgC6o7gbaQYt8/NiTMpjKqLyfvZfAQzvmRJo5SAIYjmJyaTI
BWGTs/BvDyH1qU0GeWMM90HjDN58lrpyxTKMnQH8Q+ibPPfWt1cqkeWdxusuHiYXeVo9SMYXtEn9
H8O4FfxWV3MNmTg0kgSkNJBNHWQw+lfvbevv4tdZwlgLMEPHFrDfkh5pCFVcljU+0th93dQ6gKoJ
c6LXjY10czx5JcDanPJu21Xw48d9cXUe8EufCC0OKswy4VZaDQl/tVqNaOgzbsWU4que3gt4u3dF
+3XT1Pq3e168y2WrdG+QyUPundNYYsqLW6YtJI16XdARhFz7BzLo28LqqCPDmCh0V28+kRChhoei
0U198EqyEYa9UMssZNn+GC85oLlU7kYBNH7+qLQOxoR4tou51FRy/a6cM2Q85PVc7jWAx+bVSek6
N9uwB3cjybLrziIy6KWt5duHvpHZ9QqCiT16tjd/dOH6ZAxCt/fubVpADn/OKrd45fpIxdnMw+Y/
mJ7Q7scfAWcRfTj1mjhdasq7z78viP73xR0W9f4ZnmCLZx6PmVG66laWxMKNgSN5l7UmZBZ4LE13
2IA5r8zPct5i/r9teVQHncmyfJTtGW7fKYJdIB7REukNcyU453SAhC+K/b+Gs7DRT6iyCHTmyl/8
Wl0R4z4rCXWeuUsImmBQFQB4PB2yD+xAXq0UBlWlkf8eK2OG9OMBUUFNg/vHxFcmAnt+/y5DGqez
tIV35mCCamqITm0J533viBK40f1KFVQ0Mhjtrd8KovM1ZekzxZcELu7p17Hpy1ffabSdMesxAR4k
XUa4CmE8c1YgUhHACMSp5Ix5OJitMTswGRruuEU1+UZb1Eq9WkKNNBzlSa9vm7bLNRpGEOdSPPkr
j+twmLQKedE7FVB8oAcBbMEDoeejA3hE5UO91Bts0x80JEc7NSaw5/6Vf4nIQeKVwOLv+CSKSZ3R
m3OKtCfD7F2V2g8vcodV8VhG4b7oNlkFOzTyffZ/rRWDfJv4zSV84ZDk0QkMUPWLZFyEo8w9jY6S
BEqu2q54yZH+UnCwn5abodRXOmlFBwyiIMyxD6WG+GFW8vlCTNQN+DtZ5FtnI3Lv6QU6FOL7EPjv
DpVbYfd661xhcrvvkU+9HL3mRRuuzYA7igfhYsP1rG93IKOS1/zd+tKh8PfkBxFfRNRQgE5sKpCm
O911wiDUuWnnmREnR/jwiBg/HLN0e1zXg/RHbauPZJM6VzIp8nPxb1+Ab7Wvtpb0uLNB/wPozDk3
5iT2zwE4BhqfXLHOplFXjRLd6VPfxg4RcKJEcJI90QyUD4GMo6KzuWYiPIHlxXkogxjAdiFMWAcd
jz7Bre6NKrSNfoMfO9ddA9eoE73LnbqSjPYa6Bh4dIriQGRGvTJxN5G+F8A1Ze8WSZ5nN7yBF1QE
9Sw4XgRhbocovCoemQ1h7XvpNlwHszGpm9Hxc+poU3FirDy/nPPQ9gmip8BSE92zvAIel5uK0oSh
0VfpVGMUCcRWGl2MqG5sFixIBsRQTS3i6el7axyI8bZkH4Fk/wMUQ/aOofWdjrMRE03UUWD154rW
yNScV3rDeHT0dsKpjn6MLLdvDUV2XrFfpGLavUBugeYK0tWuEhDZvjY72cUH3u6MViDRVcMTxrON
UWA4RADQVj4N9lF9HOjGfkUGPsIgM56SBbB36CJx5joxGEZtIZZcAg7uSLpufeTo1Rz4ybZx5GN8
379updfKSOXjKqEkCay1pU3A5HMoV+EAc5mGNC9JHqjOdIMDdhGMNLD9/LZIoUScZvWutVcLm/2t
zDJijSj3waG7eYSD/iS+Sj0Hfm/ecEzqLH1onZIJ28w40MSS8X+ji2CeYZMXxCHU3rHlIBNVB1l9
RJM8Uj8gLjQqUIBB6UvVnlKkgbLVYoeSKav+8Qsrc8TaQ4yjKS+2TDRh3AT9n8AnKbjkFFUJQsQ2
m2cLqTggHAEE9K3ms+piS9GibtXeR7BqTAzbUPqBbopP3jYuTROfBOYIDYDQjH39aY2Q1mPwCmL0
OiGueamk74tfWbtPYgJfcXlkTVe8mDpEiuVagWEa2IveFGJFflWgBOsf3ERG6xLpBomp6UIOqAV6
zHsVnKO3DxT0FXdjRRxLP7ELvMvAglpBBTZ5yKTIYJVteB8BjQjQAWnLHZVWwf6tehGpukCEiKs+
sgbQR+HD/J1cUaQkS1LP2ktuWsmdbKO4wPRgfPLpMzX242FFY5t83PnO91UcLT7FN6woQ+i1zl1l
XW7943lPM1BIglvMxi6Ud9tFs3arTPbRt35J9Uj6IPnA5cEHaTnWqXk7lTUH1Ka6SfOdsIFwE8Jf
t+XCjuKMW7PYCL2UJhjj5kb1jpiCcjmhi+ZPqGaYM62rcN6i5TdX4AOgQABmKfQ4PjQ2edKQznlk
3J0TAwyQbSguEpIA9vuMLwEibaB4k+ULnpITHKJnnHjd38fAzXHKNpi5N1qYR7bVBNeU4mvvzugT
dFu32F4ox8iNknc+HTwNsgIa8TvFuPausbHUroFj+NmCfiSP9w5lvSlO98NNyK1EE8Wa3hH8zq8y
uIja1L0xUI3roKAWuzcRec/gFCSDthdRATv1FVMAobII0FS72uoQAP3+e9sz4/vS3o+GLnt01T7D
v7+6jZy7C31Zqd3XyNo4d4Q3g3UGtfedobT/1BWD6cvnjesA1zAL1h1uef/Ihx9XK3Oskz6hLBbp
XhhcvZqbH/k2vz1RuqLowuHDW070P2LM1capwk13StpY3cqLWIuC3IHRTWbIhbgFbe0xpUdHh+Y3
hqQ5VoCmiqEW3WWGRsrQH4lBigxCs4emWpiSnO9E9VVmNf4/Pz02kg6UMwyduR+uDWMg4OF/tg76
ckR7cf/LcWd3D7dO8hw+Ggi3f5enoq+WNR/yQhoH3Y6siGB7+/O4RkLSv5WdR8ZB8Mx72O8kP6p0
OUz3ZXJu3do39XB6pbj1ao2O5mHWFVFJc3dMtFGoODO4kNwk4OWxAbBCbH3wR9It49ObW/crVmd8
hXyBNGXpxSi3e/rCynvR0vbzGOnOgJKu6veRdq0u7FA4iHpkRAD2/Z/yDtDySDt58gFCh8YTy+3a
/FxXW2ZRA4HF7IKYn42gtloisY6lqX8a2NGdmijZyFMZ/yFcHxGlTqE477ksVcgNuylRjGijmZji
Jq7EhJGjZ7BIFqcRUB4+CUvCHh9PDWRfuUeFV5ItOzpG0ZV3Fxe9U9O0WgNQdK5zucfGfapfUW06
ePICuKc1G04kRDgI+mPs/gAbca8Zjk8TmrlA0f1VbAR3Bw0o8+C7gjNNinlrj0Wy9I/NIFYfak2E
v2wVNur/C7aAsHajp8oWQ1Vhf1ZD0x3Twp57LNpK8+Kpshx9qDa5kgOyOuXUIjAg6Lv86EKO6Hut
6FluslLb+JxkjVuzsgqv0WoRhmG5XHRLPo7pisz/ZwkPtRoWmUJaSNbrmoSOBfXoktKm8VPOoc/w
sLuCK7jZckc7mmc0HXDMPvTyg3Pdq5HXfmnfKnqUnCigvrZM5lVyMf526bEmGAjdG47pETLWXHjt
iCROPePRGCeR0q/jxqrrtoo0MsGt8A8L5rUkYcifJlDe2KDOOUKX9A4PIrXS35qQD44FqimhCRuJ
1aRAaFTEXLKWTsCraT7eiE91jt+i/OPlEoJ2XLv9s/T26VrCapOVrjEVva1hAMfbKnFnTs0T6360
S1xMp9B0jsgHGLeAUECTRZeNZE27M0aUjS1mZkIp1OI50VoM1/knnxQ95XmDAHMGxKnPYK7AjDWj
qQOxaYrOWiz0gid/ZwohEz5mP6vy/ohoLE+h/yR73ZKUNQNtZ7NPj6MFosnoLVLwk8KZV5znh/I9
LYthBWag2xK/HHiHHt3WPKQuN5QsVKDwznR6alWeL32DZ1GkENGXr01ZaubA+WTZyF+FZ5iaWxm6
mSUR8H25phyn2RY32HgUwCEgIkty8kwSLzdQRF9zg/lQX1JBwnnkv7tQlD3N0Wg51rUeSvFUc8gK
oLtzLzWYVHdfH0uWH3TOWmmD08ouqAdNicX2OnsTOIpyck+WNtglzw7TL/3Mu1Ovv6gm0gi2AsUF
eRQck9oqldpspuNsTktcosQPIgyZZWFqoaf8VrpkUU4SRxczEkgcHfSLr3HP/Ekv/pPn9RHc2Y9w
hMcl7FmdB5OaSiamcThivGxJ1jjgyWpqPMNAKBknzGevamvXmum7VKL6vO7lefMhATyfd880ZlR6
0VDOWn+uYQ6dx6Ba7lR2Efe33MxzGaJRffn11qUTfs3kN0zagnWRdJCyecZ8DKv1snUq05FtH8G3
FeROlaQ1/f9KfGVdmqoy8igFqFz5vhhDB/aDQAATxq9rwQXJTmckZlsbmUYGhFHN2Rk9cLZt4WVK
VMdki4eUUZOtyPo0fTtHdcfnCfmn8QlU7FW4U9CJua9miLUwOs4aKjkXxAielzSHQcVAsA9QXeRd
FZCBSnos3V1XcwNK5dBKH+N073fl+ZF8nKsq2uUk4MlrHHb7B5P0IhZaqSvwqXKx+wDp5J3fWR9d
S5jrX86b7cmsoxiW48fojphVtHz6695Vx0q/F1j1lxQIXqjuWanAlhNuQtftY6n270pEHlUhcDvI
D0NzMDEwNWOH1aZxrYY95p3GSk8qCauZUAYPmBvWP8yyf/u5esaOuwJToddp4b4MGFq3Y5azLb6L
9FH2TdIlA/sIoY1lgG+5/GOwpQdNWdN7+964oHbbOCyNEZzSU1xXe0M+zjpZ3yU+pfCDSoTTwmu5
7YCLyb8ZhTAR1tp77rr0xPYqC51PsIGLBpV8VXVWOqgD1Mkgm47sC26WtjCU0jsrFYCCc8R8wQLV
eUg42DbKn9Le7gCDAc0wPSg1v59iLzvXKMIRXEHsTPgJGwLpBVPhm5YLqDzbJPdIdQQzTtj2G2+Q
sgunSJ7w2jDCuOASzApSrSDLWBCpNw1Aq3rdomhFBnaF+Jzmw9OO6dnFnNThfP8zXqTjZWeAvnJY
0kA/gjzniZYrv7hb2MFu0wtWio7XsR36brWV4AVkB5VSzV1OS7a4EN4Wqmw2giJzwuRzM02dix6i
QNHKEzRoGUpteY1wCkbcw0wMuY7lLSe7hm82ZNMytUJrt+sK8LzNIUmhnAFpOlPBmkvEcZG9hmyR
UzZg3KZIizG6Q33x5u5OB69tR+pwY2ZY+jSFch3hVY+DafyjF9k6haF1myfiCgidYAbfHJZymHGx
ytaNWQZdJAjAz25WUhqwEseKUS2y4mwAIhLUBq2LZKUqk/091jp17LJvcgwixnwcFlO35pw3atpW
Ge4MpjnbEixuh3M9ZqCN6A0IE0WkLOjmnlZyn4xywTBrua6IFd2gpIQDhK5Qo+i/cpdvhtfC2e23
KI89fJEq1HRqH1n0OZLWlA/fhPu0p1uqZf6gd8BUjmNwzXuBHeq7ox1u2u8lroF7oCdPJU3j03eq
v1lUS0oODY6mp8NsrTjU1os8WieXznH1qddWUyvSdnDHm8wcg2nYmyKr8zt4zHAwzcB8YPvq8xso
lf1LEk2NZ3opcF/QowTQC2ipdKkMtN8suPdp9iKjG/cVbDWvhbsYpESLdLghovbjml0Irxpsoq+d
AvYPfN3PIVMr7B6JZWJoSgkMmAar9W+3HYw4020mu8CF4EY5NEnsN1HssLuCnIT2s5uZyNnvSLnO
goUhBVAtoS4UXMfHuxyWE81il8XZ9XkPZA9sMWaP5KybL8j5cjJ5fP1yyMWfbLyo3RruP+HqFrUi
ts+Ff8ScyHL1KojyKKyRrBk6NFHD9ONAjJMDlFhItbAV6kS8IWICyipQUqOgHNjjzGewfrKgJ+K3
oqMkXG27TQ1TccIC2TxFKo8QhaoKuscDaNSVJFqSCQZ75UdKnQ2gqI4EJYE/aipqKQZAsIFiEcgG
Mgg+qjInvOslXaiIcztSYydThoeLaS0xW8iV1fJ78+PPav83CtJiZa4O8q6JWgarHlzdzYDNMa5x
vKQt8ITiiC4zflcpLSvGCf4f+Zpe6dwxsTMspxSPu8ZZ+1BuGQkNnnEDwHAjWIRIxVBBN5lg/AwY
A3m1C2+uc569Ze7NJEwtFRjCcteLSWs8FvxuhQ+11JsKMIpJvASYpxSjVI1tnhAyH5j397PmDSm7
vu/17LlrxAawhZvsGI0VsymuwQ5y624Hr4eLEwJVxG78lKASL9Ejm+rPpra9rccBRiVmkSWg7IqX
yQgZvjriJv+2K2WRRKdsamTV1gwgG+iiFCxJ01+O9HSltmQZZOa7Mb5ugAH//H81eNch0aEN+QGv
3kzi0TIKnL+9ro9rN9UpNpVMWDS2Z+BW3o8Pzy/z61vKyqclq8URDiedrKNMmwcAWkRMN/3pJa2P
mx3CZjDa0FQobwVRHpWsPaLWtR/2KrzQqcg1Bc8lOR7WIrNV/60rT+JFjnAZmfjPdTBdKAUVKE8m
rOrf5/f6bM3hTAJH84rCO0b81gBwazJqizlQZoB2Y4BzZuVbXtDPWsjnueiZ9BL7DGxgDI4eMugq
KIO7qwalmRhkaZV54zdfSDFeNopKWSagLMoRCF3VmliS5IZ8eTu2S0/hDdJe3zfxIlK6AIjCTl8D
0joLM2H76mKrdprfoodUWDLGzS4IIgvb+Oe39dKy6YikjDxRhCUiEgOzdcCzYuonmM6mchu6387Q
Aft8anAowl9Ki/MGAGZHUagM8cchfL0H5s06ZEFohY6hpfxOQLWjvhfkmBp9Qbo6oypsLP4K/eHO
4wgtYL5r0aJ8tYOm8uyKPhG7p9nLFLi1AXnJ2PrpHnXRGl2dmpXI3osEBvhiS60lHFMDiGF4On3U
ZeiMMYn6FD82/vIj3usOLWnhGGOF6o9w0aWLaDDACjCCM1TP9xRFDNgmZ7VMkRnWcqr5BH9g3xRU
6cu3NYTXwH2fBtdOtH9VmYgZtrHCWPcXmck1vHGXiVh4whAJdAZ6UgVMIvSOWXrtkmfIrZTYJDQb
gx27WDVyj7x36P2RsHPKGBMxLWouErhTcdo+BRlKKImy8RUg4dQHDcAHgr6XJUbTVfNZ4JuMSpb+
sKHuuyHXLqAPfBsk3uC9Jn2DYjvn2V5z8m2D3UpP1Q+bZ7USpWAGB58Jlc7qJhyzmjYfQhHh8ZZP
Cy04IgY718cT5d4Dyt4qxMcI0tE3Vwiwk/AqUVT+kQ2Yw2mVmeMb5NXUHDgpCdTFaXEA6h1EvaJb
7tkzlKMULapV9lsY65OOEEqgSfyGzEQ4J/AnGeZP8qIhzVsEw0r32BdXbDvj1ul0hcW8I5VRKbuQ
xD4RmShSi0HxupxLY1od8fIUq40IKUJdB4jnKxDUIcMFIGG3ibu4lJ+rITrtyAk6oHOhnAQaq1l6
C/F2AX9wpEJGqpkwnPhV3i/0kGqcXc+3c0rS+Cx9Jc6Vjk0ClBxPnMYBkevHy1+bZcio7XG+xine
TYwB/MotrwxHpRS++dzRBE4H3Zhsk+F/QpOBMllb9/r1k3c72m03MjTj8hDUs3IZuQmC56tQI5uK
lYlrSrJJRXKPvHeh9vndWNdAEZw7Pn6ldNXPsL52EGGg60VIEg+7ND5+dxibjeiOjjZI59+8bufG
CkRO7N2a0dFYiMbQqCDDgzSr6KLCI2QIIgjlgSSYAa+0zR5fzICUcuc9/o7hmvrOlJDqdKAT5Ldy
R2UpLa6+dO2n+eYDU3k61HGM+Xik2eYEAZ2xYgFT1XS994PtvCvkFayGDFuJGu/pjPUy5R9WgjP7
SX4tAEFxKm96jthVeI7lw4rtwOcLghquyxqGP8Vh2EAbojn3fPqJLy87mCM7ZTRXVOcSwvEW5CFD
MT2JkSxl3Q5y2vlv9e2/9ndLQuOimFG2xQTXdpNGqYCnsFjqSP1Ea5BqBkSw6YgAWflHw7XKpmcp
EuZWY3Eb7zGSOAn6vCGUUFSea4I3PChAPoBLciJ2LtUyt2Qf+BPDi8nkSt1SPkwB6lyixpp2Zy2f
Ke6tbI+UdP8wsZZxOVKoE+QBnhToAZ5xryWdkezveIUL408+ri5hmxdYpPbxTpLQBs8dV0GBCGBD
IUPmdnkspJi+l9VoIKeLuoINhv0D0UVW5oVTrU3ND3Ir/i6IkJlQQtkR8c5EPEwlHUhiWHaDlLPd
MtgK3ufML8ndR92XMtgYNvkoK52rDy7HvonmB90XLMM+bbBQa3ULqHhUM5qktod8X7iqaYBq/ZYk
rZuyEikWZB+i7BsZlMJwL0UhpMTvcIOXxli8KCG9zZzkfrUxznxdVAxYK2Nixv7WvqENJmj6TrSo
SRlivaq71Plar9yBgevpo+T5LtoOKpTI6j4vpvC4/OGEmPo8OKeafLnyiG1ps4WSYqiikSF2SFVV
7zwUZB4LJP2pj2BBJB7PAWLv0Isn6Nrep77Oy0JE+be0epdqDABwyg+MQGda+LwJwRXTb6lnGmRL
YL0iZlqBpX6u9tmJCpl6aITpoXufgdZodc8c3ghrVwJtNqpHAzq/gIyEp9VSmGo8dUx6QPvEl4dl
RVlCKWyPPdxgiGx92Ea3ubNMcgI1xnsYho7cCepd10j0FDDYyFz6K9TX00Ei1VdpxjsmHv+Ji9/I
gmGN/RmSv2VkOB94cufbqwmjNK7inKahjkUcA6OF9+bXupe383azNcYfhZMwOT2gM1eNnoqlPz7j
PWCAC0v/OdJWMUX3qqse2U0OALQaUXAjXh83eEzlUJWnevy2/usJOunnDwF8vLcXxHjC6brJl1ye
wzcqUYhLVaWc6wtQysnILauxFrs4mQFQjtFo324TUgGT5BfOeAfH6NPgKVGbO8tgIx1mnsfJz39E
2DTHYLQFPZlUZjC+xv3qKsgV6LEFdQTtGcZP+PvmjegA0gUEjFhrE3ymkxZy9ZKJsz6fnf1yW5kX
6eB2Ui0xMcSTSGAAEyPB0UTrsfA/GG2EulkilwOyFD0D9iUlgKHuGNiirOt5M4wHZK6d09S5GnZr
fVQQEpdhIWT3hYrOyP9ef6L9jQYdfVjnRBxCklk/7GY0TiBrBTLhLO01BTKaWMw5LqSCOIWhQ091
g/OojURXILa7YLqPY307SgN32ppa9hjpsaNSWNHUc5Oup7ez2oyULTbd+N3jc3aGT83ZFNo/83Co
Wutisx71CJOg8xORi6ysgiXT/jZQLyWw//YIZxHZL4XUGZIaj6JvqsnbNuFIqPspJa/ytMWTPek/
cKveRICLb5ceXORfuBT/ifz2DWKdH/3pgwybkYdCLkQmeuTtgQpZvOrStja49d7RNXFLCXLPobUI
wlZ9UtdmXC/e1UrGR61nf0Qehv1weiuq297QPbJtBK6zktnLr0msncKgv32l1LDP/wIuLJLK6Xa8
lGMRfq0CihbCWD03vGsBwrphTZZ1PS3bkrBDZ4m6kN2olMrDF/mLthm/lCyqOYlBDQbXUKMEUeCS
MOMUc+dfZt1s5+U92FnX6sMLna90lA3ezUUUmkdgfCK1xoHaaPAEL+iRmzD/k1zfr4Q0Gsuy8urZ
UCC883BKSSNHTd/23nQxeqD8Nww27ULqJgKDkQTWNCWmOipxLNG/WHlEs9EJZFLBdgSEdRr95oZo
5VCdBfRl8PnURniJHzL3Rz1kfPi7LDvgkN/zaukR2BRaprmMetczNFyEzhw/arhQcgpsf/H58rzQ
qGFrZsTsj+SF8VgoVmZL4xQgFPmgsnbPniNIURmNY77ZrRGlcsth+UERoMWChAk3B34mN/0+gJ9B
V0QTQOxgw7jcqKDJOQlM/4n6Fy/UgBgpUWnNzzpGMmWr+P92e6xtWSk61xBwcPsrZ3UPT9Y892S/
x00bXZu37Co2TjI1dG6n9A4U7RlhMfkHVPW46OrVH7d6giG2LNTk1jJAKNBtAV99e+Tk/wA6NvnW
dqtERPlFsIeeDW/TZVGEsHuabKJQH3oWQflgRcOY4RzB+BxeV6uDC6Pf+2KvwAaX5HbV/lbuZAk1
p2cagLylrN4TSoOnb34l05exPjPxvVY0smZDQWMOcwpu4EhDYf1jh6tGvOdUSGh/5ZVzQd5TDHk+
B8y7aaOTANCj2KXntWHAqH7xciqKutPQBKoCwClaabU2opRcgAZvku1OuTMSo13NJf8GDSJiXKGo
DVrF7ebCvsHBLk4K0R1wS0ybYB4p/R/JhjSVyKtx4rv/oYvKJZG5Y2T6vlyDoBAwfrdJQJxvWOb/
lZyHu4tR85dhIY1SgeGCUEdzOJSO4CbPG+WYYA9xcU02YqZT+h0F5+Ba73xr7/Bi+0G6oTFxejmA
ZvXx1hOXAwHO8+8KbgG1c5QJu76WRyc9/hMnQdTnOnn/P0OaChytO8TaLKAco5oVNvR2GFebwzTK
13qBLrzGHPsDF0O4jFqB0sAvxEX/2T9X86n2aUFRdGz1EoT4wMoDl1uwYveFWd5cjh7vNperxpNg
gFKduiAT5mwyQeUdiQWEd1m9Rp8qNhVyKvY8NWtyriu3S+xGIzeiD+OzmFJjPYDuKUWqEBo8euTy
Vx/E+93u0Mq0QBOMd9wlyjd/2+C1F9gc6vcWHXyYX1wk8GQrt4fFxFqa46b7JnIIuOlag2hiof9A
cNM32CPn7IPAJ8MwZMw/b43fRbwDSzJ6ufEL7RoPHK8dR02g8nx8iZmEq0UZPyKmoeCtFVXgO5+l
u3LdOwfJHKoV4EOCDXd6bsKMvCy62WdZxKhhllnhmyF+ugUqEvl5/CcUn98nWZNWPQqM7GdFC8K1
IXV4sP3G4a4Qos9nC4nD46VNXZnS//+aQJ3z3BDnaW0swLtwJXvVdi8Sguan1cndeFsY7pmvcy/x
QPFDFlH24KNjr8JnKg7JogoRfJeDO98utZezzO7oHFp9WkiGSTdYLBB7+nt3KwamJsC63pP6Udg4
+etgwS34RZLiC37/UKfwqyUo/D7jcG6yVHR66HwuBZKPogCOftc8xdaDXEqbQVSYA76MzNyaDwy9
XlM6PDuCc7LhDndQHwEFrbr4DU1lvpKuplS1FCGbpcpWpgtZ73SKGe1lwKNacmgXqN5rQ1Df8vuG
m0GPqPcMDYErsiNmjty0FRuUP+ggxmBTeNb1/lUmSpGGd9yLplCRppws57raIc86lxvnspFNrobA
cVnTIAeaekB4PZQtB02u8tUeOOaMJHzr1sIyNu8Pcj8n8+ezuWTd2BO7L2B/8eh8P1ArYAMa2y/7
2EwU4icm7HvEJoIWWJj9iOV7uUZLcwrozvFQDZ8m0N8h08l3z2eGxe6ltpwjuP/2d6Ky72A8IaUY
UPrx3O7YY89nZc+WVsmQGnl4bQsQ8fRN4ZexUq3s+HXOBSTmfBERMlwwvTK6LkLgz8JnuPEnAdYN
9KvtHzEXwb9sIuWNyqP7/yx4vZLU31FYfPQ4YOcDY2ajpZ4lhBYi9mFYcxzLUwQqGM9SNpGSVTx6
zqGJdtF2legb/gPRy51Yyu6nhru4wCK6d+Z97VKqe7zx8DW59iKNsr3uNArJUcPLVAJy7Cb5m2VQ
NzoH39eRQDl/fzgl/g76Y8Bo9Up2Bh3kOxFWXpvttQp5PLrvQ1aGPKomb2ovdKgFO3F0Z7wu5uBh
KVKeunrIQLlw/mvr5Tef/n4ZsFo6dpxSo8u+JkARmHcNkvcKwBfMB8k+m0bANs6aXg9/+MDfobii
boM84MdMBBmZwwYQ+heUEmv/sXSpcbNaFFOcRm/wt9wIl1E8GZ0N4Vr272OKYI1yQc6C0fhoY8PE
JBEIpU9zrIjRBBiD4d+3b1mkXzjq/0GJFWwn+yJgaRNVWn/WXX/2Abn1L2Q5savpBzZ9Rs4zU5dh
9Q9K8ASdl+ejqtGaeTHYLL9AiZboxbBBnXeqQpGbGcCzxLbHSIhTf6J/NVQLHBoftkVZMEBMB7nu
GUEr5onNkMHftcmdoaiuA/XnzMu60NVIpD7denbYpbwyF+kVlfsDToCMF+1VHfOaP7JRCyuWZDRG
CpYdqMgnnF86zbgwi6zioirLo7JaCHLye2xeThlkyEEJZ0V79R8y2C2lvz0/PM942QbUNeTtNsJ0
JEQ0FEiXaC7alUlzAk/luJMMPRAkITo9N4bBGNBCwh90AG87WBFqcHHfv20s8w9LIW1pHyXMj1Oo
IrO8qnGrz8q5Zon9Ib2m64yr92YZDWCysl3T16a2G1RefBrfvhH0EK64RRCLDzx8LbNzJ4XalBnU
j1vYI1tB5NuU7HzvNsjcnK1maC0T7jemZSqXbgtaVrnKtncvoL0KhmgAkdRpWjkdmdPPYs24Itt5
R2LgmbINM2WrRmtt7Ye74dWJN0LCzPDukMAt+rq6/odekQnrepusHLcSl7nqTP4cphEgbJBBWiK7
8qNgpNHh7Wtm+i+C885tcV9sS/3iu6cn8QIeapX5v3A4XKNNF2E/T5kALzL8dHJwQNNNPOebA6Qg
/GaEXzZ4ePohCjsJaU08bC9ZWdajt5XGJ6l6eb+5XupUBxEJYdU7KH7hI6+tF+e6nZe7wbDAbDcw
m1YphqY/nIeyuaUZGqueRGIr3XzuEwnUAHlOZoq3ZhYtcFY4Y3JGATZcAZpfKXSYLr1IqhH/KiNT
DjgEWN43tIfj0pX+sYZaDAw1Pqg60WNlOUdCH3rnmpz9PvKyjXzG47a1txE9vod/ZBZoVj6VNkxZ
fn79qnyKTQFrUxPZGRssc3iRxnGkLV+QiX5AFijffEA9CJARaqOazsV4i5KB93bJ9TiSH75wc1eM
uwrMNYS5ikFlXMDLvhhjwqLJNAZy10Pt0Z+5SNJ2CB6F5sryRTYl325gIJOxkBcWUcGnFDAOODiz
u8mWkL2diifpwfW5A831y7mDeWNPWZaI15girXkmRe7wCIOhdXOuet8oPRA8gVCBpQ+b9R6fkRpF
T1p8aHieqZtebCXjZFF+ZxzAbCHyjQiFv1hkN701n41Y9cpDXnU62gIsVdiiy+33uq994AfG94k0
VfMKCxzbBWDLRZEMyYPw0MSH2fMd15sDPfy72v5uYEF+iDiXNDZphpmKhoaSLQdcBdM9CrsAiVnk
akCwFHDjZhaJ4qJf3Ug0pRTBklTBU3tl4iC73pQgFZ3XlQ1kaoLtfq3ikoUYzgN9an8rS9fmoj4d
3a+/VvOn9kqA639Rrv10g0wgoBu3bdQcT6KU/Wy8jO2BoVD2JFOqw3PISTGCvKw0HRAXC0ObL07S
Wi+6Rn9/30lnauwKut2i/0JdllbhDwrc5826eEKS8DXJu0cWJcBOQ4IfavLm3LAPB8HCioMcIw8d
2p9Q4ph83xjMXJohasOCpagtOpK04W2xzUeY8XyyQZPeZ6skP03q3Dwqxj7yxj7FWSCI2lJO3eS+
135A8DdC1w54C7hSRkYzkXbe1imO3LrSD9xWHdXA+iNvp+3yUOgP24HxrvIlGPs2hMdQbfpSN/ge
r4uZyh8JG9vnApMl5ihen63SJESpssfbx9A+dN+pDVQFGXPhe1qu1QZ3g+Z7agyDBWWjGcpuQ42y
h4UMeTkz/ozFfjUWx91EWdDNz+lh+7uCQkD6cCVuVursabjYXO/5WbBvnXauCtR9P8pAxiQWH6vQ
jQD8my9xZCdDxmD4r8ZznDPTNBbNx67ZCQyLTI4iGH+mh9Hx9DuWSeQwcMc+FuKZj7sDYAhHdSAv
hzCqChMoOX3c893A98DG+bEmCFixogMuGnd3dnCbFbCvM2kwy07ip5U9Ekdkkm//tVhr6f0rJ6Av
dmsNacnXVLcunF3uTIaCRB79Fd5lbs/qkSq1qVmxySGKOZvlLJ7FlOTP9p7kcj6VMt9EoPZ5vRhR
QQASDP8vC7FOefBVs46rgJ/qxXC2QrNTZ10YqqzhBj8d4hQKF6phhduRJ5yvwEsgAoX7Oct812Ce
COGYDXKam6hMU4dQybznD3YAcK3+LQE65dBh3CMwjlk+e9RNAuaVFR2BNS7D6YCChi2SO18r2Xoc
8+UXLkOGF46NOcVFXywDYeyrI89NxlONUn7ldvf/Gduk0w2GatfZcWkkO/jBaaGpt5BsdoB+xub8
5rVWIYfGrDLT4FpZiIDWIVrfYgfwVoshzcKr4jtGFhxeVQoe9JZT5pTSewhTGu9LUfsJ/swPBZOh
MDovTmvSylpPC/rV3bZv1I+yYL8HwcNMZx7qMNy4AMLU+AdLWMZZn9Qsx8nJqGga9Zyq+bRb6DtE
HDenH5oI+oKO5ClpvVybR3O4gWj3j3FkFsKigtanKfr48OmsGfIXHJuCkYIrsfdbvslfaxrA+tmI
GvSom1yMFFljoou1xpqZ53ROg0Nc3LcF9FXkXbV4DE9MGWL4KY3sKgFB967ydWWa486n+h9tFJdz
LokBVaNWUNWdFIZQKyb4gKwKdn7xVXCh/QAu6+rbyZVxX0w8k4iQVJuliw16eFEgLdXOiclGdgzD
aK3hWcSNMpzqAyJels7u6R7VzpwtpW+BonLct7yc+Rzx5wSY+EHlT/+h1uXLPFS3kUzUYJi5gT9I
oa2YyRaTKWcap3EldpVXYVO2eHYjsxGGXI1VYM4Lc0XpLFy2hminqfDelNTKA3j104BpYYVRSUmC
ARK9CcR0KTQOIRjmIgUsydNPBL9UyxCxWaLyH4yhsiGD7CXGOEUTpvAZoaj01uZSMGGK2rNQ+6TZ
bQ3SwRyqeU6o1MK4T9q62Hr9qTDek7E7Qg/01hgKIqWj6F2FNwrFoaz8pxQVrYGsZImsJZQKQcy6
BnL5erK/UmABEsV34uYbuZJMdAskrLhkqIwRznWdz2DLV4BtTO72PEKvYYNyEEgHDZnlQNFKYmTx
5d0Ck4dauh5jvbHZgBGFMZjCTsdT8fUbEBJRcFYKmvAJ63zt2l97qGOGaEYwsHNlJZFXdG7iRaqc
UM5Awog01U+SrlXCHp7w5r9rdlzgt1P0gnW8SX6Or4ThC+8Ma0XFnxDfxdW9UcaOlabGZLVtkf4U
QzCcY02B2PGOgncxinR9OdDfijULKmlZliUi08zvxl5lAhTwWOSEyPQrUHBgeFVtQ1hfrgdrsMjt
u3Npls1miyj218j1jAchn5il4rxf6WWrj1ys+iGlCLq76LKYzFvtkq5Val9+T/axCFTyE65uekVq
4m/yG2FAwA0Sjf9xn0PF5Zg+v3a2B38gIwTpN+TD129w8nhEE39Yc+AqwkxLovK15ORVq/QGXkq7
zQl8nbZG4xiWbWdGcPrwgps6+AE2HnkS6KK4BRrYSJR2PuyNHMmldvLiy1Lsy+oaC3uYPfPEA/Qw
X1ELpJ74GshEDAPmEWYWD2neYf1g5uLAY2WGPLOZpthQr0ysgvLbUhVFPikrlni0kWyTMQxuVL3d
fUvUtQguHaNcm2XHNhj5mQN67lvv8VnIR2PdFqpDHbCncPD2AGmpQmXrGiVcj9IMfwqHF13vfkw8
GRd/AKRasRh9mKJES92/L2axvtLFiooMOYRARFB8CsicljUIPuCJnoo2Xm3muaLiGmsmtUozp0qQ
4xz6VP0tdHodz62ZFQtiiiHYHCuxmlxyWQc5irEPqI8i1EzkRadoAZJc+VR16RvweFQpnWQlH3CY
vu3SyXBI8uVTaF8XuVYpZ856zph1r/nf0a7tOZrG3bDBupuFI6+6NB1Hv8o1I2MRSfncG63idxXu
7BXd96N6I/oIu7cJXqwy3kff3KRa3r3rXiKnkhhvvDwjiySNQGNFrDJOFdnvVh7a2CE+wY6g1jMs
4UIsMYltiZGzO5fKE9V5jewMw8tDs+aEa2RZHND6Wn+EkcurtirWTgRQIHqu59sFNxHW4dhAAtLt
iGPRXlSX++O6615bj+mZtOdKRatV32IbC2uO5XrUeiiQyigE8O0GbnJguBEV0K/w8jaixSNjLp6p
SwvcusYWMbERaM8XmeWSCH3HqrjaHmXZI+JMpzg2bfEluVZGs2mpaL+vwD/WiB+h/UYiYrT0pp4D
9cyqf42b2445QVm2t6/0++SfDvGA6WAWCvxw9QL2iwwpU1Ea7IrmCeEI9K1X8Nky65pwH2l15CWp
FG/2HyafaZtVlTlZRFsOElykGz+kSlGPPS7YlYhxlEIjDEgQ3UbQRqsIRWKWsch5Yf30Aq41o7zC
t2vx1NEXns/wH29AghQRGQPSmfev8MkQiZrGRfHEi4Jd6ITB1LzSYV/wvmL38J4uY5CJYftnvbIc
cxtoPVtx0iE66AcLNz9Chj+kgDmbxRPWXgWqMKrvRxv0Lh0Ob016BMIJRXETZTcPzz8DkjK02kI1
Is5Gc4Ge6CrY31rm/H0qrJhyybaff0CnALPEuez0jm5JjxizkHvYocSyz7BRBGIiQEKChw3SaUWv
epuqGOtutC640NDTnVDvbX19NXL45xkjY+HyehG27Jdfh9MCqqwJDlu4VKIwOacGLSbVicuzznzK
HnsO7lN4Lg/2JzHzj2TMeeqS5B4Xp4ss5RWZDaJYBv5GWExU+reFj2q+GqX62zLsXZbdEC0HyJRv
b9jjIYrdChE+ilWkWiJfIZE27Rey8FVHRfFmqGI/HzB8bSQThLj5bJ6w0vUk+D7jLi4c36QdmySZ
pppVEjTzpski5Jz8yDLjQO1/InzlnOelQJROhBnxbtjEY1hpypS+UewmTUVb/g4QuuAcpd+gxlH4
aHpUHmwRwWNV2GbywXXrBiB+K57NZve0d3XPmOzkAwU997iFEA6v3qcxSYA657cCpEd2Flpsdozt
hvTWgSpFT11Sgd9QNCAykd6tK+BdQTPu6x8WYsZEzpATIw9Trir0Dn047drXdeuKY3zu4gHwS8rN
E0K4OaTug6ABjxFs1icR50lItaHulScOuHZw4ypRyVw4jjUHwnGoXn+lYF2x+KpAKqSU84Ocljln
7PQZZ8fysha2yUrEEEWTqmCmcZPaR4OAGdIIUPZDuMLe5Nj6gkUHO/r0Mx+JcUs3zelmlfObS3ib
HOiyC/XohmAlRXuXJhmGoMDBGLdshJI7LehZJzdgHtS3S+unoQXwSPZmpbUV9Bnob0bXEq8J28ur
YRIiR43snG8CUeQ14P6BrrS5VDow/NX6iSRrA3gZJMCMx4Cbnllnr0JcdaU6ig8RfDzq7/prtbFE
GgTs8kWf89Z6O3+fPDh0damgtFgIqAhM6nOopJPP/ZS64zmYYwH4stQ5SSM3iyM5EcG8X+GOvDgW
p2Egy9uKSWom45cMqsr3d2aDynHU9R4BIkNqVLvI+Iy41bsCG9MObJ6E3hZ9wzAZkD0nBLG9hE5a
OegY1zAzoqUWvMnvuGQKZYybZ/ddfAjXufTsACuwlDezDbWtggzeLcCoGaMcQO9etCYFp2m4wMb/
Wgxv2UE5opvr1kYKl1pGPOoWkIvraIPBNfjG4zgK7Kctm/55Grr3UhYp3bNkJxotkQ5uGp8+xtN0
uRumtBdH9MA9G69QNf69dyAKxiH0xpP/Nu4CCBsj8BTBJJgVoS1BDIAmsX7ACGysUJp756nj+mc3
K0rxGkKoMAZ31BKYYv5s2xKUm7tKRI5fbYheWeSVlNMkYiNO8d8aPUBZ9N/gcZyvb4dFfHspQwey
HJSclh/baZwk8wahLp/MuWTN76/ZgNzGCzaRVtyuBviOdSSVosZR21lOIDOf02d964SRSuwBp+Fz
QZoSJiX7sKDAIjnd9TVThRz8zIdMMYF49R7zfkMkmeBtcgJ+867MMCsy8Wk+AF+iqd5P7+dd2Qdw
1EX9RX5yJkY3XL1Bvq8TaVymOEeWRaNokNZn4E05nF7U+wXsTATrprBNiypiu2IyecYAu7Arzn8+
3Tr4go444Cj7EI0vnTLFpDc1KWXrxcCG3qr6lDkLfecieVZV7jJzD23V2gG3dtCimcp8Mk95GoED
YR99rgJOjaShBGga/tJSwnJ4k7B2j/8kRtS3jVrNyEcHojVC6ZM0jA+laUp5oi36ZS8CtzhMYxpa
ZYdaRBI2kIUNMzyttPkx8b7TAfv/x03w0LQzkoaO5YmaH26GVbJbf2MIYmmzVjusRI0AUlmRzt4W
V40qDD2Bpf7Z5P15wT1WrHwSvZS2q51rPQBo1YQqHe9o56/YxILrwwcilWxh/kvzOIOzkfmvTPsc
NkyD423QyJ7IHkUmFylBXo8KHhuIxDLGJKcVFIRMNwlkQCFHvabfNL3C3IacN7j6N5snlYcryBkn
NNOQFhZIkZnjj+/wWmqdDF9PHKdQ25uFg8GVe3qggWebndI7RK86JeUqPuPqb/lt0R2vGBD3XMky
CH8Si1LXz+NIVELCmZZJZFRgRVJLFx6eRHmgPAJE4i45Mndc369vw/WrM16ZYtoNmaQh0BIV1ZjQ
Knp5kKA3hV93p/OPzTQuRdkg1KiL7/8wQ11pIayXcpMJmY5ZoAihn0GqIPzT/30znUT5xFNYSG6u
1HHcjmdP1QYbeg/iPlXY5B6DBUmkA6scLZFs8Qvzc6pbWLT8RPj8IquX137+A1CQCQjYkLYviwgE
JzzLR7u/4+v0v4Zs7BC47jLU4n4NPGS+wAt5Mu7IgsfM5M04Nkbkrpg0zZF5Vqs9KOHKNlV2mlWC
0fJFLbvgbQBH6VHlJnOkUz4ri1+lAsT4T/SUVVDouhXaUEDF7TGFgnaPv96jhxjBW/SOobfzmq1T
hEDcz1tSK5ybWVqXktacUOKc04ArxXT8GxaassJFtSAvO8Sj/6z1FZibrIKn2l0tvXYr4KG5dxfR
JVXQLyFed6esviyT3mghc93ndT+sOVLwrUc6y84Eh9l1LFx/aC8a4nUx9BILma6LV2KltdEFhgxg
WHy2x3jKFlCOnXp3ZEh1Z3T70F8V/JEOKNqyugBZYIESJWN94o+OwV4A2FbMzg43XZkHxWvYLhGY
joo8U1LASMQzq7S/Hef/57ByYRng+yA/K3QiRkVT1y680JBFcPBPhK90MbShVyof+VQM8oXjW/KA
KIwEoyI9BG1tSuS8XlJBmDvOqIZpJXn0IAnov4M8Wf+/lkLtHOMePR3W2QEbWhPZPQOOUdjPHChu
/2dzAR+nJAGZJIpXNVYE/oL2tUbco60SGTV2HwBR81VUy3QUyuNK9bDbW4XPEwlICGhgn/dO14yl
SRJM/KAaHwSPpoKt7kyHwYuJdHi4zOqDle21t/zZigbDa4BbNXDCNFwAB9sOgxap+QZG6Dw1wP92
kmyDoviYZ0Hpjh4fmLHkgcemensqqfiAjTiKhj6HimxDviLelLt+4TiSLhbA1805PrXK4cZzopf3
suGRS3T2yDuDKwJB9tmG93/CgkeQ19D7etnoKeGR4WCgA+Jh/o8wPpD6YUipzgmiGgPhiZQXv5qo
gEx3l1I8Fse91suslP6Mu4MlLHxxruSwhufw/4KeJq0+tGypB3ZfkeiBOaPOKQjHIC5UHW0u3IGm
7O5eCR2kVdrXY7iSm/VxYNgGcYB9MBFZ224eDszD0hRjQ4oLO7D1SYNnAcUGnN3TutS2ybM/MYFN
f1KNVSAhbTqN0oatbbK4HZOEhi9W6S0mdb545uHS9EapTSrM4cmABAbJ9btu4kv1qf+hUQkefJKY
sqXpLXN1CVt4Dy84WIdRECRmRlQyPU1ECNkrslxhR6iaEJEwCbVVQXKbY0BrCZX9L4mNWql6skLQ
J3rRMkht0Z6aQ94wXpRuPi2R9wR1zyzyJAWi22LyjhLCmzGCKXxzuYXyREi6UnnyB7RaELXIuS4k
ykIIaDPVe3mO0OllhEEQceZ3MK++ynpNp9JM36rw7G0zW0ybeaWGT6WsL7wcTXzH9zfW42dDcH0+
JM/BJL+sRwQ/w2w8O2oNMfOwu22yZXn70wwVHyi5kOFiVkcYPJQUTt/jvOv8EBTMGwJriyoLfFv1
GlryVhdpF0IJnEI1UV9DqCQTKo4ABE/TBP9hD4Yu6Ge1XxZNn74trRYFy5WXQL9/nabvfQNBXE8V
iCuPAxW3hDKg43MyfB+qOZ+7ZhGtofGs62iHt3EC/gTXr0IXnr8EHkgo0wOMakQXCII1ckJVbDY3
lwGWHJzhjZavnmx5tPnPSnujAS734Cw2jwON9A9LM4icsT7GsscopfO/adi/IoFg/Rdm8cXm38UU
yU2lmMjiQDhqGg49VLhX/PBY0bFSESPQHuMazPrL2ay/mbUdGaK+BeDlJ2nF+cPyVq57oreIXs8M
mG+NtbDRFYlkGgEQdgYb8v7fConf52hvsaZW2CkSS0Ep/XTm7RlhoNKilGys0hxvw9Ccxu+5vzKQ
7nGn0/v1WeybuI7ickypNUugBx+L1177iCrdh0dg+CAAjiZ92fb7F3cd/HTArBzbVbMRTFv2NHCE
6nwk+RavxCJ0Y4phVGeC63wNT3Q8fV8V2nXUrGlDImNP+U2H78vuDQsAFX/5b0fv8i2nq2D4Ac7A
L1HzvWBbsok/R9c0bHGjPgMGwJ0f5YrjAODa1kTd8g9FOYDyLkKUNcL+VX/kmrTv9Z9gxvYzZBLq
oXFrp0KIKZz2tNZ0WdR7kJB8QsPbjLOiZ1A/NJVNBlA+GNrBAdW2bzLG5rtExDUFxZkrQFG5y893
goA6w7WB68zj5yDK4u5tSJrp9mH0gIgCGUGwEuuHbpPm0bNJ20JOmGO6LohpapSeaxxbbk3tNaVO
nUEnJjkn4sgUQ/uwrZrFlQ+xr9C0MYi76SFs5soqD2wPJ83V6WMLZz3IYL18C+hvyeqznPWttFwF
AdWW5IvBAtnX38vLtsvm1zY1i9xbcx4ho8cR0vbBAaCMv1argO3DWzYd1APZOnslECLfVL2Hr5IL
BiLosf3hpGlxrMlWhSv3rJT7pX46MWT/x8bQdZ+3QkQ39jIdgMWAkeEsJT7i+1wIwVCeVIMvRuhO
jFFhPrJZTturbwbXWZ2xg7k9po7scRsuRb8yS0BTHALOKdY/9aoirRrrt7NYhH6yJKDn1PPVBeTc
k57Zy+iMFXsASmuXo2GZ0KxMOSiWYQrr1UyGNhrbwu8pw96qY8duQMWY+1N1yCU6O9yLXEdjxDuT
w4TEmQ9Hszs2bavCSM3WXcHbGHJdF2NQ3qJzyLFISOMcIdVUbWCt3MpVQcXTEavLhg9mYoQelNJJ
RZ7jMf3fYmgBleG9XdWpbOuoC6/jCtiZGWqRE548vUbSdo80eMPtQhsYC99PV8E7hvortQ4DEXfI
VYmTH1SYqosRJRTOCfIIt/Q6gEIbcrdCgjgMfgzgTRIhobJ/mIQMqeAyfis+aMqIZ/7nsahdMVDw
smfTTxld4146zQbm27dtcyM6x1xc9DX9stHmpSqzyduuL6A/gid0awlUeWPUtGTScqIJaoOQqnJR
7X8VIpA5xAmuorMiemvW6Tqv/a/WEthjMLqGTUaZTOoi5O8mWnQB0iLFzscYYFjqNU5IEbXvQPOY
eHS8UijIUv3vcz2A5RiSMX4Af4L6UPG/EpdoO5EcyCprJMl/M4MTvOJofhrD1vq00HpN+QA+7yNb
qLVSl78J7U/9gfnp3TxaGxIEcyUahSAIWXD9SzRl9j/f7fdAw3Vp2E9bTJ0ZRs+wHkzYTyGKNDs3
4mu+1sSW6Hu+2oFsgaUHVPpWbSmtTyIIkkwUlToc9ZPx5830EunfUfq61NAZU1DPXgtdbRIr1G5u
SseLxqKasMsnh03VV5ymIYexUY9CRN9+UK9FieYgCwS9PBDBLMPgyS+vDqIXrzwI9bqdtAwYD4d2
AsBl3MVgn3xySmLMqL2jsV9z0g6PyPwNIn0U0hrVAdzTvFssJFZRx/CL3r+90B/HSr1sLmlsHrw8
h2JufHMs5DWXGgLmv1qfM+dZp06aAbaDP7AUWwyn8bVka9s5GBoeGX4ENGTiYQf0DGxFq/bTUfF/
hGHb9w+24wRoHzkE6o2wFyA/OS6H1tpALTOQd3U0uOmf2AX6+XrXQ+HzRXFzVeS5Yh0buOXIZBOW
xmN6zbpLfStDS+XL53MRXAE5NqwYKlGFGHyE/8cK3IfVRXWhMu3ncUGDiINCctOSm8KljnaL8xmd
CgyT7PvYsuJyTnmrarJCdCHz82ZlNmMEm9v42QGCQySH7gDReF1U794JUqJMnjm4LjPwlq5Jv7n7
zdAQLUzaPE/8dm0IPKqpwVb1d3sTjvXoj4ZRyiJQ+kxds/SDE2Sa49LwIVbr+ssU5bolOR9zxeYn
LXmIHOYgSZN18Oh/5HvTnG8PAqgxutE6ByRzkf3WFaBaB2S9djZNQ/nnoh4xa/KV3N3PiBZnUg0A
0HdxZoCNL3ZJ0sf6L+mSlleaaPmprMzByizqqt8JHb3VVQGH+DHrApAdrLzApooqmbBGR5erJYLR
GmDIbOid8xR0B9Wsxs/YqcupjmZEzfQeQaNRpJ6mLblSyraphmC8iCFaTnr1XAoMxxH2tE5wK7UH
BsugovvydMDp/zfNfZCA6oGU+TncuEpjN4RMF+/NK4LF+GQjEJjPCgRra69VIwC5X6Y4U+Byw/zz
KqS53yvdzRT8TZvGb1G/myB7eiWy34QouE0A2OEdz7XBFwFVkK6e7zbspp+aLnAzjnvkD8GfzzGu
pUvEh2bSYEbpd8F/0c0eUsnbJC6syJlwpAKeCj9+G4ZtfYx4mTyHjJbPNnqKa471c1qx9bfTWCwt
sxzEvSNeVupHg9LpJQ1RpjjpXMGBPbtL5hprICtQWPnWNDgJoBEoMTfXmBf8+7og7mvXcqBO3Z1R
tea9hKDkm8lx4qW3481cWQr1+C7ifTj4iyNiOIuOoQaRHaesBhu0sAvPeUOf8LdsUgkxC2OesogO
v5Ws5KF6YudcqrVGkeCVwHVnRVW1g/OSWjCYDIFnfmUm9HcT4r1MfFJuaXuX22BL7WXe1isYoTxZ
K5SvcWusSeQu7ngz9wwEuTtK5Ri0y8zVJe1PoJEYCiEwwOtuNMjb2NH7dTupjgdwCcxXfnaTaTGb
QnO+lfB04v4TfxQRF4clfQh4KxX8Per4fmmdIaUPfefg2SZNSD1TelF3WYnm+ynZD7gN/6/Ubdyx
J25iRPXwJpp4g4uGJ1hHHHq76irODu+Fap0LYG91RKhitLjZWoYqoj3Hv/DRnRuCBTafsDtMJsqu
JSiSmRH+GocMYO4/fVh7Qiq5TbwLdqD5274h5AXqlcuD5CvWDefMtwcQ7JLTH8eS9xVqYfO8ErJd
AS+TtGH8OJ/IiC+ClAurgVa4d8Thpx/zBq2QbbAu2hMXmKFnt9G6nyCFEzS3yvMXO/IzMPs93f7K
j14hQQBb+HHjPJsPCU09HJVwbOtd2PT2bwfZmceTW6HPoy/QtHEqZVP8XVaTarbh/ATnNhIwhYd1
hEHlgdqyjDf5cZsH+OwsO9M/DfEdRlND6jbh+AhCJl+BU3ilXD4LCREdDXim19ZgXKlEWSLGNtYv
XH54OhyEsumCIXgCTENlwejCP9lcqUZrsAXst5n6usP9vzvqDMQH0LMp2JmnMjSnAyTMWk/NqD5+
ys3F5JNX21LH22qu8ht9AoUfiq8bNhZB9+PUy9z7Pm7FIMYmMuormXx67EhD2YEs8TL0ivKDonul
YqehND+cCmC5AiyCEX3oxeQv+I+mbJcoinoszx+mNo2N253sn0uudVP4X7oRhvhvkz46pv4VaR55
7uryZkoaz4AyFEN1GVjDre1q7w/+5pXN1UurhKhsoBb98gq3oXzVE25R/6TZCjGk9etBL20rjrav
d4nCmeVkAqJykCywe7d960xc1AXWhghiqKj11QBzvslR3R7WS3RbbU0wiC6dIzwEUTCk3bylLDkp
p5eyOwKMeh4WyJ+kyc6dK9xSC4BcuH6UIXRGRrE7BDSIjxg+C+MCyK65Rhgn1l0XoL9jxbuKJ7EM
P/QfEwT7VmnKF+kL1ZixlgciyiRmKmO5iq4VgHUIV8tLl+mIgFfyiP2GMrBdH8EHn7bL4AmOE+X/
FxrlweOwHcrAOLRo93jGivdy8NY0HjpCp+ss7qry9yurxWukKHFFeJ0wrxSs1wc+83/ODk/AumOA
jPIw797/Bew4ZF65wYHlpIcPN779Yn551t8IfvAx7LwiIYJhIy3KmQMd/Umlw5pUpqCSPkFjTFm6
JYlHQgV6svi8d/3PjB/GcOJN2AhvZ4N0Zqz0x2HGTrq5TWijw2kibUzUTTNfP3zaHuTItAmAJOZO
ZdFMHj5Mza/+pZ8Y6Drs2ENCxGEVVpC669Qhcmg/XCYoPu1RhnyMPKq2Kd5nkVMVRNjNTG0IjOlA
Cy3LtRTc/4udcW5P+d/5eg+9ZImaK+hQ8Ki4jMiYBwE/YAiFp4wmdCo+VcMvUT1Nr6119jlLVzGh
jSl6hFsWnalbM3SZRrFjblKYUHYoGRnPmxUYtymMUeLCnwwBx7TgKa1TngTaDWeODkskFSF2IsqS
xMuFs01TXCWidd6YsPCcviIKlqL0/Ahjnn+BONz82KmNEKxZEEvLKRzf6MrKx2dbQ9XqxAlMh2yy
VIzEH+AUwBdzGC5d0JPnKCwiVMdMBwEWEOqEC+CwHbFPV4yQ1jFNzrATM8oLyWk+loAlrsqvo8Vm
okTRYyT0hLZpUP9VVmwrWH6Mi0IgGWHz7Onktp0TFnKDSID7DLlj8aQ5MO3hlmI9mq6jFu/f1tZY
WGoRLTLpsOIBwPX+f8yHNpADy7r3Kouq+4bno0crRRuLjkiRTkXgZJiLS7OquODGrZJNr6knzXPR
KiujPO5mEKUgMAHDC/UHnlWnHd+W4v7Y5JZvsxdQiz0TXeEq7O1zDByT4KjDmF3L/x6zYSRJsjjm
OS3VYORKKGB2k2pWZGjiAAfKXukqLAGQNRc5osGz2fLoiFveeLoplPcQ20MO/5knv9h3ncOxx67z
h1nQvlq/RrhszNu/ZZ0CLmqTVaZZ2AsfEr0xmnxxkGO/ysGehUb7VyinnE180zypnvxDNUyKu2Td
9eN+sJjSp0us+A2X4QBk/x/e7PswnQlAT8K+ueXu+VSTAi+F/v05dBMk+KQ4m0UK19a1lHfkS8mZ
rZwdFR1Rr3gyy5JHZZ1jLzfCzPK7ZgL3cxQb0eq9QhCvTZZnyxsUxKB4pi4ISFA/S0DseNxT+wYd
0oTp4QVSsYj2j5bfQL7Bgjlk6fTBVFFYTjxYw3iqkI0mafw7wEr11tnKFtAqTnxSzc+m/5ByOPKX
Bn08itxJkN58jHtIgI6aFcRHfyED79L9O7CFSJjrZj7jKYXCCJ+4F8p7oAmysYVfSu422yKpBRQm
Y0+4BjJQPLtoOteZoITCu+jR5yu0CmNvirtP4GMgIk4w+ivp6yMiG+ds0WHbtlm4/LKV7mwJvDh5
4Q267blu+ABySP8Uh8MrXNhZx3dZ+0CeIQ5OY1WheRCW3OG0A1wHuFwarg7TGH5U/lmCu3LfeME7
dYRdYWf6N4akOKzB5aUDnAZPyV62eYXfAvQCUQNoR8Va5gefoD/Yfpc/6bNazz9iZUApbyhUnMSS
yq3wY7qH9TdYZ3ppDjSvEoWi5BQ993DcGL5cSHtdOR699VAPogS23QS1zcJpyxVO44v+C68p0lQS
kkM6BgtKTyagKzrJov0gr513vOrQQ5psGYbBR1YUZsnoFsbzqLe6uD7kOket6s1dh2CSOzRb3/IG
ZPTuGV+C8Nd9Q6eGPVAG4gHQx+0p7BgxOuujrFAk7/RwQlI2J1mpTVsS7oH46icj+0VyZfhK27sA
nru7i5tvQVLmHF4WZnIGpqtChwiHLJTvbu2rknfn9T0wsi0m9v1cDvcxx4mthCc+nyYsw4S023Uv
K4hvdnn/dWPwvM7W2mZpB5s2OsVdOc6MqQJgFldNaYhxfD8GxDt1KlpDD5qOMA3dE0nhvyjtT9g1
yp+fA9tc/yJ5vw/O/9uxFPfQ83C5J0kL4VOaJLIa1N0c9ci6hpsjzkGjNDv8zRwXKbNNDgV6q11m
lfuexBwh8oyp6fB0hmBcdDjHtL4Dg66ny5jDnfYImAJuWU8bvJaRxJCvIFAsKK9Z7cufT28N2lrS
CPxSeckMtDbIA/jsj18xishuB2TSy9OebkR8DMbMOVL3ZN9s10bN4sXGqCdq+FTZw6T2bc7DIcrr
PL1jKa5GSJnVHNvrTTRhFLDpoccmTYP9U18G6A/8kCnLUuFhb8OvxvGAnsmAkiT48YCIxW7Cgvax
9s16D4rXxxF3UVWcPa9Vnn35sGVWB9JfOdB+A4JkVw6IZP0dMMvdRXI+UJJyJDRk0sVpWg/Z0oLf
XbtQFKkZZwCVuCYQFpUEABP0wNXN5yXW2+D/ym5hiqVu1tZt+hBhXiTJ38+aM6VJ6fBs+EQ/bWcv
evfwCdx/4dttQA1vrN6SFFqOs9GMHzlpsVqo9RQjFC8oRDsmXSacYPEqkm7ZRC9zEVCg/odEwIJw
lRd+CVFET9P+T65X3PJFpuugNySakTTvm9tqpRyR6u3K/6IvkjC9e5dpbqj+UdlssnwoL83f7DdR
FNMbMyQ2U/11vij4MvYagJNID7uvGjMgf4Ndd5saLfwFbx07G7Tv4v6t1jgFL2zZFXKpViP3ArbM
00OZZEPzACgMb1kvbUJfGSgIYYhxwHvLUGpZLREf1z5Kj0u3N2xOWQo9V3i/HnIg56+bDRg/0Yad
cI7XaImJD+PwZYwzAdBi5vKCwA7NZF6dbJhvXgiSQ5ayGgesW9ezKTYgvTM6lDhgKgsLNGbkwtYl
YxjEzUscN0N6ZZPj29j46oVkGx0fYQbNsS0KZheH9aPSoz6rbXYAGhNgCRyj0nIbkz/Fh3H6gpvy
wyNYzU2IM2bpyt0qL38Yslfb1hFC4WI9qKIPxtuuhZ8DK3fhdo2QOylj5lyiR6oDo9a3vfITueMi
B9FZbom23sS8jsSqVswpUVAhXiesG+2ZSZXfq5eYex+FK9FnhV8E216XeWq45PW21D6Pijtc+PZW
NF6TM1/IlbsigSoEP/y6g2P6wKP43IF3UFMQi0oi1mhu6eL1Rk8+rL5KUs+I0XkQd2QIbotRx0at
sBwPaYBN0xXTb9RBY3tnLs6uyYf308Nc5O3qy0l8uoS/s8r9kV28xErhblGCTSdpZd+UDnGR2ADN
53C6NvmsEeUUVaI9E7ZNAz6kR64+RWaZohK+qAtEGaszWSTyc5ukDl07OnbLg+kbx6N45II+ZuLB
v9habGWQna+5ZHIV2VJFgAGfyOk0rCDuHH9Z+FFSeMrW/yrpUQ4PuJppsYT/kA/Xi3YFdEZ8iU0h
YWWCq7XhDqylrHAkVWhbpjogY73e7wulOKmEUmKJvKF+1aLekrQudYAo284NA/W4qY0EmpKtU5Kn
SYaFKkeE1BX1fVT6QIJqxmAnHyJbocvZHNbQ5+6mIAbPsEsPx63R712rZy+Y3ubnI0o8tZoJOPHZ
lbyyj9EwHxOeIle4i/fW+OTFLHcMoR71HWD7wfmnPRoP24aNsEISc6jwwhw/W0JZrp2C06cRwCiQ
d3swxYoEGKhHyQrxUINquYgIr9AipKUE29BtYNyT5T8ROuj9uj5NI5MQp4g9rgSmZmoPmtNIcqev
B4ZGGuuPzbkI+AlCKKej7ReS5iU2kO/gjkVO4719jJnxFKnJPajDUH5xfq7D/QykGnR93D/astnU
tlnlgwCXgjsS8bDKmgDj4I+NjawtuRfW6pJFfgB8VQ2oBJgyN4WG0KhS/Z9jKEha3+2cFejDmWB/
tsHFdzAkSu/eamkr8ghY1JlXagSCFG9ePjtKVKcuS5zGHZe2FmzHbcbQrhiAaAi675uffb+PhqhY
QeLM4bvhLdcwKCTVxfgw6yyTZuWaTYYNpVIoZyAuHbk4Rs5kpIO8B+QgAIXQsr1SC1mD8uQa55kT
m4KYGik1YLkBHyi52+RALSPTPmnpZXFfct+qXzH1yYTMiTTFb3QnEn7QrFikfzlChncpxgo8Vn+A
y0N4XRhroHIhYp/ZDWneorZKb4N0enlE3IU6cZB5/PVPftLg/Pqr/ZTYKggoG1l4IDQ1SObOwMe8
5z8F2TRZJ/EvFg0N2iudX6C2k6XocfqpAkNgapW5Ws8YMbcrokOYxYiufoGJCjmuOJHv9mri+Sz5
Vpy1bzWC6lW0JuSXqRQ+IAiKVUz4I8sBC9d0ROg46tQnLNefll6cjfWc/8eFCldZIQxTAblkwyWe
hVk3lnTxYfVkflrGflLe9g+IrAZsEi46Cn1FnaUGn63Ob7qgGWpWytcnZBbSBZtK4cW/KMWmnKoo
Rk0JWRG0VlxFV618MDQbJzfGIXeabUuImwcbgHf8LnDl85RvAOoucAUUWVq0YlZTKQCdaCULFLo9
f1MswJ3zxSzyQefx2lh6iz86IjuSDvzOGuXHWleLVPyBbCR/wYx8hhpaAUEXB6MPuBXvRXjOy2qc
yqrg6qER1UUt581IKuowcyocOq3mhV7X/MTcTq+ECPUKxupJLpcYfdIAwi1Sr8FfGlfbvFV73t1v
BpTgMZa9V8gxQyT/uA3vbXoxvfxSx2p82gPaRdFWqMLkBZ7aJaTqwNSImS73GWwUdHg9TivHKtWV
Z28Lx0vh4A5DWbiL0Ja8pLS2bCK+ZVxqfrHcD/1uZWA2XYH0n0lP4ZCc+wD8iwbqcMqj4Y0HRr7I
Jc1AiGakjOYfuy9T17TLo/lx3uWTQ+xeKIxesEB0eenPZzO5Dn/1K5c3FenfL1ehblUWPNcPNy9i
mmK3IAi0iFvC5MG17G3mRrM2iG8eYrhzHnFtUnSW6YPsl+xftUFgamF399qCPg6nIb4UjacLgsAZ
913Y6GFLV/xzZUInvcR+x9ElT0U1+7hzc/bvriBDVVg/VZU2RxR/5BPifeCMTae30BkeuVyND7tW
JAkXtDJPw4JUkEt/FVH36zFimUuTySgAIbEWpyki/J3ZCBH1F28jIPcZRifM355oML86w/Rv72d7
OAM3wYXCYr7B3B9PmmeEGJCiRm2UtD+PAKIXDXvdyPtzeV8b7gfPatsOqXhNEvbe/Z8jKh6A59zz
VWfpZ5ILJ0akjqzevJJMePFJz+cR3cBog9h/Qu4iLzdYXE1MIoDY1Jiz5yk5rwjfuGDzoy1ri54f
xQ4nJQQa8xsd3KzFqbtYKeJq4gt+hhRZ77ciG7y1OhMPxnAquPJvhB2jNZBEB27nNy07hiNKs7LD
/LcLabu/hpfCpLVYR5bMsT1qyHH48loj5Qwtrz8xW99eNNCKWds7NH86Ixb3LnZaHZZDY7rMASFb
RftUfpZsAApEKBbAL6Y+jfeNo6+uR16MYROEplHDB33mj0AHPeXuw3711PGd4bBWNvjrZRRGBiti
PSnrO5gQPcvYkPvHIPFcWt0d4eKP12PwS4o7pUedvPFEHxWPYPejovkSUAFyf7L40Ge6YgANd76K
QbNTCG14XVfenSO181YsW5UbS/GJSSTM6bTw+BzOrYOvA7UoAn1bQ86TFyADcXK8HAd5264yvQzS
NkyvuCcbAAJcPl1UTwlyU9zvvUkWhnE47bGPbrrfQmTVznpxHNytsozB9CZ0XhVTp5FLcesxHhJP
pVniLeLyCjgrGDjx0YfBVj3M8Jh7Nil/vWzvcjTdVdqoUL4IB3CkeEW1VqrdHsTS5bxIfpJcmOpS
OH7u2hSxlasBdGLDYmUF5JzumOSkbdw6gX2puQ9vi8fNBc/MtySyWcE/wjgZPGHpIoXNHnvEIUfp
cQt7nuRpmv16xPut7xEwBVddwjsTBOIj+MON7SVjzygc4J9eQvmiqxR7ZHpg81Z63znukPmAxNFE
YW7+atIy6JoOsZ6tLlpxmi73qq8WE2zPfIKplDQjSMTu2w20N12WBfsjf2Cz+J0QiKK6s/+sUgfc
0zqOulfIDr8EZ6My9gejvH8LC0O+oQz1fJSp+OvUQW8V+mJQtWJ8OitLLGfdOmqSKeU1uodNdVWz
miJ29KHHD99D8Imn/X3F1UB6ZbiYgLSgkAbJCS7xjQj/LDiwABwu9nf2l2c78JQGINl+RRLpT96H
LN+ObbFaeRSMDIG1el4KmO963Unek4xKHc9d0rhr4Ul0AloNJXK7v2kl1pmssUlREtwAVjehovt0
9N9lkbyJ8XhWDxqM0HFf+Kg3LknCHJsmPUTMfsipPxm8wslOfdYn6xSrdXWd8uxZA1WVE0WbSpjx
THhndyEQdGxDyVda2RQvYDYqmhiJJsiY2dF0FDHfcf+IC+2ySOpNR32t+rGzWFw/m7hxqEraUm4q
sD974PO4neGgDKG+Jqj7N46VY/u882rS/s8lkrj+t1ntJ7xW1KXrxijDzwCePIeOiOkwDBFjCsf5
GrRvBUVDXXF4tJ+IzfSOsyHgcop48qnXlKZFWX022l9/AiXsQEbk50yr9Yip6gXbmqou41sA7MJ5
+Yp0vj75i7uBWyJASGV3yE10dxKPRlu4v3DdyEQxDeRqKjQkRPEcfIaW2ZbNeNUNjXZPmc+cX3g6
JIQWflg3wctGOcql0Bm9nRzPz6w799d1sOlIxyez6UfJbktI5ZJYTGYfgUqM8EjjFaAXCNKUhmKO
lGFOLcB4+/W3f/aa9Zlc3fc7t82/tvQB56KxwUnQ8R585ikpRXkJ3wFwmSrN8U8NUJYOeT32xmHJ
mZVVkQ9XPOtwir6zmnY8Kkwk0sxEspc5vCC95l/aR0tjuI/CosZPPPw2fahvTXA2Hw+5IMIoOUeV
at3Am3Jg8YJyvVcFQOnNAb6ReL0B9WYCA8qKTql8KGDVvAsfZTX4vGwYtJI8BZ50feVvPW+EU/oK
UzKnubsnWsg/N+b3YQf1BxiFKJBOsnKdjEiBEMlu0QYqxcBse1gVXOJJssK2eBjMAeI7tmnONriL
QpzrcjokwWjh2PFJehFVAr/cnfY5ili4h8GVveZntEFrCv5jDWUEWMSRDXpdBL0IwRRRJ35dPYhd
Rx+R38ssQx0iDt9+iWJT9BPXFxeSSCrBIi1WjHxMZJjCJ5MnYSOoantdnfZCLb/ZvFf2Z/wS3u0h
ii4/aVVg3YvS3+bXRP+cfiBhwxtRFymAcOsbeUBM44XLIHW5G461XQTmPi7ETEnnVHTmFlCEbmxK
Wvg4OheXZTxN3/RjH3BpM1LTwf1z6+LPm7TL19nnPFz5pFbjjTXECY64tW/MNoJFrMpQ8jp9HTaS
F9xFN4AXpI8AT4C6UgqGVcM0kGeZKliXBtc7M7qbGFY0cNZF4bBmNaEDdAwb5JM4QL2Rt/7z6Eqa
NzSIv45dkQLhbTNlBAxEkxdmIXkb/Nbwpr+5qqn4aJv7oMJuwUWN4Hcp5y/7B9JrZYyjacw7Hanq
25miLT18ULh2nUQRdgH6Zg00HspM3U0IjICJMCZyifrG0FD70uA5bqsq7GY1XI1kp9oFcM8OAGYo
NKA1TNaRysGGTEVp7zUZa7+DZZcvrJx032/aLNLWG8gf27m5/gIN0Fg3hso9hh2Ac6NVVnWbENzR
xSxeK58EWzVPo9LcB/GRhDi749lysIZ+bdRAYI9q7xhTkOzObW1z+QmMH0pcMoC5/+F/vA4tWFy5
EthhS4pZuvdz3lJ54aOEItEGBDIUV5VeymscsfYmoO6YRcod7rmzwVDpoGVKphuT9qBdzGs05HPq
J+ZCxhK3lC11bhDyM7jznGuAqqe6CzfMCAWFhfAU/YnxN03bTCpZWvuSJI1luMICmSB9NGRv93Lx
rGdWjjUVEJFygxT+b9cHltzeracoZe3M9wKnrNCgvOOaksUHoDa7O4KYEbVslzjF3tIPG0HU0/RC
URk35O6wTx1rNQ3cPy9uz6ePYVos+GCoPLrwGDYuBgK81+2/pKJKXPgVOeTfmpNxu1Xrl2gVLOzY
DGp4sxfb6VL9mPuDjI5E035y+JmxPPxsC2XMRcBmBWM4heJoGU5RT/1t6LWEdMmz5X6jSG3lc8Pf
0WwrVtdMXGk4fcxgJjM/OLtwjU72xAiXvgG2TLPitlqO3vygJ4sLpQH52vM4nIeeI6bEGJttFzXB
mPenyDz+hSskIR+jJATHL3Wvs7r51zaESjBn3rbJ3Yv3UviUDTY6QGrhEprjmgs19APbVw3FcIeB
8IY5cAaLac3nn5rtFc8/NCjjoF8U/69G0xXGSSAYNAt0U+Yri+Pc6rVPEUPB4U2A5keQijGMa4TQ
/6/2IboKxcSeqIM+3d3K/xRQmXL0m+rrRv0iNwPdH5Y5Ygo4p67w6R/rUFdhzdpqgYhRmjD4fKj+
wejLTcni/xR/rLfp5WmMRzbUk2N2MujSI2ym45vgYrQI3wPmgAWnjQs8en96Tek6s6AI9Oxkwxs0
+WX4kzfPXryuZsbbzyB/MedzN8vkrbskTidXtU5MyQAdJr5WUuf0pIRPQT1LZif2bdCkO6S/O/t+
ehcefh4nXNULewcfXhS3nrgGjhrMwBpKXwDKz+BPZLxPkCBnP1A2bPHhR703yzk3bkXmFIxHHSks
g+wGkgi+PopuXk5aYx47TtXoSNVzfigP5ZoYvJfH0F4gCvPv7xpTZFAZXI4+Jhk+LXF1WQutjsFq
cBoptgpj6AB6pDJM3OMX7YZa4PUQNSVJ3zhrrW2SvAMdstqwPnvjBta0Lef3U9tMVkwPAoibZYzZ
0TL+c/Oe0gmt5hV8lkZBx3sOQjVZYTRnw4dx1FzXmu8JWRAUSiAN85IuLxvZh5RoGJRSFw+4fV9j
LEBfFNzfWvuBV+U8WlSTlNZSeF6/BjGC3VkrJPge2QHxcOVvXlJl+VthbHEHezmkMtHy6/522R80
BRdXKOQOL3moNpWHpzPT4xIO50jbpkCvrb6Xwh4KMA8bIGB/1WMOJXTVOmZAM2qg3e3KOJSuknqg
LxU7oSw0PpZbwZpFLm3OeMrRZAJAVYn/rsiMis8RXgRdtx7z1tJgOBi6ukv3kQx02+DpjjOeRcnp
CbRdptD/KgIOOuK6O97+HqTwAWoriBzfVAzR0DZWw7F6dyToWCrz/hf04MRpJTi7o6P9MWaJ+FyH
dSq+cTgUpZTUPl7yiWzF5NQal+O723CuOoixqLLZE2Qh0hwqdsDUyP70XdzSxc4rtyOwCDiiPxDn
Mphca+RFJHJBjRDBRpi8Vh18ni2ADF4pBagf3M2gnjtl5Vg25hBIFEh39Df/MkTdeB6w7jWPfduf
Oo+vWzGFPyagr/MdDNWBRq8qRniW3OtJzYemjs3ZM/UBt958A4ev3RA2p30laLVi+Mp/9Jloqf1y
tU5Q6/Aj7Px8lBKYBiLOb1sjkEldWnRJYHGIn2umuWoZn3DIiy+MqpMOp1E+jmdhbiceDdgvhhsS
mgxWkBOrtV/xvlfNFxiVoqQWkFfkqDlGTZWMb/OadEJBQ7+GBOWceh8D5MNz4mskHd+flFqTBCgk
bPkxkflWnvOAcbbnmp9WYE90GGTsJhURHv++b4uZlMZVkvZXk7oZUfKIHNsR2LDr1GCvYrc3nN3/
pt7X5WJ1FMjyTqBSrhBRlmMzk+08EEVFxxgML8zGmozQkQAlUi0oHwj2CWwDl7FCL0E24S4Jvvyu
cYd3exVhn2NER5jLqYkRFqw6ZbuegDltH8Plj5jx9JFgLsaCM44Rt/YshJa3JGvxvHGr9bS0Jk3R
3ML0gdHsyuvG7A4cSfd82xRWpl9gcpu9g/YMtB5V5uG7jnf+6HWT3rHgYMUZiSfcqUTDZtyZg/47
A7lLVZ4PGuuye5aB7rj+Qg6/BjYHzP6ETYG1toR5LA/J+m0Ovr1nxW9TNFOMblcVZBXqyTuAYfon
hyNJdcjUH01K3+wxfc7l2Qrf4hlacEZjzXiTBqQoXwWjmaFLQgjAZv+/x82ebOivenXHKxh1bcJo
qJ4YTOckPNFStNfKM8DdQLPtm/MGDvsQzpWxcqIV4aPTIHjZjQa7DpugNJjVD0BUpV/+hhidUhpe
ntMpR4b77ULbIod98gV60SvdmTAi0FkSLOTHb9ubkrE0E9eZ2gEBwnNKk7N6WEuTCj6j8tEG+692
o1ZlUYDGX30FslD/o5Gdgnoi1JaGlAYciUvKqqwFpy8Fxgx+MIP9SOKc45Nse4VwdTJQVyrwunnI
eALTWfNpMKXYL1199Ba05KN7pDY64QmkMqgYVUQyx0hJna1473D9JIioZWaIfMwVfwzRMWrc+/ut
YAPYGLL2Gq1nC6KaJ+JuHxsnbdYLPoOugyFZIDxxvvx+NMpX5pYByki3wofinzMMWY9Dl1HiDWu7
aKJN43Eiyr9cr9AUN4lDsawWezIDd8FZzwY4NWzQb2tOF9/CqVO+lqvrhfrgMAXFqc9Qlf7euWZ+
gLzeHoloZj3Oac3MoVgRwNOXHa43tZWdZABiJcRfA3+R2f94q+KtI+W8EzmwEwtxqm2S7YmbXJtb
+pu3UXdFWAZMtJ8oF9hStMM2CPrXoKYSGIQSwnSE6lpxW/1a/FR7+Cq9WtC+lE3TTmsLzNJa/i+R
ELpVMzIJdgpMxieyRyeSVqpZdxnVUxpPoajPr3Otpxuv/V9MUCgDtmphfjbYLK1MQ6Jil2PSEcYK
UhfLvNDVO22S2lgxYJRVxkPy9QxgI7DkjHrMgLgy4MnvzMU8Ld0USUYN6OtH41OiPq7hIl/a9K4k
Wg2vIt9N1uTZfExt58JFV6idPOVDtWf5qrZvjVd0PaNKL5VedfuxVkeba07yLGpZnXkH6xcNn6b/
7y96WCJomrId4QoCFvJWAVrgCVNstdO6QwzWXCHb2HRrI7WP/lncvuQarfgX/4J4c3/3tNABAwTO
RVBnmtrinTSJ/3dowHLxpJ6HO5VKyRFakkwD8XRCV2PWv7cTWwkkggWz+2KR3+yCTKOVtt7UgtsP
Y+5kM/b8y0eqmv311uz6Vpd5SFoUJsmctp0L6kkDv/RscKbHmjC2DwDkCXCDugCzlERyUqxoa6HI
YWj/yjJ0Plkhj6Nm6Y8QfSYHt+h2Mkzfdmhc/uzJHNWhp4zelcBwvsFABBC5QNPVYoNx50pku5Ap
2xDtyIjmjGjGZ5KrWm/wjlZwaLqtWniIkNFgNfHcqXzUxsEx5PM54PqDw6J0W2mYcpE8rZbPjELG
hOBoCpmY0z0WsS26O1M/HYw8Wl6YSIlXPK6JZ/+maBQMZeWbfbyUu+o93mPLEpLVG95c7LdiHwYm
dmxWTmBWA4DuGgsTwiZzZKg/mOk9W2iR2qzrqaFK+gBLg1n2vXPGs2pycEkNj/k3Bi9i/f0UWw0x
c4n5pwDu1/k35Ghp14QDgHzUGTFqe5k1EbjkzKJXsR2Wj7XPdnKwRX+6iRBPNZ/oHMNXGx9I3pak
XBg0dCK8lse3CWcaxUQyJXcB6ftffkVu7XBRf6ymF/mnH4kMP348eLyvgphFwW9xadFWlLdSGAnf
xVSRBli3CoPK2+7Kcy64wM4usxDYYaaIRzkEkx2F5YBoOkGnaW+yMCCo3urC8bXJxq5mNBSQJAGw
LDltUvb/fJBRJ+a5u6Da4ESYqyRH4Zp8Nv/a56U9iVCnMuaIbWWwbNrVZC6nD9AXH7mXiPlluaWX
ryhm1Zh90D52c7tSiz/t95riX3WUeIRouPVU/NjF5SSwUGEuZvbRO4iGw7aHv04dwxd1V4eySlYZ
xZ7sY9IzGwObWfwvZQeXGPZU/VCFRL0EecnE367dv2u9i0LnlNvDjqUWH2Q48dE22MgXQr/50qBL
E8kslX+cCn/G5saNOkDipIfkEuYur35hV88CpJ/UV360prQuIBZTRvnSCIv9ImGDnManrdnDSMWY
q89wOnQcpwXOJX4MPXiUU/na8mgMvRwiZC8zBlWA7FL3H+n4jdo462TxBNvuLUGJDeWaDUxwk7nb
hiBnD29FgMeOMmpSd4ApcfNZVO8X9yf9eVchlKLoNOCB6vMiUQks6rCyrPLa3cq4bGgZx5bS0bFy
BsiV9H4mdiqSldsw1VZKykIGor+bnT9rBMUbD4a7N+69+n/Sd7+byErrc+GjsId8tMRXFeA5bQzk
J1N6SC7WRPy8NmHlFiY3tRsSE4Nou2YfcGYMK2BBxwQIJB3UjV5RnV3RcBECXTglpsor9/X8AsSL
Tds+sDWNTrhJfTcVVzr9NwVFkMY6C7/DTSmYBtjN4Je627n1dgb8JfI+VLBD5n4OjheOQUS+Zqcw
YxQd4hJNEHSk48sU2f4DgVtE7xcbVr1nF5LgtS9hpyjhmMdyUMRu6aG/Gi3XLgk5qa4Go6W3DSU0
/v8I+IXMIWxtv1VitIPL+e2NcVRLXiDiGyhR5BldGyF3MmAmeyy/mRb7++xHXxkO9T2NhGGtV3ok
t0iriKJmQj2+cCYmOrwB4p4pRPEtt1NsGQ1vrsU0ENog/nNUUClQFzSUi4DlyXSnrmlP3onIi2we
vlcEorHDbZjuAJvj3Ypq0FOfOBo3CRuCiKT1BQTF8GtiCyzdNxSDIRqRQLWN7ovFMgKdt4StpV/5
phSWM4nQg/MQdSU06OergMJOlgPyafGeQaUBzlmYl0+jSmX2qRi9f99iFOCf9V/wEtt9YELzRlG0
sU+8+ORtNSy7jd7Hs2wkwCyaK90P+v/SuaFYiLUYtKP+8/58UeOqVXLTlVZfqUIilVVo3CChBole
AvT9rN/URYcU3CMpACg0kS7Lsnoe2e/wbzNePfk6Q0JY0JknWRV0vK+QFaO/G0+t30hRlIxKP4oc
gp5ZrzEx5zTby1zVoxOWLvHLP0e/FW2neXdtdQW31bk+TffyW/gFLrh+B/zBUOuN+Wo5bbVpxamM
tTm2PM6uLDmQZbZnYHFVKOm9Mq/2HyyxScwTjBccp0XYuTIN1ljSwof6V9kEc9ECIPaTNVPg1Piz
Ksoop4R7uW5j5Zx8xBgn45pvc1A88MVajOY+c/Ruiuz5yAkRSv544Kku78l2Iijwl231CQoQqbJL
ioBJ+Mx4UqcQLwGq/y7ygHH1ycRQErcI0DIRZXpI1UoQx96ENn4GOF2rMHVSVyxwoDK6Y0knuOEW
h6fuj49md+gMI4lHaB2g3Nen3sTLbsCDX46qXfo/RaJi+9YzwzJi2wb0/yX8qUNhquRc0MQ9cD5M
MY8MqkTkzrzpHAem0oyP/UqPRdyAM7/HSDuEur9Ywy9jLAHd7UOZqdx0V4nxu69nHwVvk41Iz1LE
J9r7p4b4tjzFn2jHr6/N+1ZECtxAI0irNLFq9iSUWkp7mTb+TzMNm+KTqbE+vVT6bReISoq58QHh
E8fu/z25OAIHlEmJPYntI73iFAmC9KBVxR73zSDsW5j7642O3W4qVUGMQEKuiT1hTPEn1o6rlixI
DbXdjv74LPaHPNyF8hlUymP2p7T4EE2iSkxZgY98627DoG6jEuXvO7yDQWc9bt8AoUGIPIjCITgt
nNHDOtPhEyyUxw1m2nDqUvIO8wrVC4f13OOOnGCUdQ1sEdT8c8uvjwZYMMFWT/6puw3XBy7/3Y2i
ML4OGheOJST2opcVsAIA63jAq87ljFbQes6RvPlwlgK9JQaFesoi8o92YqIjRPuK8LEvrcPFhPo1
OCo5kA2IYwGiFS9R/2Yv7HFl9+UfNr3DRU5UYkaxdYOQOGwck/zHwMtynWrX3jgmrXei0ioZH1H9
w3XO6QRZ1eZZewTel3GseubwEaJDtX1ht+UuVZG+yXyHqruyP62Pe3Mk5HFWaiqWuZUKH9tpbvMj
BfFloW124QLV4JgahsOpAfhIf2VkKlVb81XT/9A3A319OKg9LXbBycZXqSBgCVAsSO4vTQWGVz2V
K2HxWeA0oTuunbhl9FUBafUr3T5WiP4NMDas80h3cg2tcXmyZotTAIU9si6zR+69PchohAzDGF3b
ns5yFTdh3cnYzR+qjsqA5iziKF9GqJzC5Zza9TFT9QLKmWBh1D50MVhNXeWD3Bkg1M+tcy88ZW03
ZUtlCxTGjB/oqjJcRv/rG9cAQazi/uU/hHaMae2wvQdRhwoVXP/vTcG7irmrilssgePLFNGGSDIB
hLW/KlxzVRtic/vcBVWRmEFDHoopqp9YHgAXw/gd0857MLUvqbiFY0OXasqC1wsjhM6rgcx/C4hY
wNwTwBve/l7ZZu24FQqt9sGpkmy6oGch0Do7EDcpDBu/C4sCX41Toxt+A62tsDKqlXSw1bTo1T96
xOLk2g1+XaEfdbRTKRB6TOBtZcVUpAVAoW8SnGuvDpmdUPesTNQ+bFSzx+5Is45tp5WLTDzFIRxf
8dVjDuw7aDBbSKxkTzEgEX+n9T2UHewEMnUU3g4SPZVUEtqdAE6pBuYFqjd3zF5CeQE1Pd3xAMKW
CJeZ4ejQ/Xp3Em7tP5BnWWXwcZbqE3vtA610/UjSdmb689WwIVWjnzDCd9nNAg8br3Wz/BU7s5X7
ZSmi1yaz0Shdg27byqwD00+bfPbiCo9Y2DV60WTo+/NAzeAa5xNfs6JlpTn2USEqaI7k8qePLClG
EwconJ9wMGMtBXlSKUukxKbjYL8T63Q+he+wsX5qpAFVAxhGWpg/HageN2D9yY5oh5Jz45fCKune
rEeObZCc3zHv2SFA4FCTq1ykkLb04KaC8qVM0uktF5FDUgRo8KqFeUcmHZn59eNNAYMe7jaaFUCu
GtvVCChq/cRhdWz9fZqW3zeFSWdgrgnLqfmCAK2m8v/IlO2abHwesjnTHDCpH/ajj951qtCaBL+N
6zd6QkzhxL1C6IB4pVTtOLkSXgeI/o9P4SlXwkdTF8cX52lz6ioyuZ4aAGBRyViSJ8RNzu8OpypS
4GWSXQ9DZ9M3mLum/E0R24nTi8i9UQ5KAsuNYkj6VnEMETaZxOsw8Kq5uSHpwWZGt6PLGQz9RWVv
DloBRqcFo0g4s5w+a6RpeBMetwDdjnzbXfa3FzScMaOrL6CHEF5YNd72xAHRogz0LEtfbq6r/znd
KgMP1VDbtMxa5itIjid6ONWIYG1EcB5AFosxKTplwLg30m6g+DIb0xmth1ocDwzg3w4Ofbi6V+Qi
/27y5GZeJYjSRa5pnT0YFj7t6JrSTSPeAtYODP9AeLEudL1+QiH0j+Jxo0QaxXeRa0KkFlWNHF2H
f6jidDoeAfWaICmrdJhmy7CBnv5JN6v6Ezk1gB6MY+YY6UfDxioXvWbPeqb4EzMn321hMZwdIjbl
nxr+a73imJoFCmxT49xJhaDpuSb+Qs4bc19jpOGP+UFGFk+Sc2MTGxQWAuPym9JIsQab90z9YaeR
NHdYyomcC/Lz95dqc2KFKBEku2mP92gkjt7hjEzgQSMp+j+eYfHAzJ2CExWgEWwHpCSwU1CGRmXW
xvUotVLRvI+aMwqB+tLeZF7SlX8LQ//mbot39aHY4kMoApQ/vQUUij5b/xgB6n8idnZ7UFCLQcBk
xjx6nr71Z8XapL1FVg6MQY2iMFw3is3rd9NnV8UXO3PUhwdMOaFRX6kG6AMAMUH9rY7fCsbRXEOX
qOLs/guOutUL503GIx+cObuYGKdByXN6050rrQfb+dmmwNR/jRvbwAf0QoNlqNR4rloZpgH7V9Lp
ll2bbU1juaCRMnrEg03+wrD7j+ztTiCYN6CaBQRKi/cgACamBfBM4bfN3D+JeXF2CZ1J7NugI+a8
V3Om9MFb0Qnq/l+ggvvFzDlf+99MkTQDFxtEvTErVqbDcwXOwbHMWARwsuPYqv4oJZ4rbUk7HdTJ
5mNb7F7zZF8w/0PAB9IRIH0FNiKbSaX1ZqybkZ2fFfgRsdOujBz9/ZBW69ELjSI1uFoTihxgsex2
Vr4toVVKXBlIZFXdTd3myJtMnu0Y2CuWMKeNDhYGyOy7Ym0uIU17+656G4WEPQJBJOUIEy7dRmuV
lcfaIffpzj78x3/Ri94kOm7BegowrZOCcsilJyo5vynTWcX4foOkTiUus7C1I8ZmXtdidbFS/aDd
i7LYLCtwh3Ii7yK7UoajNBRxpA3R/jNoOhZ2IWcaenH6f9Ei+4nCIvyFeRj9b8rcAP+hP2+Es1IN
JkeNneSeHy/Htr5Oi2fridBTVKrU71tBkcb7UTy1a8Nid2Zuj8W+WaqPJ+IK8nUudKI/3aiIvKTj
H/MVXQ1krWE9sCfg8OqCH6KaHGRSYFKAsXbhUnr+fa14pJ/MBaw00MiV+KDmCdb1pBL/ef4sijn8
xZyN5N1hp4Wo2LcFBLahSsEaMJVz9vFbgW/6g3MBkc5VV3g/jguBpMMln2C8FL7stXvLtUaIpDWl
z9luDJ5mj7MjHgF8WC5uNanXRFoes6HCUo6IXps3O8fphWR3q4RKs9hkYUAOIy5TPhFXgIxffTD4
hiFFOEscNbjMIng6bnY0UnvraXVgfEbhGKO/4v3U8ri9Pi7zj9ApRqX4wRqZ2kgm6Q27pAooXNiD
VF7kR9muCU7pY6sZRiK3I55oSHPHkKbdt9tyujMCeC3+OgsTGWXGjz+x008d1S6MEt0Mbg0Ofw1W
1CA/MTOEJEVIJywA2WlSI0pSj0gt1r9hx43/MVDGW+y9lsJrcuraA9PjUrS6yblg5a3+9Vjzb8Ck
PIQrWacARV661NEEQ4iySccSliC9glwKRJlgdVllNxwfJV1PNYOnedven6eVzepyekQq3dS54+Kj
Oj9k2DYLnDLajpIJvU189+L+wq6qKhyWPP4q/8fAxkcIqu1AvnX6XAOyEFRRoZ5OY7eFKLLdL6I2
+JH8bhPhLWKp01rtIdvEheyXXjFu7OVBSm7EF3eIu4WIjZPwH3GMtacS2kxyfIalZnvKJWtv7xKK
TFhQymVybvS+hwF7/odwtPbbJNjQG0fZE4fP6FtqRX3nwg3rgsu7Zo262Jtd0nnoRpWavZxtZn7b
njwacjEwaImDzszECE6THpfpW/AqiTE1Q7hzLnFgCm5TiY7fmWMakg7w8MQTla7VcVmSFj/rewvd
5uJV95yosDerp+300/uii/GdTulA9RRrH9SkZYP5URDI1XRzBpXOHTW5qzMxoL0nlr6KRFq4tNYW
xeZac2sFYb3JrTPs8KZmEZzT2rQv+KBtEQEhz0u7JP2xUzmNo6c5V2DbV++GT/gpV4kOyx/ITEeN
g+7hBxaO5QUyFETwZVklKE2/bemG2b30NzM9Cxf90bQAUsNdByV2UhsnCA8gmfieIAtt9tcYNls/
J808Vjq0Keyi7xRTCz5N4ormaHn5TT38HTLRu09EPMrrAk4NTYz62HQlvr2yGFcCUNHjAejkq6ix
B3pES44yQiN8TJRGyx41DH+mGfim/p6VQyuQCUG0h9Z3bHeywSPCbW1ts3+q13LGfRJfGwZzPErT
lZEYlUGd4tFjfs/eR6HkUTWzQMbN+dcWo5lnA4Zpz0qi+QlCzYnk2afdk70gyqyY9nPWU/U9NtOS
SFURMolaO+3JGzb3z01nK+8DaCygBzL/I1R6zELtZY4bMsohdaWwaSBkN0Sa6CLLgSKc0NQc2DGX
qROHsZ3mBFE/6bF/TB2DGe4OzkWC8tibY27OINGjvhbNOk4UeBNQvpgrXmoh+tqake9ClfpZuZDf
I0gu5W9cNKUb1TY9XXIcrGrflUoAfKF+pDilJn/vCpeMkH5nKMyXesWhQAWInGh3iRynSUlr+FPO
k6SShM6q86H2BCMUEzTINVOeAZyXngLlxa3Ipr+Dy7j34amD28JfHuvWgpNWAYAXOL1C6nMx/z/v
POHrLmRNWwuvtGPN590rG5rdsqFhEWwH2MnVtT17RrRxH/6u029yqvN1uuVPrBqpCePte21vBPtp
TF6Zb37fkYEiIzkO2yBKXytKvCdtw3Zr60bwcA0vOye5RNn/YWJILPezRT3ISt72le7s5x6HtocD
/RD5wo5q6V4m8fkJf17MKMziKvJQciz2vOqIYxw68pCQRqLIrNbRe46oRjv8yeZnXvOVAOky+khd
OePYHR5yLWMfRMWuJEBZkk97grsQGVeKui0+9sjHRQQ6zzyjT/WBdfbRvqRgLNL5Io6WrESWmehb
20G7flEdemawj76C4G+Y/0VyugKISG6OWCXmvEZbQaqmVNPL9gw94VMPA4+90y2MyQIxWFaeehL7
Ql3bS4zaWfBTH1yvPoIOMijrRegnJdt+ClhUqtLdwVL5XSIw71BoN3Hy4dfvi10GruAQr0bn5Djo
LK/XUaX/znAlJr4QC/0oZMhw8/oCHzyBTTaGDQS3H73P87fZkas13ZHHTUEppMN6t6S69rFMob/H
k7wDKxVNbZhSkfH9Rt82qaVHGXE1yMrGiFzI+FsJnoKNu4RavLCsdk6IbA91YOAhIi+0PPubTQsd
rWLbTEx79aws5/lFIibMxwKA9KDWAE397cZ73oj4J18qHYRQeztvH9GuXJVOAQO/VhMv0tyNV/Tm
oEfHF4wcsycrshf48roS58S5A7cbqjIO6gigqJ5GxXLbAwEf5PeHH6Hmf9wXeUthNPMBsQL/QZtW
RVegLp4kqggGyMFPDqftYwTA0XOdee+9JdkGiXsHzq/JzED/5zDFzkWQ5vacj+4egLBQhm+PsIXS
3lWC7aCXB91RWxIJdqKtbHwb2VVQvpg6UnmCT+Rd7ws1JFeWBwJTY3TUANpKtkzqD0GEdqTwRwRA
DHlxRYwVieNReAWVO9ckTmju6Zfic0vtu+47hAZZVhzkWu8fpMHje23cKKZ9DJ0RZ/6xwzuXLYT4
ItW4m6NHqUyTjuffLGxJ1P8JmlEtsMBD3zDAsV+OtYxM/Be+CxiyXgTDdR3tp278NFJ+v/bBL+lw
NaoU16XOdR+nigkmBnd/T7bZ99QKSDKzkoA6kCvHi0yqcCZ2LmNIqCdL3AAn/bXxet9Rt2wZPrxb
WdkwJ0ItTGF0oNbdWGXBDQyDrO+CDKuXw4dsLafOvPd1+CT4vvQGoCYaNEPrqbFPElFEMMD8m5lF
eKsGbVjHnYfqVmqcbpzCpW6S+gOtkDUNUU7WRewHZwhT8ABqj76nBp48L/s6E08lKuoOQmLurS1p
hMyXufphT1R/TzrmEkXiRht+1QTfCadwZ74I3CtpOzqfLSBiL7v7wUAkLy82OVSze7VJNva6rpaF
OFeYc/VlGpH1mi3uJiUv37vN316x9ZXMQZKpeYy5R0Wms6P5T6R4iFAnYx3NmRzvQ2Uq0W11IFo0
zDSi5IclxrjaCGNrLs4mVMeRf1yt4MOWjmA26SclLvw8wHUCxPQ6/SBYlykxwG9/oCLkfJ+QSwCs
V39RJlv9Bmr/DV5xPivj2g8mUZa9wninLcwcExd+XeZt4MY0MB8M9/YzMfjMaQ/DExLT/Bxot8tX
zOsNAlBw7M2g6NzRi1OF+i3Rpa64WafKr04eSWUwmTAhytVs5DQ2AwE3h0wqG6pJ8hBFVoVcSUYT
fveGX995MkaxhueayAGA/UGhIOcxLgY+3iLpJWlQapzyumnZ9Kf1TlVk4FkfxlBUSKysec/96YM8
E30QQlhki8nkfslflAVih3PI+ikcjFgfpVJXY+iDM2VBErikjZMYOGF6zleRvmXSiHn1aKrJ0YtC
d/4nYvuSS7W/sd31XSFUQ31uzQ5hc+OnGtVdGIquXJMw9BoLQuLhYfSjqW8e+6wDzS8Gl6Ag/h3q
P/l3Bv20GG2jBVbOsovF+GcTtssqB4LuhdzICLWCLbINZc6kU6MMLHRhYXIiyLQq5DKuw8mGkeff
dHOaG1ZA14PxKZIaudy0Zo6qKAhPFKUbzuKdzAa1jQClCZDfk9/dYfzYs2/sH9P5EX8MOzrmDPKj
03LJSWBQ5HwWFPDnyLYgvf1EGvI3zo4WjBCXxlGviwpAzVz+0MxZOPGisItoLlAR1oO3Ip7Iu3fq
ak/hinW0m4QsfXz2wQKXnb0AVGUw6pQ9AWQJijlHwzX3Y2jpDcp+61BLOrZTeZG9dulntJbWBpoL
ltmh75LRxlQuQQBlv/j9lEi6zcdmpqmzbuk3m8MfAsZCOlgpSQvK460MS68haKw1cAiYm9dYCJ52
RGJJkV6EBbDsG2LNtpIwON8hnJYhPAJuGuQu1uTsIB2cI+tHCi/OmcICfW/702BR4E/FWqONg2Ao
zDaGEyLSysulDJhsAI47xoSF+mgNZcutB/az2RXd46nd/wWyDhmfwaiUWhX/ZSjU1efaIEKZT7A9
DEPVKOgeDRPgfKrX6KnBpcmCT+WiYGCsWhbbJ+EQb14+2OhqlBnWNL0tVG6QiBb3DVvMmdPt8MC1
UiaBLMrW67YxzFFMPEtK6R7sdDH9TXQQepbyEbXhJKkGZ08OYQ9/mPZb+0UHHv7cgF5KK6jn/P9d
vftpxVDzYzYQZJUAEMamcRVP3QJN74KpmnGBP0P1O/A8tFdTs648NE9ZQ7/b9VE9iQb6ZxR+yUTV
srvglRwj9zoep4WYIgW9VUP/YLRsnOlK5TqEs2ohj1Lazi+++SO1pcEU6vLu40MysiZaZm0qVxrh
edUEay3nSM+X/YZ9eWtcZ30iQ9nAr0fU0UtW9Ut0yF6DrMmmYahDKSzTI/HSeAQi3zWRxL3WsUIa
2LKqoZyxG7rqflNeEKeRHEPrDJXZ4/TRFrr9NmYduo1rTjFAOdWbxKkyqKidy20NqPwZiOgMd8hZ
fAlsDcFyUco4XXNAbxZbWeUYqkjIERKwvQ71kIM9QWF96ctiYG2UO9GlYSBAd36ntqISURQhDa0w
TS1Q390ZAgZwld6NxToevwcYViCfQs50+u0ePs4ljT1kHnOtcE9PW5Sh+vRC1wdNCH3Nn5fjUy4G
gfzFk/4UhTy2xgY+NSYeqjG/5zt6XNTE7fonbFIpn1usGSQS29wXe88B/GmfWG9UJO6fYfhDmtxX
J64AhQKlbJWpOuOII0ASplQmLSIw4QKd4mdMMukr1PdRNe8dM/DPhN7ZYtuDoNPGYHCbamAtexcx
Jde/CtXTEcU5I08EwQ5YUkHn5nmPCQWrQtBtsaC7tnqeT42i36e6dM2bbai8r3Osp8PGdc5IUA7S
jw1vbwwX387j3plUFmadmatAyANlcsPCeM3YPTSLrMV1nyibwXzEaGZ+5vJTcED/nxNTaHczVdxh
OHlfc31AeoR8qbuRrZ+bWkjMrJYiW+PCgewg5zf/fxVid2xPnYKBuDCmRrV649YxxOKKr9HrhxHk
NfoCBdhX2UhyVpbYurLRmzBw6bPS4+rJwoqGQ8pXt69moxzn35RWTswXtBbMKdLQ+0UfOMJwPHLg
nobr1BR0qZhoecOYDToHaCHlcD+GXYlVslyCekShHSS66LhQtDgAHZ1XzbuENswuuZerq9cUHTjL
96G91qyeXPk5mRogpDlvwTN5HVEgR+hyps+pJ8WTsJxjBxN+OflWEg4Seo+7LQJiYdqo5z58970R
QYjtRX32maTL7z63dXT0DEvvYfNPCQCiUgefrsfVwz+6kcWmAof47VS64/VajyGoGGzTnkOTq4ao
rx4u8yg+FoaYDNIWc4dNoAGnRX8icYWiagPdffZsitBwI7SimFd+BaZdHgoI337PyGGioV/DGBbL
zZ8dtEdp+1jm2RZHHyX1uxfvVgNtBgEfyHsaks5ussF6msjjQfgJAkgwo+r+5awKmIw6Wa6PVcv/
gOrCf1xn+SDIwqr8jxlOVAyvLhXP4lJMF0eIPv/v5sqlSa+YCdtLOam7dRVZca5WUadBcv1bqMb1
FAVOJALC2hmTxc/OaWn4nt8qBYI5Px7ptIwCIsCEAogmXFIpWaDY+R8JqNzJ9KWiBAUijelvRvub
iriCTTJKeDZMYFVQI052rtgBuHyaYWRt/yWPveDjqIQgSGdk5TvgaAXQ+hfzwJoWrdl6mTJr9BSr
7snOS012VZHw5vgYsFOSMG4YqwP6iMjFRDi/8QzUe4MI1KwNFV50f6NN67Sctz14Gjz7aO/5it46
+8RWhIC4HbnYpuKwbyg0xFZD0WO3nutWlcKtXl3saxyJMlbnQRsWoqXJnoc8ckB/PXwkFSJ9pd/O
EUMvxjr78iqWJxUVs4u7YgFomuEvKCSqEdONsUtHMY54RMdNEqKLH0MdDKYRkEWEROLA2JU7Exee
fEb0btn/F3J7XPyfg01aiSbfjxN0668SfAvd+pMqjk7+aCYJg4XthOW9BaYGnoldKDF0uh+Uer+m
VfOEROWLATpIZXwVDRgeIubEVNp8xa6X+QnSX5qCcALb0iBO/zw46H2Yq4NI/AtMdU7jmF1TIJL3
0B9zmtNTgANAI0W85NDKLp8huJqOBJpapWgA7j3WJjB/hrzSzq2f72HaH2yBEW29CWbhspavaI8Q
FsEbViOysLhuSxv/AcNMnL7fe+tmVUB3xwCixv7Sh0zvKZ81j4uoPRrja6hxgT0NFsuYJJuiF8Yo
RLH0Hkj3ylkIhrdZzPNF3FYyqZt7/vI3j/QNQy/wGrJVrpQlLfAYTvWVCDrH5+N/q7v6yEv0cdGA
frsOAAqyz5/BLL7y9ReaMsP6CpPuRbBrhE+hQuQbXKIYGVRBo8j2IIwwGojNeub1rB22kXEL16B4
g6/QGQnxaQ7LuOqsDeyBjsykOtu40rE1WurWlBVj+HbfsdwHephz/PQRbrnD8O39ECK01k0WjSD5
Zb5doWQE4407exTqyY/YbRWAB9gEWcipGiE6WTPyc4UcEaB2UEknmcEgxH8HJDlDw4ciQgbMikOt
P3JutN08Ex4TMtbZOwZ3l0g6b3pHn37cSd5nKhR1lfIVLypYSphoHjQf+HWjedEDtwvPdO7ElcIW
c+4+ZZvUpPHu+PaemN43oEkaIepQq5cS5YG6XL3lyx4y7+sBOoeFxxUGTAnInQiCHnSAGCSvwoi/
Ej+kEuY41FV0jy8HNFC3KPfaaUGCp2SZztUJ96Fmj9QNo0QRFyzbOwvWIsC4vLiIaGUmyQjzhwXO
6YNw+nvpMf8WByvDS+AawXpv/Y+27aB2M2z7l6P4ZM/3es9Qyk9C4xpqwgkepWFt35oiLtdhOG9S
LXHKL2+3MwWxYTPruEKVO0ZpQPlqkrnVQqsqIZwHDmFYOyVUrmpfxaOEC4khRthI8MSkWwikOBmH
HrUrUU5AsxvtI58jx5X44GsKFHEomUI2jC2eERYjhfW5gDThdmzJLAM5n0HcUs/1gy9fqiJQqbxh
gSJW32DfY+7/EANjcgwlL8Dp4q/Dd/UDldCAHbVwYJBMdaBRW40AUJKg0dZtUyouyvVNTGcLf17t
GShBBkk+NPww4XJXDFe7s0KrvHlePjETYxcAzvp6CNPVgCb1TZslg2EgdpwjLO4bAjLTPNVjgvCG
rxA2bKdsFBLbtUyOB3rArteao7JHweknpWAkqCKoCIUI+YWTD0YIK3y4GnJ5G007lG5Kvyvzpfxx
L+K6xX8hSOf7kj6MnLzmuPs6lFTWQuWCajd52WSuF3Jp0Cj5nzy9bGf26AVlhtdVdhRq1MQi+IC4
X1E3mQV7InlUhHHTCTPqg6BG8PsFryxAkCI1dbhoa/030B8h1A/YOkj2fGUkTwBsIW1B1XqytxPM
//bn3rnWod3tX4Su9ebIngti6GegqQyDWgFdYr/qs4QPLaQBY2S4tYgnEaRi3ijX06quJzxcNs6h
+Dwcn5MDuPpJE+0u928qpod0qHX02ySYzol4Vo47DaN6leuTQNxS250A5u2D+38AgMCoJtdqiPrL
o2pPa7aB/Prvn7iHXwt85dQD+gZ47mhJOiac51LJYEYcRg+DC59Mno1l8cKvP99cqB/sWFE6kDa2
uG0oS4dsrb1fcRdYFOXZNFuDAC4NkxzJ0OTtfk8GzT7MUQZ1bEvEmEJ7WCq7g37R+Kzpnv7quMjU
3fw72VyeycuO3vHCRnR5l7iJB4VlJJL/3D21lWzbwfKe8rYpkIkknDQtzcLcVtlvIOFU8TFBsVoc
cZL5rNcQJzX+NT/gfpQ1Yz08XN0EVPVQJFWR9K9sqoF1oh6k6Qo3pBGAjbYe5l4u82oSUjtXoIJP
ReBGezN1mSNLiQabap9NEB02R6lnU5n2XMGke3byQKPckqllvx0bgBA3r1Au0r1ohqqk8GFLPpJr
wuC4k6e1SZv4r42OGgvApxwwJcqXDadU3m9cBO1fOEvu/5ZVfyQLubPB0k8NfipISARF5ONIBPgD
3GjUxyCOdB1Lw7B2JRrkQyNLE/4tKnKtnxqNOze+Wynh0RxzmwowQIT/04Je5Ql3a1kk74FHCl5n
wtJGC/ZcyRA7QauniCzzL0jiSfU8BdFOXe01H7z0FZ2B2x+X5NdqgTak5DgbyXHA0hFD9Jkp95iC
71xpvyBIbEqDv7zSSE9a3UcWNgnlb8DHPGjM5llBwRQOgMoDZ/I53MwY6DaU4nccANATboilGFFY
aRhP9eEYodzTltH9rEtkcuxBTAcIYra0wL9FF88U3cZ6JHt87kkKjdFw7w1t5w6j9JheuMcixqct
v6QrwNQc1wedSooD8gWZyk/BkWc5zW5g64y+/kN/IBuGE2Ma1HdOkOxbFuxuCrIZqJhij8vXKxjp
iS372c93IRDg8ktYPHerZFzpRFP1jG967O3KwhOgjaCQvFHVA3wdVSpWcrfC2mnlgk9YqWHRX3bu
XKOrev6fftJbuYJ7txH9TSzvIhBUT7JM10yw4ERbF35ENW6UhQ8EF2PsRFm/xS0qlwnHFDuFFMur
Ke4Nrb6hR/ER63dEfN5Wul4L/IvdI5/3uxI9aVG7gtwqj+qDumXuWe/DJ6gVFmaCNny2eH+Ag4jL
L3CjN4X7ezxZ3Op9qP/zTj9LOzlCEmYlVNpgouKhu4Y2KEyrQIZvk1RgDiPVZDhpQW5wF8L/NmS4
I6Om6+s54CHytLO9Ale2bbj+kT4nWMqnpfp7p8aPkzS8QTjlId/nj9uxPHVGBY2cToAI5pSnl59f
OpH4+4xp2TefXBvcur5RKKTdRwCYNIJRvzOrbv5oLr3O4dBeEL24J9iASe6yVM+zPDIa1kS6fKGX
G4Q4WKCkKX9A8C7AWt25WT4dtf1YtNAOHmQmeFMq1SsjzYbTaT0ONeMgpAGzFz/wTzoAeS8p/lUC
xvymVBFC5q1N4SEi7XmU+Igk0Shl72VbCcbqsicO8M2l1tONHiY5szaVoSJM2dsWtIeC2y7//Lqo
MIyZPrbUaBR/JarneGoBYgRRGcPFqKd+q6lzmb4G0XEXUkLW5VxXy1LHqaw9ePvxxcnu5xJgFsyn
DKNJnDab90FphX0SOcLQE4CVtidlnDynrC5kD0u3jYe+NRblGL78SurH/rMzIEhs1+srKDF2LDAe
QSY6BOlTjufNHpn1Oi8ok5baNMMf91SUUxVX5mFP9T8cGfHf6fs1UUl+R7r8kvfcZBsWinQYO5cW
vElk3+nzH4ERCXmsr65iGnC8MJP+ve3j3X7yiBm/Ap0P7Wf3IV54vZDNnpYcx5LHKA8PVucG7rQR
yYfEWikCLCUY4HWEUNohpvRqCBufYY3WzMDCru87PXXPHCqNjEszZJ9CE9ZVOAbOO9+EAUIGxdxO
N6he8otKxlgUg1A0V1maRWV6tz2NseZ58GM59B/bhO+kwDwfLXFAgHYa0wBgZPbMbbxToU3EtS5a
CZ2hTj/nWYStmILl9MY5u7Ipb0+lt6Y9qTpgv/pYWKC83Y+m2Nus+4KKPr+e3O75kI5cFyloLpwY
K7u9A9UQK11PTaHSqs3VK3xF81sshhdYLBuS78KyOA0xrgdCNfVm/FJ3u+P+8UvCNbaahPViHeUJ
yiyY7hYS/QcYBKwCZgntNsSp3oYwe2KNzc5m7ocX7arcej65jJ51cPKUJQKWSG+ZBIMUR2tOhvCn
HSoyJE0p3zoKSDCeulORPazbvq21gdxFGLX++8C4w5OK2FEaL/mHULNTHpGc5rSXHcIAfztUwC+H
gag4HhMxUy/ccgw0ezaUeErGDTbYUTldttPpzayB8y8H+8jj3TGNxYe2Vkez+G1hInwce3yj/ckx
68E+WLgdkqckjb6rvgqQVe7IDP2xcGwy4Ka2/wiXI8JEg6oRljry5VzQIDFxbBnwi1M51bJ75r0K
jzVhrkZqz+6aqo1RT1j49VdDQE2Izv/r/UhuogXP0lzEtV2QBL7zBSL+vB9HYq5w7A8O5ee2RlTT
3GqY+uE49EiRnKbCcJ/6LPdKICgK7N/wuqsVnjPKNLrWLkcdcdguHaavW6m2si02iRBajADzSk1P
KkLZ8hw0PSNISn2peJ8//gnWIqb2HhooAhMbMUHn+AMPmaUNTOLDk5H7/aj2d0vjYCjkgMYXkcTQ
U3SEV27vabrbETc3znoZqMX279dKUbJe5H8reqqo41zh8L6U/+MncpMuhH+lThP/g+QXfhnjW2l7
ZkiWtsg8QiN5VXvdZBi4dE0vl3pblHKNt3dYU9fR18LNGgx50ZzaoXR9nAc9T6kB0UyMCLMUo2ND
Qmaj9YsfE6o6Go2OkCL73u0N17jiA65wcwUrDH1Jz/ECHnhVapZ4pi5se1b4HrKeeYN/tus4rqST
bFpXlWOXCQAk/LCppY2hBwIFP1yQi/dT2sQMo/wEoHuTKa2qXzlWdk/gWj51dlkwKLz6sl/3RA2D
TLm46P0j/DxPT09ayjfOXPZRRXnV5FT+drqniiijUVDuB5Du+ZF70C3DUNZpeXmkKYkANOaX2wXR
SyGev6b6IYTr9uwXMSvZDCmRVjArIPQ+TXI/cRRLD9H3TmnaItSOMhaSqyI9ou5xJD5fnCJKKkVT
iVtjnVS8QzLSq+6avqUT7WU8S8Vb0Nu0GUp7aBNxYM1oVhUOyjsbahB5Ilc9vqUnpycdktySn8SC
hr1K6ZBInjMnWOZUnG8jZWh0CuQeBaASgJ5GlawV0bFxatK/RnFVxYJd4aikjdmvMM1Olg26eS6f
S9zSGqAkY8oToDGa7DEZ9L7CbhjPRvAzLDjuVhQDXoU+BNpm2N4qi/3Zq8Np4ZvTH1UrUfmHleke
A+ilgWdS+PFZnKWmSND2tQHgugnZdT8useGJfeAgRUQ50JkUJlfopORG8ag2naVpHqqZh+vuouO8
/D+jkK9u4ifAJKn70zcY/Yl8SSTxKa2HtNHOmfJcQjoSLvkam1Ikotq3LDmRlPD0/6K84TDCqAAo
UUWnAmvB4yZmPBjmOWGyUHsSengvnDjTfGdhyFazYOt5ygdAyWqyKSG3HmGjoWvyuXZIuor0KaBk
AFmviWax1YSD6k8m0LmBslSMgVTIjWywSrbSNhaExFwOaTYF2YlmvWa3i4IwLzIRuQEacumyZLYn
j4+ZB3j2LiWkhnf6PRHV45yDA17FNwlzxcerSnXQmbyoU5TF5G5AVxXC0HEebZCDPQrqJb2XcyhV
wtcDdlapM18lf9Tl7q7OLCNvgPxA1Llt5U1NVDiMrRdGZ47KwpRmlmKdBTNgl0Qeof/7KKii5O8R
AuB9bckAQPm9HNYvjeSxvsrY3XvZSdXavtm+WHCmjXOKa/WKhtLOw4/gSJM60iiAnBNUCawwdrCt
459PaALJidKApb+Md9rmrfXGoOMooVtU1WmSee+pRr5fhC+b+XmGjai7jviHRX1TfFWBMmLdBZdG
bZaSuCLmE2QsH/Yed5QloSNDaOTyik1wstFdo7jaanPHQq7zFLtYzpHDg3WctwgzmPzYOFQlD/fx
5g/85XWMrHqci621N+rvg0CncnJFrA6fXumAYM10OGIxU3PC830vu4wYrvU21ISEunjczvU0SyDK
tIeZH/pjaf1YpgmFb0hEOOTIep7IoZhHArydRIZSyNoFAh9nxmGnK9D1fM9Ksou4zwi2EVD72jjY
wt91o7C6uBHKBixFU7LIELPUd+Ak0qxBJxI8Qd45jlYbgCxOwC2cCaexWZJB/VyT7LNZyjJva3yZ
pRQ/g8zz6Kb3MSbO2WuVqrlMovFmcQUFk0e0Xp1kjFTKZ+B1KJ5G1Qsit51wdCarWPAPYThNXzjY
aK5Up/Y2sVp3goDutDHQUqfFHiliGcAXZzjwQ0SlMY4OlzZwNvWnqOdkJVXC1YUmQtyCJBJscTNb
jjcTDL5BxtN39G5NqKX9M74YEm6ML8WUYsCUOPOumMPv+D/YcwsTeHH/J+jo+zsc4cxzvGV93ltx
ZyQ1zvnNbKEe62soh9QWwlgdiDuGr4OmsV1QJhnQQbPEf90/tZ+CP2TSXTwO+KIRK0OmXb4WhZyz
4yxPmGGjGx03vQrrYlT/57E+UvlGR0SweYIR2XWnpOgK1c5kO4a/ou7w0Z9Rk4so3y2jgXUwBKiz
qanRN234J8bsS0vTLzoubr3NiNo+Y0LB07VU+cFd53cfnYAq1zH1yktXXjjN9Masaln4OOU8Guq1
6i2+WUDtVFrRw3kB3r2ESTwPF1wzf+KjlUthtN0Fw5dU2eRsc6JJS5oQBOEWtaJ/f24xZxibhTpo
6hmBKvqxCpJAA+x+KxEvO30BATBdlkkVxQB+XAMMGinjm2Eyns1k9G5f9NhL9w2YlmdRypT+FmM/
Jpxq+SdCWqu6jBxei7uC1c1fpiOVWWgyffbKys4XUHtUgFF9goM+FqDWhcgqIDJhDd8QRT1teFQA
GHSV4YV9SmA/6bQ6PvvfObDVMLDmuXPeSptkvBY5s5k/4l6U7JsDnyCcc82AEVqkzjOfVoSWgK2I
kzk9jsQZkFbvmrbAJj/HDLrn3HBYDRLsJSnbWAP38o3AY8zAmt0zNg8g3e2ML+JgzFrLP0Ry619V
YjP/928wM4+/uBiA5qmDjI8/2C74YxWadfwVIKEx2N2l5sBWwMjhHWYH31yKPm4nFOT5VS9muhhD
xp9bXBTM8Rv+tOed1auAHedBvMeStrMOCpnpMbpPNWpHWRet6iecMwibwV8nbi7Xi5Kvzc6yEn6l
fQ1PB0BYLGQpSimDir9OxMFFnp1EJn0USzqGOisg6seS7Dzk9sdy4G6FR4T908995NSLQhtNQOQT
Nzxfh2vNvbKTgReWmgSMbtZMwrNB1dQv0+uAhREP2BKFB+vNEEv+QGIJmWsaon9kAw0LzviKC/i6
IaZIT3onguNcLjiKRYQdL7EXl7qt0iUge93h+Z7IDMElwBcauAkXmvI0Q+iAPUklnCHF22In9cJz
aGERdvmtEnzliRJ1qvsVlFihO7i5O7Mqe4Op3gHaWExYt4y/ieyGaNbbBlf9cRMi32WmiphjWfe8
VpyfZ56OrQMWru7Q+ePyAI1Jdv+CVJEpxDd8AAXB5+t7PtuGyQ8f5OWGHo4D+QsOZmh3mPlR7nYl
8+SzQlS6MtbbEB+G84PwLmWBfBGpmuSbYHwwtgNXzWrvqIblp6Q5Qr2c7kvSXXA+LuIxJDIHexdR
DVlBgIfOVAA6SHYKv3KbeYVQ9Lqk7VdkEniMT0oVQvIWCTpigUIxGN1bf9VqGzN1Aqd3kWtj39qM
T1Y8aMa6m7S+mq91n+kHnqv0kdZpiu5c+bHbywWjaOOVFBLQ0dZVNM5y2HRREI0Ef+BVyOJ+Hemo
xva2x3uNCdPU0M8yAgVqiZuCZ3OU8Oj983acDeLquI1uUaM3QW5B/+uDAvDwOHJkALEtQQimcviM
m5CGTTMUTCN2Wk7TvZqJuDlOHvO8qvL87q7Y8grJO7+wHwUFGTJMRoFo9T3ccZHFKgGMlmfLF/wd
uDBfaSx8jHhaMp9igv4U0Z/xPQSanKk4cIGf80hg0Yv36KlxKvgQqUNXrK1GGG8xqR+TWa1tKS1T
G/UY2/cK6m+TjLjicsV5xfKgctPcNyjTXf1metlux4rk9HSoL3OhD6cFvu43L5YgcbszRagHRJ84
WGJrUVe8cEI6KkDRaE3v2F800iEl2MJlw+2oiDmGG4jD1MoYe0e8QXOzrGfY7pnoJDXOeUC5v6it
gp4zwYfFb69I8culLRRyxpGslrjec6gBUtLuRwAxxDoX2EkrE4NefJQGrcpIOwEphR0OKu4AmMjz
4nlX8pxyH0Lf0a27RKv3bLsqCfiC/Pdaq4k+aKtHzMwm+MKS28dR1UPEzd1rzHsx7HszFTgLn3oj
DdIruk0zh9qeRuVcWXepM067/rqKEhrfMcVxSPF4pd3a9Y8H/zvx+WxCDs66upjcsnpABxDi6uuN
k9kZISolpTmS3M4jksDFut0+FG/OKr8rzZx6tn1reez8MxzgEd/otVdILtAIY0UQ4dRa7ffHgloJ
lcY9hifecFdwd86zd4BOn2PbIiC11tfnY9aEWCF4G8ZsQWlznLSKrq9C9XSqD2dEcIK04MosopD3
OeO++hHbZOLq9PTpP1oqO0yigF05TTqbkJDSVDdcQfF8rQHzBiVal7VGxqeSf3FcErUYCwEuq95b
dAalMJN2L/RhXWKCURc8QXaAjf5rPqsiOb6mRpIsnlJuiU0T9otCCS88LNhIQRfqdXDJdvGE4pYf
60fVrSE9QgT0au8/OckAdYh+Xpgxzhr4S+O7/7lrXKrWJM1fVzgYNm604ENHqo/SAt7r4GyQAMl6
oZO6zOnRJd2LtLRmaVt6UAfLabHLADiZttOEYpwzfeL+S5bgiySSzBvAN5blboKJ+l4Y//k1WDwc
xMnIun35bmeedzM6zmZPN37uUvhRdpDh7VXNvDH5738in44rbASS3TqtcWOcmUwEnCSCTCj+B20r
8RL/7NfBsbwjgqtM2wdZEdWvVlc6W1bz8zeMsAc7ifjux7t5sSgwdYhcH3pELvCe+0NxJtNV7Jc0
VW5cVw/WzYxOaHzCoq+bTCCRwluAISEmtAoIM36cB8HO1n5xcp85ItfEFvUqTMbVQjj4MXfQJ7pd
nvGvrXWCgO8debYT9EnsbQzDKnL8R2QQUquk7/LTeAfVRzS3Vvs8V3wXLotR1XZzoUrKqH/IvYsV
/10WqRrUIGUuquy+tqV/JCbtrs4GdECjSu0zXe0MKrs7kZjqWfJPKKADHRSWW8GMXb9wW4jgxW8K
gqOuDDc2iEm38It+Pp1jZ0CyYkgQTh1xbzFWZjRb+stDNyU7POUX3ADo2AB0C0oa0oAnYm0W6a5q
6itFUWthWBux/XiKtvHnMuJPYjjbYoSmYcTjwFu+uwl7RJXf7KQXFBNTBPKdlqCWVMNqfFK6f92o
zX0AWOS8ybIR9fxGg6EAy3hwz7onb+RwZly9fvsctFpsUnW2CObNxl00tqK56x+CTAVc9d+viL2S
v223EAOw/12x/yhROiENPxl1+KIGwklCwesVQlnZKJ3JSAR9G6vNYzcEQJOg7l7bs4yJlvwWd18a
QE32KwFg9TucS8zD4FGYJmKX+2XULqfN0uIM44PON5MHqYpOe8Zvs8zBMsGnlv/9B3WA8McfW54M
5ppBUkMKrq8XU+m7vkAsgw4OhI0OfXspgznmJKEr0OMTH7CUMWk/WeCEAw/GMesz5yqKE7eAhhfH
0pNKGHcxvL0+RJCv59haG8slMTz0Z9nAp3UWa9/Pk1vQ0d05H5xebJNah/4GH8YO6zIeXL8XoGVT
Rxa6Q0p3HXMabeFMUummLhtH4weVibVUZJH4qbbeRv7L874Z1dckEM52ThXnUV+WeZClp3fPAzMo
jfQP9+nBKwtX0G95yDGy5kFhR4WrLqPA7N69xMCporbK1FXFzp7o1g1gQ3CgBZtZqI+uFzSTq6zu
YeB2ZRSCHFK5U1MhyAhVs/LjEGd9scWd5oD/lboYdDWMnvJzv49DZrEn07zCeeL5icYkWzciS1k/
2bE2SrijzqOgMEPMqmgULewhs/2Emusbh7GWamWUud6UrWbt9uEyOHYRNfsXRJyFosQXk3TzCVpJ
gbb2oRWP914Gf0337NYxGGWt8eumzcEY7CNVB1FxKBmpdq+PaGuRSTQcsXRgV7bWfcC+A08bSSFY
X8wyvtR4FPJrYUH02cvjaEzVbJTHcsoLD/g/l70vOzRCugrun6J2J3Ac8rbc9FpSnOUXATAqCxdx
mmlCc8eQBxH/Bot8oZNMEwQAIZA6KMZxJ8/m+LtLJlOB+bG6JZaetsRW/JB5N+0GHflF/annYDJq
iL6V32ylq5e1yARQ8Yq5pPT8l4ASffkq3+RUs+E68aY3hGJp6IjRRYqOrQn2IIzgEOXdubeH4XYe
ja7LY28lj23MBXzjCXS2DI6RxSc6M+HEZSfULKwtg7R7VmRXdVnPPGHCNhOcjqvnDSTacjEvwkYv
mVjOSqXR2Ut8wL/fo7zc4+MN8JdpISKCQ80IvsOoF3F053LDG+l5mG9Eftv8pMg5P2nfLwv96euc
ilrEbVRwfHmg9bXVqzt6B9v38prkgIiPpVZZ06Abwm8Z+xpidRNAfaVrm/WAx3PEy/1XveLlBaWC
044QIy7bcYrJecgYA4gJoin0C2ngT4vOerwQxspBjz1EJpgOMUOw4vJQol6gEXEXDqo77e9oae6M
0uA9P6gN3+7+Fcszht7eJHo4/mH0DEil0/A2grol1CToa0nswj/ccM6uQOd1tRstsKTAtqKPX1U3
Vz1SJsQX0XMqhKMa+i/DuJxwC0PXg8wtnt/5uJkKVljMGfd+TwDpuBgeKvOBSsh6vomSUiKWVvm4
SaIrGcsoWOKM7dvxPC4HNhl1bWLlN5bzrPJWuezrqAp4Z9WXlnloMxxW9UejrPiaZbq0iPFO5XBv
NUAnrhnga1J5WMQWpFWusCOdFpfkmLMDqIjYCcsdJeBx0PKzyXMLAdt0oi57P1w6Jw3XQAsaXtEC
6ctyCNfoR/FgIxiSZZJSiXP9yL47ihAq/0XjDK/mqjk/b8AKQwv0jII2ECBePtlYhRfWb8JcjWwf
KsXVle/IOZKn98GcmLs6JXJFUkz6qs7HavD/ieylUmxQvJkZsiRKq9J63WEhVIZMa/h9IJh5ud06
Ld2ehESyl00Tn72LvmBNtuNFWSCvbGOop0Lx5037zDLKWsTDvb4adJLSUAfMcmInHjn6R7Pik3yJ
lb58QsJw/Jy258IJUrsyf8aXj0NU6dH39l1IChS1pGjd56EbWXvfgTpXjUcGDQLDsZ1+kTnhz5j2
MM9k7Xz6b8gnS5TwHJss980D9r6Gbl4hdgFqrUN50B+R0MEbuqKALzKjkC+MWBub6r8586AUE8eG
I1dUN258F+3XnxtzuPbF3pp2WDtWFXCAUwoovXbaiXCetjBIRbBnqeNSyiotzDsrGeInf4CZ8ZZI
hhDNLLOt4Qdbf9e8KPcKqq/+8SFbqma9lB4WWQBDrdMlhmrSCf+esmhsH6ZU+WEY8/z/sw45OOiF
Wy+I+r0ioWJfccF9k4KdWZwUnibgZRkxFm8rPIEnEuv8oL6l22LumLoYzPpSpq0p/TMePEXxQXkk
Jj9qjh8rYnhs+uX5VfQuQISE/IhZclevWIBeii8m62oIT8X0Tu+L3u8vyUmfhWu1lwe+pJPzIdFI
IFmi66w73JhkNDnZVyJOgSUpG9lXrAgQ7s8FCmTXD88HG8ZpmhC3hIjW48VqS7vtOhPf+qg//mvr
qYYhccsZurX9hEWUDlw+op3KJpCN/zzeKBML1kngBLbX+iMh2RWdAHD7kpVHsLvcufH2UBJA5c62
NeeYYbMRdnU2gzQ3xndaalzViSoSDg+7e8d3tSxRHlL4vfUf3maf1XuFvSAmQXpd3zGVHr9gkjhU
1GxnULqD7SFhCzODknvgDmfpBDTQw0GSE5VdgUfxXddX0ERr/5NGjR4YJQL6ogB1LRFo1h2n4fSb
FuEWsMxPP52b30xG3PoPVAehe9E9SoU5DM9/9IeOO1ON76Y31kc/EFVtz1eugjig3zX5Fs5HouCv
dxzpFIMcP52aSCkoWUCRcgFRI7BGjp36FbQxv/MAh1fqRucPRUqvNaNk0tP46N441nORXpk+ue4e
PA31r+wFTZU2QIxctuXq/HmyI587waB4MYIrBg+3Vd/i3bbhNf+HR65l2gWZ2P5qCpPyTNheNTo0
l48/FI3fGGdo56oPp1iGbytMBN4o/i8NZE8IZf9BHL+VQiRY8Xgmv3epR7Yu6kLYlZwcDcQ0NZdc
b8HtxyVE6BiQy26CYU8MDOX6STmvwJYHVGKb8672uDFN0+avhIbqftiSzMLMcNuiPimTJ+enFqOv
cGCBoLCvRy7oCMsrVJ8mDZulHb7oKzU5ii4zE302ajlPG2+aB1gDoJm/69kYhYCzhS4LDvAmbmUA
g9xlNPDJrc2+Cjf/ci9Cbs3+HcfsTD2VStNENPQiXYXypmhRcNLZoFrRfKu3vKNh/yRCh/XCWSL/
DT07G6W+5LOL2ZM8mF9Ij8cygn6HquNoJ5seCuVW5DdrDw5QgKgee5rN/oSfIGPRX/zpegOdtYiE
4jJH6HWiCLNMTF21exZNLTBZDa2lw/vbl4rbWp4dOvOFKWjRjtNs6f5ILAUBSQSyiySVz9WpD8e/
00s3q1+peRaeO5vX6a2e/AyyN8/mWSFUxtFT738/TBLykbBVq98hyeNXg6bpw50s95Ir1K2V3unc
yOwrUmsHkGfzAoQHIsHXobeQA1rv5ShRL9B8gOyXAqhgWaCy9vPCOLsOo0tai3IthGjZLsUTYKln
6ynRCfOWto2Zw9wcuzp9XwLyp4bmgYDPO3ttrNzjY3ApWuu41yKVG8fc4AmzJrXErjgON3OTJDS5
/jg95BjqfjAYGkIYUUpX1x5A1nOe65OWeZcctZZSy+q5tAm0q6JgKdxh0AQUZRTA7ENaChpy9Tgd
zSw5bZOlI9W7rbFAL5XuLLVt+sDnotf+hBSF6RCusb6sTBptxNxBRcWPAbabQmP/h798Aay/zXAy
TsJQ99rKPsRSla/AKUZ0AnUsDKilN2CJe5uLTMoXZ/QnyAzC6L+AEz0elSC4vyWkqy8uMfLsn0Lc
IaPGqxK8h+8j/wxgFNBitGiHUDEgBRYglPBuBTIshwoC27TD1wec5pnZyG2Fjej02M+hCL5fIVQh
qR4ddaJYpxux4qbUcDk8noqzLVLeb3wrhlMkqYI9k0UDoBX6wLy7iwPCHq7qcQG+/2Jk1vhiYtPm
Ryud7974r2LeuwTR2VL6m1X1G3uFTyQkQp6Q6iitqyWyTcUHUY5MztGL40kJQhh/hL4aMKFKtk1n
SAGHyq44F7gMC9a3nu7yunoiCxjVmaDrEAaoCrZkdJUysvgOKtJtl/nPXAt9IjvtORm5fTd5MbGC
PqMTbIOgb0tzGNH36teqf3ROeA/aL4JLdQrTzWyKsVvBuM37KBxT0ysolY3oXoXWKv1Y81+dlBir
VciGgyS3d5g3/E4XpobpwK3rT3y3hNWBRdkndsdpjyLb5MHyuzE+x7LjdRCITPKITess1P/lthj4
MAe66h7zCvaw4TD7XsUEvQJ23NttIzUXRHybR9PVKxgP6yOOREcY4Q9wOgu1E92ZiPdWHQ61CjlU
WzCLFRWnFIlYRTHmHxAUSzTOUECdSCE47sgmZFkHSgaX7xIECGeIzYAabkA/PtMhCQfgzOJg3gD6
RHHawbUAEJyaLp0D7dWECeO/eRZdt1TuozlW1hZSfNeXSdNQbmkNe+5gDkKWtV9blUGpH9oaCafK
jn90Lf+Y1QcNEId574bx+Qn31L1DoaKiSz9K29b7ahSLoybTTYtZhUrhpgXApw9/NRNNsL8chlQe
Ioj4VAIZw5/5tSPFCEYFo1PZrLFIPE6M8Vn8OJYRRuqfNj1nSd+kEeTmbgSFwLioeitJPi/zn83I
Nu51yUsv+8CWotfadUaWwR86OBof0rFrux3pfIH4Xcrdbsa5e1TayBq+1KvGTZ7Ma9IVYDNSWHUb
Qny4AJ/4ZPXUQGIRQWrjZ/JbhF02ghtS/YRgYFTSScOnMMwfigUnAYw3PQ/jDKe48LRFl+eYFVse
k8zBFwVExTKySVrNzS8Bs0Gi5kg8X8l2DXLwd1T/CkKNbZRDaL3rwGSfeZhAXX0hEzAHO52yi8kT
nhYoV1qCDxZi3xb6DJBLFjmB6t5ACb4u55kDdA5zKXqTerWFJxgJ6DpyXNRHsUZzpoIPwg913FLG
1KlmdTAu7WlFW+ZMnKJSWt8kpVZSRtndZ2htprJ7g8iyenq20LiEU2GXES4EGZs8cmO/5k6A1Pu4
MjsbSIJWEwHYi8Is+RCEJ7Pt1j/BZEXCckIe3ZaKXkKtH5k/EPOScOWoKSZxOtLh7Z14qrGuH/qS
CbUP1JB8uyC81rpoObleo4epEWJmce1FWYrqEuWQv/dL4UDY+BWNuxG445frj6cgOXmRUr7XMrFp
J9iYUerWpw+UrTbJTXsgvGuR4BVf5ky67VEH0QIqf1fQLdR/GQzMd8+aHSkbof7hRXN3eRnmEAh0
8hdy9D4k0DPAieI1ctCVzyNO9u1fCXA032ivoWGO1x/oLH1TC7VNk6lkYB3T6z4e/ZcL+35ttqJl
9ENbWlQYPiGBTUM14KWuDrd/LJv0k8tOz0fzVG5r/0Yk7KL1bE7iqd2ZewE/jHWnc6i8X38O5+ux
D1n1KrWwI+jgw79SWZtwS1flYuAlzujXz/TckYvR6NG2E+vElavAOgz3bhGyqTf2D6gnZonCrCsI
ivMxUw87TU99DfgcGRXHx/a+tj89LaSYI6g6pCuOnLimZZm6LYD1csa/zxesPbsEbfWewgER2PaA
ObyaUBejCm8pqTCIwVG1y+39/GvWEKWwCkEibw3n3W6Y541hVfAHFdeAtbES9/DzbfHdHH5aHeI2
jr1kUxyagy1fDy5NylJoOOUoZc9yquYoukEclS10ZMEw7SPj349B/K2O+DELe+SETsIhi9p1C+/u
sV9eceRcgHhmPe89ekjo8NpuTJTl3+iIAQL5Op4jqaidQYn7u2G4IHgQr56LdefFaxKWWYfMgjTM
M3iWcoFh89iBQeekxA6zs4VwlvofBVdwOCr8rGnf646MCTX5bsu5OknXdeDPf/pPMVCyzthukEMN
mjoOXxxb8SXsyqLLdjkX2msCwqmEDXpXk3TvP8XEjTVZunjuADEAUUJjbRctgSgwVFEjxwDFiNC2
AZNdGnTQb+0Dflh89qwfyHFDUtI3UOyrfh1/qwRy3Lm424vZr8Cks28gj/XTGmww0exEG88/7wIY
Evqa9HETHLVIzvMChmA4Qezfp5ImGph8nqTOCdp0/Sf63bW+p4/r8MjJcOKjps4STkWmDVbQZ/9A
K4/yCrW7cGvy0i4iaTEvsoSZciZuvXuMqYJkS+5Q6Qpgo+8S0PWrndsL0kviqDbrAJ0Ql9BF4mIm
vak7nAp0FL9YvmWk4KND49qQcEr/EVAPTQ8MaIxT8H93hPEOVrbsoHl0ppctFdhvO/XmyGdmzcUX
ZO/CSlXm56Ir4/m3cDnJxL2qqpsEJhqPpQozSoBSEbZh6+0C8ZZFiXvRGECNcfkBVgxRGLA+ry/o
/u7aVXtKaxy5el09NHWr9lRHbeneIwGs+Wv8TJVqbkIW0FUE+wyu5Sl+a9PLZ7a9PuJthsi+jb1j
exqRvIG6c2EarrG2dgs/s5TWsC6EsgBwyRT2un/x5MM9FTS/i4Ff88IowDhM648DczWrrdi2A1s7
ZhQKgFAGdjXDuI36Z4T77UPXcL/rHaftF6BMQM0kpYcmIi+Z3hj2yCTviaTXpDSz9xJejr+YZBRA
KDHpykB7dyL8VvDqma4njUKyjSCBdX8uY3lQ1c5E2EBY6QYK8bUXM39b0JeLD+TowZpj0hox61Ex
CwiPGAsvY6KR6gI8pnRP01qNBRwak8hIZmVqxZhdIzJKCnhDRSo8baM3qq9HQYc0+DIsnoJVT38Z
z0QtaylT7443AZ9Jgk6+i+ROEafHweDFuA6skLi/zQ52HpB3XA5DEfC29cq4Xo0MqAVBwvA8Zlw9
+nUszZZoXkDehK29E+TmXcBpmDQDdaR1ypoGLBRV3YPqA53f8k1JHs+OK04Qzy3+EFdbPNJT66wt
maxbT6Z4rXFU9ZL5f+LzKj+4eZ5ra8KxEabTYjZOHSnlhn1OkPAI08ZtqXbbVug7QKBuZQ0Pu6Nv
pyyRgdD7EeOPdEbUyXfov9nRrKxKIpWSfC0ZdMzbbFKY56+gSiqqxktbXKYIxU6IrMvo/tOKTsf5
fBxICCZm5O7kkoGK+2JjEjWbAk6ttN0nZDe+BDmkrSeak58M/tR6yVnO7+wn7fsxTS4Hi1uVLuig
CSIA4ER5ScI+0AUPVT5HriQg4K0+sYK1gH/cPNeBS1m9OoSEebbeTf1NC1TJFv5SA703fEBY8Vgj
w1ilGxOpXTNlVe8I/5SCnHYokFZO2UfPL78RI/mLZNkISCiijtX4Sw/XFUoioAdxeT8IJMAj+C7P
+C4faw6kbdu9ll8qfCuNkTCOgKrWmsgfCr/yigEKBzGoMnACLAXH4TGF/vxueFR9HizPJwATn3s2
p+WZc5plgmaBrflTsWhMY3+k3ufBR8gRPw3TwhNShDativLgC4W1PhuD43Jwg5VYIYifzWrcRo0s
gYvJqnDLKPSaNaVekhoCa5PbUWcuOh815Wx1cm/ZUrXj3sdpeVUjWA/ia3XV2UMG7QBKc67iYHJG
jnJwwjSJvsYGqKSiuoPSLHMSZs7A93UHFwvvWVKuEhna1Ne+Eop0u7hY4/wyQXhugdfV0iHjNJtB
laX82wmnZgPlC9O2voGrN0viAsydSXXLugtH1XfMzdAoKYqbxdoIqJ/4Jv7ItOjx37Ao0iVrOGVN
IHARfFmfkC+9MbSawWvWcMfjFtRAlTgQcbjYidhDF/fMtVxVIeHNHSU8HoFUmopk2SPHfoPZC/mX
mYsTPFPuCX2E1eRRv/jhXMoCiC/+onIfsYf2oGYXBNY7BUAP8zDK5Q3mA2YVAjGNtRo5uGoDtKhf
lf6hoVDLUlf5hqE8lyDszEZ7VE4U7SvIFYd8vhyhWlmJeBdr5D0x62N+G4OHlnkQJ1Kqg/C7BMiO
rxy9k1FVWXBpfSqcxATEh70xlS2UyNfdjfVsSZIBMBlH4bHn8GqDjMlTXJ7HUtr/D1Lw1jV3O0LV
GjyrXxjPFU9g7Y6sv1OAMwyqoYfH17m/pCCCK01Jy/TCArnpY+XEZh5a85P8q1Uv8uQjUZfsXtIz
TamrNyycOi6pU4n76/Sfgms7AFyafyxxcfTt+yum02fI8mVaMG6BJGXqle85Kg/7D1Yn21qvNAlC
2MkbFFebG5I/y2gUnWFqnPAN/gH6LUoBkvo5wBlPO6hh7/x3mhVqHOzWUH8oxjrYoe3sfIQw8WeV
aMKvIfUXNmAxlRBi/sNBw764FQAIuCVDtS6m2O/O64bqu5pAnCnyQHJxDm4dqgaqtyeohc2tL6LM
0jWV2n3MF8Ff0oPLKZohgPitKNh1QTOtaqwBhS7kjXWL7WuzqP18zTS7dgX0oMfEkXcHnYgXYszz
n4Z/iUAyT65jsgMqkk4Q/8ojXNfVvYRIQGT5Iwcs3ujBR2jsqudTxk9YKF+gURhR4uwD+WDW/9vk
vLU63lXpnqo0CDMMBcSLoVjS1CkLuEwv9yuB/TALqVdoiso54i1J1jdNiOg7KgOdrx1vRaoW+mmu
t2IdZdiWPk0sK6ZivQaSQ4NPm3mk7u9brRZ3Ua4W3gyRvlvqxgfb/fh85jtTRxNHzC8n77sbpo8U
Q+adYUu3N6iRnl5cwxnyMh4l+2h8YRWmGfKIIY8vLFjEc08O68w44fu5ZCfPFABe7sCXMB1J1Nzp
T2GoGLRqmMqosxm2zlzRN14dQ6BJa8NB+UlOaQFSBksmCov4oTYKFZAAV0yDPVp6v6lvRvLeP+/O
2nl9e39NjsCCPCPK1omtqCFiuoEp1adkQYGm2XQCb4rTsJHlV7qYpvg0ddKJRoNxrugatkK+FrHT
FL/wa8BEe3ST3/yxl1LpRb9eUPJToRT7lPaRw4cKgLbv6/KVWB04ecjthtQXEd4Ay6Su9OWVTXsO
nEOe73u4pjI3v3ilvidgWb4NBCwLQ2jxU3aWvtEh7cT5c7qnlhPfmkilE4nkHJsGtNgOYWjYtzVU
1aX30fdwlPzwZn2TL3rKM3diMT7DCCO5MZ99OZzIbWZVeb5o5vwou8puwmAmTpOFE/TWbVBXtwjw
dkpeIhoK59MfQdBnyRpOhXO+G46a3UFdjdrprzZv75ZXklxx3OOfXqFmKGHob2GMLc53EtnB+hS3
hRveMcP9y6wpewVII7VrFwWLNothnayqwUO/RIk2RlZxXxjr9BwLVe2za8ZAPe7zkejcQ/jXBAZk
WfIrQR3U04NLqQXhlHnnpvx9sk6EoDqmaOoT5+jeaE9JaxRSrQyhjP8u+XmuyWbju3izd7OYGjXm
YF/Fcyj8aCFBk3t8dre4buwkmOLKNV3SZlMSDeW1/DP/ihPqkA3QulZtWZsQ7IkDgn+LzHSxw9tt
eooyGapUdV2d0/Vixvi6jkv7uaeYDy20jwvMEU5KCP6pZgDMRiBCYQq2mQp5TPFDEcnIHifEPZ3/
63Mb3zwH5NtR2qgeBGE4qiQ0EtEvWm/A0WcUra6kfMTbq+ni2UhPHdLYVrTe+Mg4jPU5Vlx7cGoA
Us3mwvTL0U6eYLO/RlV++Gev1KgCrrWcTrg28Czipm10bPhm/MEEnS4yN49Ic1h+PvMNdUZTVWXE
ZPUOxig1URA5naPpmXy2u74kzcbmnLqDOXdK/7eqKKdrtyHYolORVIy1YCAyge3LTXaVshXgqOW5
po659Q0I930IdYbTXREnUOWeMDRhpqXm94/kYS7F+7EkXbFmzg6M4lN3WKvxV5z30+Fg4LmttmX4
WFw+jL9qbmlm6JOASRKDgJy23MgccKEDaT+LypJ2rLyutjL7LKSm+tWKBoQpMWqDjp2vhUN+g0hf
DsUriXXSU7XmfXAs6V16quZc7C6jFugpl7j0yWl4HaKFbwVH6Arr/h5pfbvXaKqmvf2EPxs8r1uu
yBqPdwZA7NwnhOIlTVrXWR4HpmQvnjV2zEtm1fm1sZBGMcIkCem4/z9gD7Xdx2Nvvo+M2IcLmi5W
ACCPZ+i4foffN3P7V0Sww3uZaXGikg5iwzoHHRZlnB4xG3OQcGzOKGMRjvkFtGB3VG3Aws2Md+eo
RUQiKtwjjNBp5qMAu2Icy1SBAdmgaAtfDpGd7POvsfGXCeSDaInDV02DyMVqoU65c7GT012/huZ4
rhB7I/HPCO5kqGx8EHLj7P9gxdR+Sx3ktVxiSqSJ0785lALHXYsweZDUvr7hvuDhWS5OkC83b6zx
mXdLda655Yjg+eZNNKtc9D5YGxGsoy3P2jlDzRureM3ZRbZ0rZ/itbLHPm/Ifi//3tqEGjwqnawp
3CUaDG62uKRsBUzOYax5aXinZZzoTOpJX0lURXSohajES6pBfB4NvSQ8WuJVx6V56E+ZFMaEDJ5q
yAQHGYjQ2FW4cLbijrQrPS3eo8AJmVdzMLJucVjuPghAVNt7uKjrmzzrxdI8zT66MmwIvCQDyuW3
zCtzfgoFLlVCADP8yjKO6pQGI8IKQQvBbMDagbWB5XIWMoFqey2YpWHKWtYAdY+C6KoX8kF4T3u9
H8WkDNAYVjia//oBo7cPEhT5jfCBl4wCgp7ycoTqC62nAz8jv/wbggNTtdKfZ1y1p+O+YL6YKNMt
yejVrpLBS6upXj5xQLKtcjUWJXaqZzvXcJa2xale1W1dDSfYzQcDPV/E1oHBB+1CVVp9y57kgHc3
meqfImWjkljUX5QV2U+gtixZ0vhMyXtvtd03He/u96NEBCyNWzal6SPE+18g+jLbM5Rwt6XheC3H
2HVjtdqfMQR2hPTQXmkuJezWrb4u3HvBoJojwqbY2J2cn3MVw3bod7BNIx5LBA1BexxPfCPugG9W
djlI9/fcOPLuo1fuiIGfRPTFE/vW/Ro4bbGbgk6s3ih85pAFfh3u8UjJPYMq6wCPe3onnSAnuuHf
L2kJBy4YemgVPXD77dM3jGlg/yFV+WmCJdyOYbuiY3HpNKFbina+Dvu9e1Ejpqn7W7oOba3Px01N
Z8HJy0h1htaQO4kpzW+VfvcGh0TUrZXP4Oyf6tdnnp0oTPY6h5N0+VGkai6z1ufDcDUMiWGTykXu
RUFqaffP3PZm4JDrtPGVQ+bEdmKcJwLlrF0FsUzwjxxSFl9G8F9yu54fgqusevyMxSboi7iNCyKy
I12FDmknHOCD9RLbtPrbUzzTp+ZD+lPHlYymyeWuauDUWzkuYum4bgoG6HXTMO9IGVZN7QOg4sXO
w5PJbw0KDJraZmP8aPBi81ukWrQ988/Ou2oLwLV37FyCqn8lP5Tt0AaKk7GRLoi8GW93GBf6zuY4
T4/raQp2LbhdR3QHAE3P848EusXScbU1nI2Ae1bkiBPcxSxRmVcRx3o4w0lz3QgCP3Ba5YD8dzLb
H/DPI/aZWHHedYxi2nYP74ts4+PbJRoQYDCZsNpVo8hI99tufeiT4g+dNzZTvkU6e1ZYVMpVj5Pi
RzrCSOwuG2i29TjuzML3EBPIEWzqWiUS5w+ateJlfd/vSA7shNQi49ZIDqiyIeWHEtodYVnZtn41
ye6BSO4UUH5E2JMQUuyGcwauv7Nl+RsqylriM7gAYhM+hKvdg25ZY+cTjuZilILhqkdfcDL+PCAU
x0zZETiLwkTryes22suf5aeQ57vvd/t7vvd3adSCrTt7JdxKG72lgprqcqsdhQcCOssC4p3omdix
t25yhWHWWGvtkBVBB7FKoMNkXAnHf6ll51byC7O0Lm4MyWKckSeLf40umb+Dz3a0fsaiUR8FCMoL
UNHnXte9wykA2qso/JkSzh9SocYyUaU3Z6zPAcdSZeVcPPYk7ggYYB0law8PNXy1BL7gg9twXxBP
pwKJQggNCPLO9mKQgulyqIbJvGkSlsLdVvTNXfX6ibNGujLyMUTFomtXOkLhsMMZ8VdvE2XITF4W
4Bg5fIIn6oAlso0/zCq8aERvddUfKSxtJLT3r/PUhEyOYRF6GuqVkFjfrMuAw4KExOh0NhOdWsOb
7zgUTUKMJjMUTwSAhKXFCKC+JebnM1nXrlQbT/tvpmuJt2DECWz9Te6Mr3Pj4Ao4wRYspVco7Yno
22BR1TGlFAtOhchqzZZqh+jsP3l9dhV8bm3JvggzxiFqZ3XKOTmUtPB/5EtE8JWzwc0wfTWjwvAc
RDpFY7NSjy1y/hUm2K29lIPjFQtcFrD0zf7ihSTlwx4yLXYeWHyZn58NN3oSjUYmJlOBrXRO/v0P
+sCbCC4LijL8KMGpi/i4RzydU32cyc+At8Z5rbaQpsOA+Y4igEp9lbH20JVfrHe0qJQncZ2wdlxs
sXiNnUVT/vjgV6/TnBwpwYjDO3IB2IcvGsozznMTJlhInFgGW0tb3nqVNgEsDi9v2wxTCR9d3r6p
n6x1WHw/eTjfr5vF7xaV3+l41foXVAhMthcrwG/06rICaNgXzX355IMfdlwIrLAE8HK1SL0oEWmz
qr0fSFig15vdms3N0zfyVQZ0iV5/dWd6Sgi+uJPN4GjYjJbxOC/OL4yi+O3ecMEGUSNouXn9Nf+z
Y0gUrWWPENJive6A3tDE23/dPpLBCx35lbMfE5lt330rg9jEjAFvcyhRyJuwYmCtYiTs7K1uo/SQ
IRYbPclGjN1Xn0TjrEAruOGO0YO4WDmIogFdQygl5pgKBO5mR+b4Qm/miOH7fzeAYRljwdjgt/Xc
BgcLlMy3mclhmB+Js8WwXld8tCJLJCTgrP8SO3tljf15qck4lGv22vCMNkEoikwMmRwNRzG192P3
ZLCL/oJe5+/fFAqpdFaiDWpFvXXcMQXcqGE5smVluxPI5cM8d+GwF+yx/77aofdQ2zcQF+Mm5wYv
1chCBjVwNYyeO0LvwY/lg0x+Tt16ZtCTEbPZAU18V17pAp88OyCmHOnLeRx2SuvMUjKH8TTMI4fV
BJ5waAeJia8C/OpANLgSG9WChBoxWzHN3HLsT9l+EZcInGcvxeiLT+4iPIDdyGXTvEomMyjR4tDx
Mq3lAe3N8LbJexGm5TDNepd4JEFVSs0mMJpzzlqMcLsmd+WiajlVKmcX0N3rCcyY2ULSFX/nDRjU
grnYGz2vwY1iiTZj+VjWdH/bCHG5yKl1vbW8rocb8dPGIsCgAXOboWOcfqDn8giRPcIewuHrw3OB
74/1fPpEQS0+bPYQG2jUM5SfPqTQf+q5D1NMnaH+ySN6lhvSD0Bdb3NdXFBphDJnZ7/D8fVEtcAZ
KrWOliHYSpn6MObm0aWGIK4DlNxxnvFf+GJGFYzszoySYkvSNiWwBjbUfFLQptd/7aecqFAsO7KD
LilXCq6MRIccyo4LdAR6gsWkNXuQ6IVf3BsltTSE7IGAMNHYWuRTwakBdXDn1gRQX4m7t9TkAK/c
K48luPWcz3zRbtxQq3frUKo1krB8yuQ0PIvpCiHq+CLgo4VvXmaHRhutOMmnzMf9In7PKOBigPm+
D9zj5Ek4nwX9h6W57QjJS/Se/C0zTG00ex+CDB9kZtymzQY07Z2O2EJ1KEpinnsCE6l5itbu/1XD
FNVMYUQNcSjw9druaMPuRerW8+ssEJBbWW7rYNrtxDNz6t+GYwYoJ1pNlNUxQxmpgkEETGDDQgPw
J0l4UQsgUttIDQ3WGcNRHu01EeCDeWCn/TZ02cYyJmeaGZXugNEqVDqyTMG04Un3K/fBnUeU+aI9
JrOaTp3eHkXd9lXwVe+VsCykiYdTtXzrh9Xkbdj0LsLqiOP9xa29RhdMynkSBzNYk/ZFmpzVZWXW
52oeEm2xjnCYqvVFjO9p4SF0mFfHAksvVMECNxlN5NCr/M/vaZV6N+LUvWcro0lMF7/dyqdhsV11
8q9BpMFOcGkYHAVjv61ZJX3B3KsRgYnMVBYfJ7Kt8I8NaFurNivGu4H+J3u6ofPxqe/3S5x1yljZ
NnWZEsM22yNI4hwWUAmpJL3MRL8ESxyBr1c1zIGnIFxXLzFpyTyTgSWZELKf/fRuvjdUaIXTHZJB
UE8O3vDwenijxiCapXmAueKdTy+MAcGqSBrfS4QmU7qZpDjHfj7ZCwIVCeYPlMw1XprvA11Uvq4y
yNlvN8PKga5M21CRCimf28c4cI+LEYkzDeGSt9+WYI7JlQSsG9JlX3c/wML9CKPyZe9F1NcKBfzE
TSfuYYOCQuUlCor9mYDuVX3loWN3jbDP/yFAdoRLRNTxuH/+pD6dgAcpjHefx17ZBzT2tu/wX8Zf
9ddHeZooGsyLqAMkdS5TInB8hPeI/tzBtEtVW+CBNH5mJUwWe4+fVKVv++LX8hNQkCHT0E9Q+dCk
QivcHhJgMEUffv2qCUhhKz1Sv9VK0Gv+Jvk8WV500BwkGyyv/wnRHX6v+O++WJfqxjAur9bToXDh
NrJDOIJJwm0ow2Fco/Na8AYAxQmlT9E7mz3vaRCQU7I0YwWR7+fm9JXMg/EFKQUQfAO4GKOd8IQS
Xfh2SppA+KbuMD+wbZU5xFYZGntGzedRupZdu17o7y1tzuNSSxXf0R++6T6qpcwxPRpYoVJvBbZy
LxS9I36NdXGasb3dZtGWa0LCtjk2i+Z5AATjlp46AJa/ZtHwEPE1XNe2iUqSsaJL73hi+r6c3gev
CttQSeX4oMU1D8Zb/F9MtY2AIZYfT9q2rLk4WiUR5qebbOND/iJaSUE/NoBUiHTUMTZaMJRS4grr
5zKCLziGrCQ9lPBU4BSC3JYkhP1XILfsgSy9orRXfLKVthMUoeAYKrq8yIWAfKOfVwPcGNt7hpPQ
SutqvR0W9HqzjGL1oJ/f9/JpdGdzzT92aT/6gGotBWhp3TP0+vGUmm0uKZ38DHLZiRnJM8NFI8hO
ZOIKKdtnxN8pjkvLIlA5vzA7viZ8EINpA3PZT/xKqkhfqQJRp9krFtAOQuVZFpnG5ZjDwEoMbF2j
Sjrs1r4UkuwhQBeHqS+FUSprGXd+5eFAfLvhiKWk9ubjA4kYq1aNntTWU2o8z1lFP7J3TL1oukPt
ZgPnXVj7GwA2aHVfKpAJzspfOI3S7fqZtg2P10+nyno2UEbpWp0Z2ar+7yHi1KUl62fufNn5dRiC
D1xvkFXdovLl2llsz90dyQxJhRpqXKs4fslhjuy/km6P1svvaVbzr1CCWHe9xx15oXEq/VpQQt/4
JVck0vsVMLyDlDn8AQdVg1+bGgcWXQY4SbvqXyL79cg9PLh1YKr+6Z1zFCNYBp11REL8WgoEkKQr
SOcag9zFlIIoNirSqRCo9pk2sK3/p3IbWNY5u54BHTvHxO030TpZTAMCeLWCUJ9tPu/Rr9SDInLL
zTp8iIhWAvc7clHzAC7TBgPlPootqBxo4h5ptfi37+psoJB6xZOROI5h8z2vRwf7IgAYOliPu9wA
8i6godTCqTJ9Pl6KV4TAuEvCxXCmM5mA208Fvkg7nMRo/8Y9NUGJ8BUU9gvsrZ6Zri8Y/WkzgiCf
sieZX078mS9c8rmAB02olQ7a8DiMFEnAaI9gnzhgHUc+LdHkEeMFryh/GwvRjK2NNugCjns4FStC
kTksoUpekWCrqmdnR/LwizC3sx5nHDmPINhyZOwbGv4cYEQIqknYNsc43YUbMPPwMV0WwB1QtJKl
l2SPV331f5Hk70mC7qeyFXUMZwtBGNTVQkd/IWygWFWZDJxOC4hKUsJ4ffGA7mXyD06hzLM6ynEA
smxCSYpHev/mBbDKEEaGChdPy14tNdrvlkCDxYf+wOch6lDof0mY6bX6WI4oz3OhnXG4/kNBhfaF
0d8hzOxc/oSDpbhbmRycoincLkW++jHXSR9WCMUSWp0s3EFqT2TayTIgLvX5yx8RxyHZ/Dzr/mqk
jHbvBzIH60H/K9oMV1J6P0uFW32eB2jYY2nW3HbsrHYE/p2t+lDJDkC8wYMF7PAxZmWZQFDn4Y+8
v+b4XlBVscBovxBR5kSWwjI4wUPbmvQ2KsNRlvdiGR69BRwaJ6SJT7+nJDeumCRcvH1w8J5yHE1t
ONoUS+jMwfySBKtD1uXs+XJEsYYfpAY1zVA60HK0if/gC7+25RDjn2WLU0HD0v/CfkVuuXYwBTj9
/nCbBF7qAhK/gmTY3RYXlY2fuPlxAXNTZI7x96Lzvrk/LbRJIIrSKcg0BpiuNp6GT6c0SBuY/Vfx
1szTteBe3icZE3s5535pn3c2ozW5Z1W6yCPFaNiXHY5yitZr1QFIIly4rAjXOqFQFCt3GH1K69aZ
reugi6JeLxmmvH1NvHyywL0IYK5KgqobBl3ewx5kKO/+lMOI+lQf7tnr5rE9yZp0PWxnwuMglZOD
cbp9e2LG7TOizmXQy5A7tz3PAgfgvLqn4iT/62cNWh798SbQn8ym/CWazOxRxBQgeGHHCG/dzqWT
eo0cLMJYME3vHWnhAYTAWDTaIRUZrLXH9k5mOvcKRdCPzRRP3Ic5J9DeR+tsbbTYYDjSLBDfdwqC
LvmZLM57yCmrzcqTzkpL6bMdsb9QO0A8sEuFveecOAEkJEVz52lzioSS5o3mmZP9YEYByx16jnci
lJMBVDRZr4w2rAjHxF5wuukfhYRx9G4+Z7pxzBGFfGHBPGDSLmPVOd2XceARxwxEpkabZ8eQzvsS
Jo7M+Mw5lZ9GLa+Ns+8F0FR4xnvWN67QKXp/us/BquRmNwNL8xZfTlS+cQKUWnLB2fqNYKSM1Fm7
ptlwWwp25Lncyb2o6G2WyNhHsFBvkuNPB7mwq4OCwaf9IeHFn21h6Wb9nrnv/JJRKINoa8xoSU2x
qEqp2yZ509C+Z7ZCukKmfqKgm/BRNiv6cOWYyJiJbFJqoeqtju+ShvkS6TwXs/bbrNYrEKbUtjDx
oZ2CVsM985ip3EP1TPGiu7dNS3oPvHm/vtQWgjvYbirD/mABqd9bz8Xvj8xyXDH/r582WM4+KfN6
NVdKUgKX5imo4PDhj5IjOTrlREbKZBbAsJyIct1nw7x7K1XVheCT62hbwSLuZeDVevkiYFC7kL/S
1HCGIl1qKDlGbDomh8tTRrxxuSBHeCyC+V6v0h91EH5NNOcv2kVBiTjs0jdhDc55zT+VSor+JwGg
vv+GHy3qQSFABTlGcxN06twpETShI/aDvKWtYPPA+SzfSip8br5KdqxuVL9XpoPoqCT3xiBTGVyr
92Kqk+tuNr+MUqEcbzSZ4LbTSUpIL/ul+CRWBaA6WY5tYSYazm+uKYxnfKXS0GnLy6TORIvLXUBk
TaroIVEUSdsizFEJttBvnNBJZsfOOCcMga10EJPBi8+fhn4c/LNOzj9E/8rmsCC7CGqRPSkVhQDp
twmTqBXlZYMfG/YDB2hLpzCZlQyxmQUD8U7OykyqQaD3ZG8ENr+ePzSrAVs7MIC3iLoZxs8GAQAt
SnrRil5TjlMtSgfBfXjamjlLdtoAPgKX8MbIRtYfdVwyz9LI6NeXevCMmeP5k5i4x+yAlSOdFtVR
eBjVmMOYtQU5uZAD88l4DPzz9rNgvMwKXLvqy7zS2tndWbVexQIS3nyW3DS6iuUcBIJo0aVMfr/w
vdFBP1R1/fZRUIAfNen5QK/9QxF59YsTqZAinq1dFEdoXTdGgsLf8zfQmQkgYw6BjmgkN10085wD
/Eeh42Y2R7jvWq4ShEHHX+9Ighwx6t+BylNmPt2DkLrdlmR3rM1zSjtvX3PEuNl53rkc5dBKE77W
I+eR2wUth6QML/46uPKk7MeQrrKSNOhMLtm1Jlc9S849XdNjyhciisybLmpKbcS2CN0THgAgKw57
EdnO3wsCehFjzDwU0MyJrNqUZXYQr+p+cTlMyI6olYFSwo8J5nRt4P1YXJQkH/VnNYfBSOQK81+O
xLAqe2bSm+G0UAFIhnN/u7Wg5gMafyCVyCll/aRPEhVivq8LFipI2jG1tDX7oyiV2K3f3OKPPXu2
o4upxP1IXFQX7hzIcHk33GCIL5NfhMHX2IiYhP9cffokD050+2zOUg6lAVeRygsY95owujSl58CC
zPd9/HEqqv7sDUryM0fJAO6yMEn9i7MEvImzBJDgUsWG9roW2MOdsT4QGuHo0igWv5a/XoR3QOnQ
lt50LouLVIblrkmXHiIeFxv1SkiBYowxTvruqE8+Vr9zVeTCigplmQFid0gE5q7jyZi/8cKSvOKx
/aai8diJAA0y5hhq0tRYARxq6oiT86gZPgm9elFJodYLzKiSV/59hVa9NKzIyXMs+23+uV+ZaEwL
QEdVFnZQlbejW6KEhyKyLBfiVuOqrCy9ELuZISnYO+3O5ar+Kjcj1rpY8zO2sAWWaIP7YZ8gP54a
Ksx8o7ZelTFzziw7IP9ljNz5BU/62P23nxLspNfJS2Z2Gj8/gTaIUGxUbcSgTPiU7o33ZO7iwRUZ
x0qTw1YUGlKbxXyFVAEU5NOFiu9KRvgX1cmKZYOkzJhgAEId53VxhUaq+HrpOsXS0gWKztMV9/jI
u7dDw5vKjyiw4a2hr+710ZKQQvbcLu2VBInXrzMPXQkx9AjGyeXEYNyOZCtG+OZoHYYgRuna0Vgv
ZdyV7ihGHA62OPRROo3L5mkRatP0KuIqR2wJFTz74dgMJJTxzYfK5wByphbh3wLUJa+zqKe1DdKY
KEhjRhTiQ7b18njhG+qQaFpnCp+1I3yNsKRyqMFr/hAJpmxei/vtIyIXF5PVjaRglGd9exXog11g
aNzEm+J/+cv1aZENnoLs1QtMgDNm2gIqxva5O7TGTR8xl/fxEdj7te1yMp5voCd6vqaIVNIlVhdN
gU4sXErBmZLl+ZSbnxzLy8/dOSdj+aFO9BjcvRKcWnOk4Zroa1aMEXR6DlPKGyQSHm+FHP/ePStE
XP9gdcCAaabfIacEeK4/2LKGufIu7oGzb259v1yhSKBMJiL+O1QP/mO5FrOWa0h5pPVr7NZw0zVF
LLQBO6BV4JVKZJ59T+ViHDZD8zkgbce1Tws76VpjwgOLKC20We0f6GsWoeJ7g1qYQSHd78T6S+hD
p9e9UOprz1vrTlmRzYgu66ercx0z8AHDCT6Y0SKuu3/RxnAKWyWcCAKdyrL0d7bX1O/aWTF6GwT6
wtKT0lYJTwYhjfB6Y/+Y2+2q6NcZUCxBGzcB7I9Niclz8U6Nx3IFT0yy4LvQ0oKCQTfP8PFQ7ewx
GqgQz/wbITSBIqKOVOON/LsCFJrjh0nm3qCDUtj66+ivB8MZZ2ohjylFm/pAFtiqTyO1rxK3q/qU
E3uhnyz9i+zt/NquV688qcoaxbnjrdRmoM9cwx4CuD11PDVlJuKOy5dQ4BhVZvGqX9B2uYTLn8+q
fpOvqwRZdPpoRdXJFH1s++l842wBc50EZHHK4PL/YhgBXxxJPvQLDhO+8/X3t/4y8mrwyIM6FhMI
d0kJTFZARq+pUkHO5egWd3g2HZ3THvE5PgJWILDzujFszcqHqFVMUAPAJavGHPPvrF0NVj2scuRC
MaJQrbCf49cPTTxqqh0UBByz4EdX07hmOeBZ7KWewVySf5EYS+Hmo0kgrUjfwIxfpOB/F+CPfLB2
xOnefIXKJZ8aEM9CLnN15dU8Yjpg7r2rooEi/o2XHtoqZen1WqCHk24IHKvOIXtP1/DGMc3279hf
bHptJ61eoEhoNSGYHjYoxigYvZ3eJzKY27vN/KGdS7is03+NfKDXxaBcacPpStiuYBsgGsGxpIKR
g+0gQf7mEeFzy4zJFwT+0ACeDxoRK0ILKJQ2MWJAv6kK9a7VCwgdaxhtNJZloOqDdwJQDBw62ANA
Gta9EWBbwM8rvfKxTXS4Px2tcuA6usyOrWRJ5kUzcm4yhb+bv23jT2q89h4DoopginVIDgMLT9DP
BcdjwfREcdq5jkFsFYRzC/r/VTaXCtZCkHewEAju2STtu7o1wR1GThMHRyhmwXAoBEcUHDmlAQZY
YtEZA4SfD7i1hoT+/GPubnO81ek26Ez6kZf3ezicrWxix0uC02n8JW8xFysR77+qhXB77L2QZtq4
cFNivTQzEeyUqHrADrE+//mZn5vW7fUPEz4ZIp+OhRdAfIt7zZ2rgPLEkzj5bu/CfTdEKf9jNSol
vC3MI1duKNcNzV8GkTipqBrvYQet6w9Yjw8VIdkLyKJWAo8aJS3vvVUJr3AWwYty+IIuWWUK+ErT
gOD41+9U/8nJSF4iOVQaBm9rKOdlLqZ0qknT7rjpkxzV23je+lJ5WaX5bnie0DPoBvIKRzUVAKU6
g1d2D0qkMTF582wC+oxy/+WqM8H8UZzttIiPT3FjVIvHOgh5/kBtZjeJbfxbZroWZTlSPCcraOiS
MXUBn3j4H+YOPQs5cWsXV75t1mTNlYOSAZ3HXzksuSlumSXqlDISmpXo1vKXNa7LWJEun/yKNC9/
vic4myR6FkIA/9GEFb7uj3AsfVsVCiH6zrlq9WL5Q0fD+9m6CruUWOAyvodg5kQIBDpvqbRUFB47
jVk4+oeOqOjTM+WKYoN2w20u3+jCp72p6z7q5JxK+N0fD8dsSwl1AfRdGnQ/qWZaneymATQaTJiQ
EN12xj3Onx/+frwFse+iL0NXdyNXbmeuhzvu/fcn6BHDXaz+KmRICJgZgHDmvSmmo85I1Cul2Ohm
xj+UbDa5St5rPsRIQxsGOZ5o6DOzWflFjGHPFiij9wevV5AO4vTTYpiHgXpy0m76aMR/C7hi3PQT
mB0R0SO4YfX8R7EO1wrcX7PxgjN3YWCJKEK3SeCNvOlVS31MOLFszFDv0m6Qq+8y8IWUvBFCRzHZ
Uwdol6SSWGDaK0P72KO2OfdFu9pKmNOYYznOsuLrBQGALVyzdNd4pu4Anet9J3SjIutcY77bV0x5
SjvpY0xgf4Y04XipddXVVRc4FugD9y4USqdXPY0ePLa633/z60T9+Nisxco3c3kaUWDG0x2fXYYh
pLUsnBGDt3kkPQVCkkhyjQzoLtWDE3PVKQTn3MpKzA4L6TFjR3/Nvi2Jczhkb/lqb2U5cVnk3WvJ
4VCa7OB/+AcKEQgkefDP9e0k7zZFZRnkJmNwPwN49vH1YVRrkxKgiTXHNAWXwzx6dpZGwV3Md1YS
mLMK3F16L3dPeukhulR2neO6Lmye9hiuz5IkTUh0fZA/+QtG+5wh6vn+anO+sxU97LeG4pISZ8Yk
ggASzrEmHb47WVJ/sT9Pa/qvIX+6ls4Bx4bQnKXxsfRxzU7ZPBCW4/hBrJTuol+12J6sSh/UreD8
Wb3TznfP3eubSH3IiOLJZs8PGGCSrMEXdZaBjSfM9yWuQiteoErkZwKuPpzm5Wdrw6j2jNLzgjE6
U/ggNG0a4zIYqTMUOSSYcpemVUeTohNhXw1wnESxGIFZL2d1G8wv4pc2cn6aQlp9LhFZJEX9Rdc8
fhjccHrNjY1h88j2ReijYuYgWS1VhmBy/q2F1GVoLZLD/GvHb2b1j/lAs2h4067Qq/NvRuw9BaxK
n59mazNBQpiaN6G1aZxdQO00zIjgxKNOSekq2FhK1L9oFvXRnZlYVNsIHbZUJzxkYoSAbLV7QxxB
bF9um3GQasEitYu3V8OISCahihC1klWcTH3/QAVP9Rs4V8DZlWtA/OakbMVA0zDWRHGujN7kRRBo
WOog6OSUzmVT3Vxs5JIdzUSDu0gLeewRDdUayZoEVWifBjwUjYLb2BMxhkwK0TENvSQuDnqvTDjB
LnFL/ZjZlnJkrIWCPQh0ySIpfSMucNtjJdFFr2udf5qiSTrK9Tk9KrQ05/Y8J1Fagsp6TD5sKta2
gYBKAEB/YzY0SHynu15yBBvdGJQUkGxeuqBW+M5zM8DumgLuofcNLfXhcBU1Uli9eNzTNpgBQlA1
/A6o3nDLib86VoMAsvun6iGJQcxiG55R8eZfALL721m9AnR74uzCI/bb5liyRP2cyiG6ZbSX3m4x
ymg6BtdStGUSaNSinTOUF7nY+4Q1pQdVqRk35vNggZLKO0OvoGdwE4RNkSj+a/G9HX8c5R1znHkA
fNOGjrGOY6+3y1bhtXHTs7qWSJ1RjYqm6+y95xLDMbWu2isxw7a49cofOsNRP6qBvKbkIqonpgCr
pdtn3M80Gmg6QVORPnlSShobTG/C+X5GxCdMV8BoC6PCIzRxqjeqdT01Pe5XBXJaNC0OD26tgUR4
odTNq6ucl2EtWKKYxYtC/ZtAXrB7FZfYYI9DMydnykdItOBIYEPrfkOoS+fJhjE+Ir9jwyvwUhMA
i+ayvqwPdz+wH0FCbkmiS8o+4dR4PqFMWvRDp0g7n9osxhhoDl5vLh+loVUksYibU2RTPeN6JKYJ
xG/KnTh52iubj848EuElByzgwzRp8MDOVlyuq+ZA42O7YxIcCTWzdjEHPeLVy1lezkquqtpIY8yN
TPrmgl0BYeSbBs8O24JsN3xBzFxAXSrQ1o743o5bbrzu42xYpWGTYjDs6fGpC1rmYMi9WolCLUhz
NKpqB8JLBXOe3g/aVMuuxrZoFz4LWN/vIc5S1IvfZgABMOZPa+v18eed8Des30nbL4W3uZl7i0s1
iIi3kkXsIa+541aaYNBEgc/LC3QryCyCWFPVCOH4bNdogo5Wu1e1O45kjAx0Iq4OKS0SHk0KYCJS
vjtefjJN7BOCF5HHWTDQ0mYgGcUv/SDHO1hWLR1mw7HZscu6KOg5Ha2fuYXTjdowJmV0mBRxdt3g
cU+CFV7Ieh4IiZkjQ/xV1z/doh6A87QGP3sEdKrpqMIuFR4hAc07uiJKL4OomXGOOAlUZzuuCLVv
0o4fszRf7Dyd6lwTZvn7wBi1nR+B7K1wvLQbx/ZSAW2CfRtHBAnffuAWoxkFwMuPfj/84kSy96sB
UcBfiZc8kklOcTJJTjE0/Jp8oHFqLjL9C3P4wyf6oMFfLDykw1Mi//pnZVirZscMOvcX0RYIVBZ0
IwWODogUC6RmQt0N6C5qENRNaqzff71hqkLyaZ1t+2mYGKo/BucGwg+jqlKGfCk1IuxB50Y9Hg5Q
ECXE4qBYou621pG3aE9D2om5vZLv+sGY+NXElHSHduPjMe5qbV+LfsvU+s3pJvXtDnrmd3RSlOSq
xjPD1ipKNLbAvEJeKNag1LluFC7NI6JaDYIGaG90df/eosNKV6RfytuJoUhit+0EpcE460vZBVb/
Gx3B9yZKJ7XeOp6aOuxr03YUK+fHlHS6q9oDOjEWloJs21VBwaGuzvIoti0+DHj63WGkeHW+U/xs
hcm7gMGsJGpDBWkuSrI/X1E4B71XJ9nXLiuSOpgX2zxmYnUhtvigNL+HBQkjWR1HO48lxjqKk/29
4SZQd9qwUh+YLXpvYcqGcMSE8AYL5yjfyuUmoMftwwiM5s1SbqNTC4wrP2dhIzddd2OaWRrGzMiG
n9cC4giLvxiU67hEez83bQv39tuPf9MobQLpaS1Vzy8kQ516MuwnaD0gVESvWYPYZwvjVz1DjFPB
KTJDClfVPZ2uFcYNBHWaBF55sfNFNH1xaw23/ku3x7GYYMdIBns/hwDhTWhyhyI5/STyIKHK1oUv
GF4JcC0DuEjg9sKqKaf7abf9NchYQ8ZrSx1BZ5JDjVdrjwl6tW+kmjhU6xLoNwIMvjktJKPcXsE1
AOIWQYiRdYSK6MdZ5rpgsJzgOpyclIcvXqGWzT/bdrUTA8kat3lZR2uX0BrvlzqQkPmeG4jHGDQf
hs490OSiwx/uIpATzchBI9BNhPXErN0VMCHWMsy9PivuTrE5RFXewxLEtliINPeCsW6uZIBS5Fyo
f0MDWOaL1oZl1z4xhirJeOWc26GHCqgyRI/xkzIyV1sCzYFJrArYooA3PWqdCCRFOoALxgBGDSaN
CwHclIxZyYtCfhx1hZOD/YZXrbn3GUDGFwpx4j61wf0SxVCft46y1wygjKETBm2jZZYNCtzvnaMv
H05D6n7egd1G8n75WkUJ/3mJGrT5/c0y5cdULlpu+WZ2IjZbgxSdkzlUz1k1FCQsef/aFFQCX7aU
9msIhAetaTlyoAkDtOE9ISSSMSybzP/jhscWptTrESFlvE/OqtVcY73ar2tsr14HgVbO6CBeGyKx
kKVBcexIV8veVSjkxxVueRTZXUWs16DHir2MV3T/bcnR0LIjFZ5tpwZRu4E38iNeJ+9EmVp7b91Y
vVgwpdUbYo8M+HnAPiB/AsrFxhQxe+cIVg4rYCruhfW3bsg+FHC0EnrOAeTEKgRspoiE3DL30kRz
4FU4wTM7lDlyXtUt4CyKKLBmUfrmmUR/ITfihJ5yDDZXDimwNQopV0IQ3icS50ff55KYyVHCXiKj
w+UXo/IzdQwqypXSCeG81a3XDtTU+Xw+GaXmZnZaaAIyPppJq2uCCH2oBxgkppe1YEyFq64GCqWa
LdsO2frADwFFTzl8S1TGPdn7dR7deOnnxHE3ZgromPbQDoS/rjoUoeAPrAOj4vUaN5zpWxD4XL0i
kYN9Pu3u9rWrDATChVoWjx9jm3HwmYwROi9TFDkPDjn9fFR3DeUopXb4NsiM59AeAc6rM+w8BDtA
rW2op37l/OyB7rq/Z0lWtCS87YDCvqCGcKEmdVt1o48Qo9wwMHkn/gcf2yYtl/0Qs2OLyA81ulDM
b93NYLnB3Fb9EmvhZZSoRQGfoGVGh4mCeN2qC/cw1fjNnLL1m5egjfZtWC2W9a/sDzbPt4N4fRPL
hZ25z7QsMo4klcxomND66BiieTMRvBWXfGEOJqzGNsumMSL+xOg6XfoYWkxlgntSukRCSCv8IVnJ
hEyGRwKcgIivOYoBbjsaXAdVxZyZGmQhhrtCNOJuTuOZiWPg1zW4ilxUZjBwV5kGpBrb8+Snr4z3
KCaAS/hLhCLHTVNF/BCXqqHsy0kgrghi2K68FdlGhmZh8nTp1GcKJREKvk8zI0Q0Vu/cnjOEapyA
GgbYQq5+2UT76TsMPAgEJaWIcvvWeUilYPGKbol07DZE+aimpWHOgXz8x2oa+7SfV3V8S88lMdFa
R7H0jXvcftVG1Th6+XlkIIP3+TrcbXTuqKbzJs+C+VEWbzZgHBS3Z9eANEqOIM+Q1/EN46xH1ZCS
RcttUEDzF8Hx1MJdfTft/BWwlRzpinigB7NwHxIbxcvKTfaQ6Yk5TUIH8giVXniKVvUhzk4JDoiS
ECcAgD1LT0OMrP6RZ4PwXogHvTtR2LsjHlYx9066zdvdbNtqKWY1SAp0kxCc+jSpGZUaDVxbm0gl
U3UU4Irwpej31WNt6/ambdaZMWpeBER+eA7vXf9J2OCYM1xcxzXD0w6d2SUK2UXuOx3e0uogVySL
zjP6eB3bQ6XyjyHikVV0/VStDm587LlWx6C5pnLpOUUYO/cQBHQ+DYt6umSwsgpk14qjKWtsMYTA
z/ue4nWWHdhh0wjEAqswbqa2lPF+OpAJb2wr5ect8LPWS6ul5JbH0j46+Sfzn/UUmQNnmn/thBW6
pU4ZFQkQjYu6nCZQigj6aUpU4IFop3k1n9/GSWmHpbHJtg887bYuh83l9ojzMaw/le/s3ptSEka5
hC9moSJdKky4+qvPVHFU0AMyd9Dta6H7ZyaHXi2y8Y8iw4hO5mx2Bd854UlT1HHmEvEsPDFLovLT
Ob14RGQjW+No/AVLJneJelSuKEQu5Q3m9bhKXP8U1+J30orWc2sQfdPFZs9gDE7HGsfoQInmZweQ
DKeucBEkSYk9URLbsLENg8CQXzLLKQ3ECzcNKk6j5VJkM3N++f0A3geRnsDY78u4FeH0ULbVIfZu
kuAHWj9AmiGL8HQpfQepOAxJo0ICLYQLqn1duiiUhjVjHAoz3poZUYqFZNlga4x7+79MYUjRwPsk
FT0+9VxGZw6VJsmpoq7kHr96d8fx0eznBALZBgJ425FfYFMIFZqdRIYKFVLxTAoH/HtjjfmewyQp
z3q1YUVReRDpAoajO4/gyQfPAk3sesuvcqdhcLTEFlBckeMhsE3r4FsmJLcZhE5EYDwYp0hKa8JN
cm2hTNZJdwm4OQEMNdQpw+3HyU+s8eKEXzJSO2aJ23aTFEbNNeGv3Rjb1TiXdaH13AlbcRvE/dKb
8m9+7utAgXcK8jVBcOKf2udxi+SYG6X5t4HzS5d5kKEp+TCENoZWYkNACkrFfTaxt7nj2DLxqtag
IfEiz1M+HDkdvD+CZx80ls8WSJRqyuw0RsSrbsHZa4QeyhiGhbEN3VA4T+h/T3634P9ch5/c9aJ1
siydUZh7WDbF5qmK3l7e+CRyCC3TMzIOK0/xbvS6IYKjPVTJQScTA9K8L66Low3ssB00fYolXvY0
1EmtOMxS+cCcEDoTOf+Ifyc+O1ytVlFTUS9vJ8u0+7T2zIhiyGlZRX7nQsjA01Ss8fWiD+a2Dhox
a/3/EpHIisVY1UtB5t/D183WaNBE3kxWHaRDAC72wX3psA1GjI3MRXIOd8IjxxYjDWxYdUpL4xAs
tRFcOe9tC/dsR3zI2qyJD0AurRlDUGuchPGgmv0gqrwZDdegg8U1e6oVDhDScZ3qA7z48tj/kwNt
FHRiTVVdP/G1yistEJ6wvxXIBx9BgRZO+yG4RICc36xZUoTjMM37QjDKjB9oAF69mrCXhNLzRItR
eZ4zsLyjY538Ou1B6kM+zre2fsjzmFE+URnDLOg2YpszhJGlNjAwD0EJN+fJv1j5Sd+j0+7wZ6sT
ZniLWAn8uq/xtz0Nf1jHfC0mJ/6gImafl8B/iHe2a+wWHxmJ4Hz1lQoXQFYtSXVaZAcxjNeU7/4e
WgGJ4K3Acf9Qu12O2TjJ5ajslOwUH+moVE2dd6R+1wp1icHUbSrMkx3wGCnv6akpmpDhcAbVKwC5
wMQ3g6foCBLHdo0MpmQDq9nWcMjNSak5Qfn6ETuDhsKNImNhaMvwgzCg4J1/og6QfRL49Mw+WeNe
5BhKjGIvBUzRtqYrdEep6/d2XJeskpxzET3OH8hPAI9NIv5culAgFzlR4+BOZmPm+SxGbzEffGy5
lHDrfNh/GjOJ1kak62sQAPabboX1f7KjbfOyk9I/wPikDLC4xbQGk07u2s6ieBU4h4N1LWOXvVtt
oigTbDBcdmSsEpHXANpNxE12/hbaMjpQjwx9Si0oksApouv2PC6y2cW8cB715jjE5ShISHOBE+/s
sv7ATYam5HJNdoAdqI2y8Ufofmz9JNKEnSHUQZYuxwFIrSX2KygFKFGRVfpckZGrxYf91uOEe3+9
dNCMQE39w6ItSLvIeAGhct+Vz0oZ05KKTJUD3U6vQTOsWVVBKHvI8URW25ItbXzIz51bYRZUxdRd
iqYf+Qm1tQK0t7gjbJesMr4O1lpgGftEr7Z4aZcpKCRscu4J5xTOfCahLFHEM5VHz/huUEbPheca
RH38rm7FV2BWAvY7fQTzkSM44kmD9R9q8nDZW4SL7n01OqcJp5hy5CVg8t2iURmYZqx1pT1l373y
wJnsMrn1Sy4snxBOMQD8Sqd7qBv9sYYusSU8ipuVRs8W6Smw7eKK0xuZs1bn7jE5H9Fpv+SeV9n3
+bfit0vjfVMeqREzTDzZnedOnSKoQxFdF+ZigZ5dov5Gv7+FD2vWHez+fduc/uM0OFM6a1MEKr9G
b1x6IO9/vu9+Hbn9yDDiUIH2l9EmwmrZVuyyIy0hGDfSv3/sB7mPNK60ejL1yShDV3y1b1+lSCne
OQmu9YTpu/V3a6ZlZw0TsxzUXtBLUKCuq2cw9ZucS1W7tvKXmPxVmPKfjMTAm8k1pfre2qsCCDiN
7m2sAAgnFwQnhwpPyers0wsT/S3i+MOjfCeXQoQv4ec8ksGT6vsCEXsQAw3OTaK6Lbei1W7O03OH
Vje8KQ87DdT+jkdiDL8pV9cv5aawWjzYJNFatsjSGe3UnbiZEd1htze650c8D4uENytnuZAIwHpG
zzckfGYsT9LAMpgdDnJiicky+2Td+zrgwPQM5TTseFekDaq/ZC3N1XXbqLCXMlrKMu720SLkpXfd
gc/usUASQru6Ugc3dBaTQLQ190v1aWHDxoG2tE+w+fROjY8pIGI+RKBJTWKuvyDNqGRkHq9wP3c4
SRGQu+M2ctPRtGr0eGcaYFChb5LmjGcTHqmnrRUIw5PFVhvxdfKGlqo8paZcRvbDfFHvKVB06D/6
9jt/WAVGUaxXUsOqIcMpt7Fb6e8qu5n6aJVbOPLE1MbCNzD9AL+IacRHyoMTAy4hDfcSXNFYnVe7
cYJIJR21SCxWPbD8BjyGnts+molrnFU+PrD0AaNLg9KWgHQwvwXn86EuYf/6kEO1j/KTRRQPdSO4
zw6AyqCk4WLvv4bEJXfu3wFOykNAMdZRrTn3E2D0lDi+9KzAluylwUuQrWy4i73a7JQZEfXyP6iy
pdk4GfcnsCfer4wlR/QHOF78WpEODA7rEAQVYNCeQYoNHEp+5q4z2+AXJV6hO6qb5CCo+UpSGp+C
YJu/+WkWPI9wdLrgJ81C51ew2sTm2yRQ/e5h9MwyZw/UxhEsOJNXDd2A1NvCyjnCgytRzdIeKKLU
PdywevC+s97d58KkagenbBkuPIxCJu6K2gqySsn79nAksC04VrwDKeqPclYCZpgLTRGENgUI9qkO
w8CFOQ/WZJhUbbwbJDHWn6likPJKIVaMrZu7xW1RbUfs/mt0+JUaxfsYbuB5l8fLuwhXqqRhjplE
6bJx3tHrdzRpFEBfiNqe5Tfg1RDi7sMu80bLfcKeF3hEfqsVEBHTzbt2scC7gKsHJT+lFDlnnEgr
3jFszhdY9Ux/ySn+1jtLeTbghZa2EvR1h526g6rGTXvMdKi5tuQn+N0mVKUTjLxmpvAB1LVWGnvG
i/J6TtWmi69XSqCWTMaRVw/0JFiR8c7fn0e0+XH0KphTAXePUtZ4QnNRCciCMN2c/yxn8u+FQCsn
VLE+/G7DqHUMtQABxcRIfYo4Dm1eIkgnoi0R/iVkzdIegy7Kc/xCmjSPA+5bLEvaAes7ru4VGqdr
B/06OInkTBVQ2xgOv84buFUnotl2SXT4NItzDIXziQovL03Uo2QiNBwn9JXpr6wL8nW/qIqXWbx3
Crfg1MZd4MHW1TKlnrOpv/LvlW+qBfDnbaohU/S6OLT/SXfp9taPUAJt7rdYFZXuhf8ujbxzUQtD
BxZU94pwZDP6lqo9MeF1GE4qJMvpMVpXe1QqODQPnEYiF/FqDcyJ+jFQPyCF1dah6n8s8cDn7oWg
1Zn9M+lZyDSM1Yi2rFpCIBR9rp+4wga7yKQ1CE1OPNh47bfOTsnItosoIOWMc7T9TT6Qsci7ifQ3
d4VvVRxrtlICP5wzl1IHwaz9WC0+iUctDjm2yCVfjqT76DSg1gelg7lx0xnuOGRengtoDBtp4Y0h
7dxiykHgxEK+PoclkdMSdy+I9ILeSgVFdGz+4J3ZI8n6DA3rvPpYDP7l0AhvQfx7T7kuAKJR5+s1
3F11zQ3nIyu1IAsrHrgzWVgiNCqr5pnzIcEKW7qNpQ8H+EE9BSXRA7+9WlrYaWzS9xaFCXx3ghvI
Z+F81a9MhOIn3t81dosFPpHo9zuGA1pxSSnerUyn54L0q98OUlibpOEsH1mLp2lxAHknpOtd6c1A
WQ1LjcmsHeB54CdcciYWzk6YcZu2/G9LBupShjWdvE7qQC35w4YwRK01TNtnposYDbj1zloWYypm
/mNiUuHifcZFSjV30gYSt20XR+PPlbeCv/05cruTMi/8t/U3CUpG7G+sP4XZpH8lEA7keGtgFlQa
pB1Ln2xQj66xWBRZ9ps7oT1krvDF504i08j8v6HhjxnrtcZ8w9m5edXUx72Hos/MSFmZhidVvgMr
pJbSnH/VoaAnZTv0U6IBiBu6qa82cy8RVYWHwJV2QsANpeQ3HEjDLksJf5AP5TnqaANw3Y0p+AaY
iTaIdcx0EuKNGvkatSSgmAOM3ECOdfU4J0/ev/DrBDJvPxYI3j81FSkTZmbDTqBrNZ+ekzmP2UDP
GlrUiK1BXpLMQ6AXF7t18qFcfOnJZrQYOc4ZJscwCW+1YnoUbeATD08+1kSx5/FUNw+Hi/kyC4GN
MywXDMHnpooKkewv/Q3EFdlxG6sd3mR4QALtlq3VZiXYANdCGVvDBBVbxrqmkdRbNJ5YzcpNkBjh
Xl9LyzVJtDMQN0MSj1xYAulZTYATTeFOF6uY6COCsWtomECH1XpzDUauJF4F1JrmSYo6oSFhSvHV
bmNkbxlgwo2UVoiooX+S+EcLl+bicSljtjPgxOcXNjXEhWSKysojwGM4wuM9yfw2YH0/KvkiU0lJ
109O0+MvbNPFGyyBe82QI+ufqdTIe5Dusmz4ouSSxbY/n3M6rlSIvD/LUGgAaOZm5M8htPPLolbC
HZTxJnrPTRa3Yad200n43nZieEkPwHbJVXVQC0cjEietWKZvXK6xcJZ+VR4GZvQizugWxG8rGGtG
NpQeX827L8TYwQyzGR8oQEJayr9hbgMg7ODWxw6lgA0U5RkaJhnDoUyNnKHjM3XvMKya/30HIpx/
1YHd/7cagjO1Z/6tDOh/FBKVOobTlA0v/9ikxLKgdP+6kZK7U26TaE8ptn3R5a/CSBivI8YlT9nk
uFRTSAbxEO+SfALfvVUDCuMwTyzDxHQIbCm5WcBmunYZmOFyxvYjmE86G7IZEd0kl1OIbvLTGtHr
gVGDTw5juDDv9PksxZx8+R9C3/UUcvRhN+XXCoEy8WekuD5E94j/NUy2IS26Xuw0qbJYwrGj91+/
/LQY8lkgDlDTzGTwukt3i2G9CjPubiOr/66exlJwzt8mBLTIF1Rl7yhJQ9M4+0iFHhE2XGNB67YO
j5Uzigl8b/uM6HXFdfS4Sgiw2AlShq6d+Vz/2jd0o6oYzceJhgd/tjZXMvC7f15QhsmrqsCDvbBx
FElcpkx3+MZHxF2V5Ksc42qp5UFYteHvXUrAivv3gpTVZzIEym+zf3bNVUexGl0QR61HLVSP4SUK
mrFeXJx9CLmbDptoNdV3N/tjzKW0LTbnOlafPQ3yTFJbAm13xw2BgNi0dN1m1CNSDW1wQ034iqGL
fuMa4WdmuweHcNSATclRrkTBA9/hK3QcLkEkvXpty7Iym495kxcrKUrSE/d8BzeuQ+wyHjz6baRz
RNfuKPUitOgzLoVqMpPEjx5YZFZNQ25xsR1FnLMMIwFSB3j0gQhPFpijCRR9aOx5bvv1Ue97eYGl
GYHOw+Ll7pUXg1koUwEnvmoul7sfdeLh/0pRwyeZMQNz5Bdtf4RmIJEXmt1Rj90yXMQzEn3oI6gc
sdSwsGWXR8kaLLf6G3zNS68Jysmk5dYsYU8CBb6vzEwOma6mFYf14ZLzWpzPTBBsERbXqpYeb7qJ
ID05DQxeHB7NCLlILAPXFX+vnT84g4AnWAFNnL6bvwkX/+dkBRiCRJT48/NUd/q95admtJXV8co8
+W6PyfTViNiVHDsm/qYqi/4knOJkTM0RHVycFXJBIS17dfP82equBDwM9RjLRSP82CjU6PyN1J8T
rg7WM4TaMVuVG6xQNGnrhn6yAyKw5swnUQPUmJOyxar6cC9VnZ6UppSn3CCdbTlyy98JU7S4XwH7
kDjCUeN50bHFggC5NfBkVlDz6UNsC+q3xoGOs2dBXHUHF3AiX3wJRZ89j3aabSWkSHU8d9/eAV62
2OolmnoT5AHQULOJRrkslB3Rik98RyE39ZhSRTbfor81eIcVS4Kj2cM2j0DDOwSW6vDLvukkdlwC
qw+zkWTNGXzGDyEk4hCSThR74VeZFjSdKbuDqxsktrgc9OfZhqWT7rH4Lt4VNpFAPlitmndcbqpW
+sfgWgomf+56Dsaqj3RaKZk/tjyp7OmSx0HknV3QUtX61WJQNjBNRZd/E30YskmPrX/LII7f83zy
fbllnJRWiC/qPU+OH1yJTlNI2eaPq9hm4uEKckhjVQlnRgtDRq5HR+AgMqn/PlCmpXktZ9LXDByZ
mYpENJUpkzsySPRVepF4thKXsxE6Kq10FTG0vlIt9i6Ptd5/Li2WQltAXplJTnzMb7BVKD8tvTWb
WoUaMIMOy+rSZfvNeGHKRkiqx0PgxlVyXy/5lFTz9WxtgZYrXNT4ZU1VAiFnjYygx8PCH06tOdb1
jQFF6IltPYIJO+UXKMEgQCzJpT7y2q6NZTPID6Df/V3kvTX9ef29j7TO3wBka6cgOBBlbu9b0nkq
QL7uxyaaO0z+7KbEF56p5xwuI01bDDS6B+NStSwnlfrgGykJKXLYhpy2RccOfWv3JwIgHr+MszCo
twH6JouTkZepVXeQmTXbdRv8Em2L4XcLaosEsCUERDwHFTJ8aMXxV2A5z32Y1qF9xlbe/ySv+mx7
/ncZ74gaFXHlDRfjQuYXGnD41KHwpgFw8Ewpscvd5hyrWh3kRx1KfnGWQChCaV+uZpaLDJb6Pa/o
THaLbNeJGNcFvsPgvhqdg+tXxDi5fqpK/xIR8Zr+02lWrj0pM7gGFhpIyUdcM3ExI9QutoXTrvv1
el6ZdNnR3a3ERXqjmqef2pnlSFv781svJgmVvzKMZFGqDJ+/dzxTWQGFHztCEMkHgR3EDmYpXld9
TENSdCEAvjBBlxT3+Ac8URpxH/9YO/V8YTrPuMY1JklbEVRkWG5NcWg0qi884vU6j0vC9gYbzZwS
i8zTmLdvqtZQhwT0ID+RO8RllwB5YUvTy3sgf0ZXv4VIs9kWrShmMjAwy6DzNYgYHZyMeh8TFJD5
JS2WICSE+08RN7MyTqht5M5G7PbtVcgdcQcrG8BwAzbcI85Xgii/etdq6HaZ+qFvKVvm1WZ1Wcml
0BEJ4alR1stJGWKJrpkJ+cbJA7WkbjWHHftYjnmuLoEznBoyVVQCKe1QYwptZOzzkcusYbd7T6Kt
LAXvxSgqoe3dYqBqxCUdwNmH1G6yZCMfLaF1HE8ShMDrT3SJKkvCEJlP/LdBZo0V8QrxSUsEr9CH
juyaUekR0TFLHj/K7akfcfDGR+LFNKLMSynGmgFPTXIPLJNDRRLuvDNSCe7VEBGzxCNBtorIakez
t1kamS0vOaXzDoBHsS1f7VA0Qw+59unlTlVn1btSOBEu+S3ZdgHIfXxm6/Ri/LyZRp6FrR/eg1Z4
O3UzXS1Hotq3Dbz2d+7AV7yuKQDrmgZnOL0QN/Op1ErlcJw/s4rSKSHpfSqxUiFPqgWIvDzHt3OT
CKUQjTabHrtxArfNt2TcuPwt56eI3SPSY7R+74cgNd6JnjQRg9iSjHQjX2P6KXj0UPhIdzQpFssj
LsIoXSPKqzQHgZxenJg99mhqaA0CXeBc7h/uwC9YyJlnImG/k31nb0QeHlYZIik2BuyUOl1RXP2J
WIzmmlOV4Ob8MDj2pPN3mOziNPu/+zKo42br646Dlf//umyEH/F61Em3WST9N0a2PeEQ3PrJLRhI
E1awngv+4AULpD0K/tw5+vopR0cCUifKCCmqFZv3/lG4Xk3L4BYrpHei68mOShTiXLeQ8H+unAtX
90iTv/LUOnyvyIgkhQfTgP+dSJ5iawhCSL67hSzbryz6Q8uW0LSbfo2kg7EXKJPFqC4m5ZxxS8ZO
n+1F66yA9Z3mgoLWUnvHFbeOwz/RJj2WOpIN0IJxoD2o53lGLBGPOuQVABrRcVII0xaVwy+ux+sz
GX/wPt/gNwvPNQ8PlFDPnA/xCKqKcpDdyA/Es5PCc2w3wSn1cXXueN2u0mYDG8MOWi3AfkHNzI26
lPaJWlCde3EvcowEFDBXaKEmLlJIXRnAlrsZo1pdNrxITbOHAD41EefMfBpNvaOLfO3FV4TnnGn1
+x5A8xJv9/SGBZIiOtzeOUgFfAckTh5a2TAnBTHwQKjHDr0mB3W65SlsxdO6+5iqDnc0K73aJVje
b650BWvbys9zBvt+bMYrVaGLeJOGW+iV6TZjq6PawgvK7d/sRQ8cLTECtaKE9ae8A4yfinZ8Tnca
L7nbG8d7/bl4NJYYBM8Ffxblb4cQ+k1wgaQBQTl1yxlVcCF/BS+ZYMw+CvSpxVpjpGO33ttX3gWZ
BRXz/bBwlX1Y2QP4etwdNwz0t89UyHQVmQqd78FbRgfBZ9qabNdFr2gtHA4FBDBJHYE5ze86Afus
8etW9wsn7DOYJyuJyelAhBzGHZuoEFIF7Y7ZtN3LfnQqWnFK5DqUZe1qZ5O//J3xMvN0CUI2XiKL
BPqVQ7iOSEt0aljPB+eBpNFmzcWfZ2zQ1LwCJqzuBnJO0rhStii6UR+lTqBGoXpfZL7hPmejxOuh
M+TlDP4RQO+OmRP4NWf3bs0w2Wya4C/h6wSYG4Kj0KiUBzlXPKLj5GXSpg+VAxF6eTm6/yXxl8M6
CPSP0Kra4DEoJZ/lkGbRuNCU/ALXOcsfIrq4q68CB7xc5GQenEmc09OffMsR3mpx0PQEE4GQqVg7
bW5UzWjMW3+8WSsdrBWEbURbiCjjOTtflE7s2Id6pId4WDwvC922UygkeW6nN4sN2ZKDpjxwL1JZ
Vuwljfz/BKvksarVwFwYaUz3LGAs1hmCAQeKg5nqkBU0RwtGbQ27BWjp/hP/yvLZCU9z7xHbyP+9
xFX6IDQQBMfokLI9dh0lqOiFlUO3/ngwHlnYkgvivnA1E+ixGZTDfki9CQg5wO7DRLjyQUFvpiAI
lY7z3r/OJvLgcIfUSHly0Mn6RnL6Vg/T6XdLxewX8sLXTRbhfC+nGJtNk1wX0X11kFEy7VaShnPo
b6JD4yPeiZ9Ziygjbe94krL/xIUfGurmxTDAarW8nfnSmOCkz8nROhBaD96Nd8aRWor68cnCNR5h
KrvVlJnsj/ss/B9/dk8rONUQU6RagYyO+rmHvGwwKYshlVYhEz8UrcJcSEYHJw0H8wYgNBRhqjGY
XlMFUbjbv4qD0dBYPI7W55Gei+QzLaMiCf+bsG4iRW3r3aIvcR2xtMrkaciFB6B37c31s4aAAEod
jopzFiSc3W2fMpDCenAZQk/XILeKBiqpwSkqEm+oVOFCWeuhTKRAy5hs6kyebcEPGlKY+42q0BsQ
nAeDfeYwAxKQHuKs8IE+bFFrsUMWeYwSqqKk81s2IkKHbSrm+eW/4vfpBr2w0b8tR+JyjEV/MytD
WxFc7tlslxvLJOb0b5VL+KExQPhJdP+WQVVfyLu0AH6UkKbNbLSKJF/WTVNdLmSqJJfXtrj/Hfec
7to6C7DEdmCJ0FKiIKY+sZ6faP/2+Ou0EtGZqG88n+iEcFfrlIC5+hSkXVstZQ94CKvpccbuO7+1
igac6udDbmll1Ed+3tGP4UmiTal4LBlpMwSLSO70SbgRpqaHKYuceyFpFDlOeCQfg0eGITO6pBHm
04G5GWIwnyWWUtaWgzxJ3jr9wRj/VBkvu6yb+znmZbXjwkYd2EmePqqrm87k5H7fWH3xHtfr6vRu
FfAguD8YFzN7C0TQ8et/5UOofUjI0No1My1q/ulioRK4vXsyyI+R0uVnJ7onUTqBrxsqcgxv1IUx
MQ794q9c+Yd3WLfKBtuQqng4cGfhQoM1I3D6G42DXcxke7lpqsbbG35q/Vfmi0CxASwLtN/S+K+M
gyuHbqdPjpMnqSseVNWp4/ogqoQOXLai51erIiGs/U8+I3lmbi/KqM4UKGLiZfeMSJAXljWF9Leu
D8fJiMBmBWRNr9FYFPXimE+FzcetNQ7hlSABE7k9U5C+D69GAhKM4WhvfeKcZ7p4ZycQNz9BQkwc
Mhx0Xs6g/bdNTI31kAQUjMp5HWKjKP04bMbC/NHtO1jpNz+GEuYx3REluHkbesgRcSYP4KOTb7Ea
anCDwUA/6NmRSWGXqDcPTwBMUGkxB6AlJWwsUW4J8CtpIQiINEgxh0MJkhMxJy83BR0poqpZWq0h
HH5Pd8UR7rzH+DPOiw0qvMUO1YPpgO8BCfQXAdyoxxfN/gIBN1lKbX4Wn/Pa0fGv6ivPixMdkZ3N
1R65k889BvHuc83mi2LOkseHEETtPmZrj7RrTHWxXhGftI0CBr8mPXkI5Lsni8mcpL306rXzKLrf
gm7F8W839RJpzhvfc5oqe4zgGPFr7P++H1rm0i6bdHPxHkXgfLvHe2f9d+pMxVuGfOZcHNL4XNYL
7511oK/0Qu+5GdLDpiaTjsA0+0BmDBZiCayUWIlRufrPwa3gYPjRenibpPLH64Av9Z5/e8e0NOJ6
35Uo34sx5G0Dr+hyMzmXst+bvpyaZa3ZBCkDWu+bUzLU45y3pwYfCZwVuPeEBLZJl2XZ7nquGG+F
PTwcZfY4eGgvJ0BP1Sn3dAUdu+33TZQSXRtKdMMYA0U64rfXoCQQVV1iFkNnaOHCUFZVY+luxNA6
MK6jqsbRH3qYoM9ChtxxGWaxKSES5fJHHBCh3wgwsprSjgrdtKZ7y5B0+1tpmFJfKx2LiZNwe+R1
YW6iUqPGJR+Lg48oSvn7bq3eZoxPzfQS9WkjimppjSdL2Dgd81yDCN1jC+I6Phl/apWya0EVLvmh
WP1asou92ElwkF/iOf0+SDUItmPZVnKbElNtRLVsp2SoPayzPeKXcEmQIJTb/YmaYO4CaXv78xZz
XgAfxIqAW2h/MRMeTFDTluMQ9zNfjBjn8xkPtAXji/2dLZr93La31uuX7oLalXiMLprjwtti7r6V
y03MFUpHUv6sU4uvbyu6GhtfXfbcUjlRKideuAgmtiuugYi7MMCXDW41HHk6YxquFeQMNmEQJ7Mj
eueI+JY2XzkaVa1aHU7tVkWCFGmh97J8yL0f0YhsC2rm5KcOf26/+k905lm6kKhnoc9VmFXFS36m
FRgbdVKJ+dLeD9IRv7sqqToU0FutEzWzf1Eg1Ht8R3q6KR3xNuacHPrgG95A0l5gFG7Lm7C+d5JT
y0nmdrEA8quc5GfS0hWseBuBO5TB4q64oAY6p8O0S2xjI9cYUOmCNq/CcwYDFBdfNgDSGK00q8Fb
zX+8Gr1zZaAeKhKf6LS4Bezsz9D3nO81LvDi7X3vdSeGG79Ev8WIJkz+UAT9nG7FDWgYaW/tVh/R
WMa9XG7dbkjqccVoALCmYiFO4kbeMhPjcWFI26os2S75dkq4p+HZijk/r9hEM0Mb8vKA9UXCRZDD
AWSp4uOEUstFG+ks+6X09WPLrX6h6kjzObxR4KB4T/8/8Epezzx+CIs2YryUP2iFPN/9H2zgFdGW
zCy4JRo17XQcTIXXg1H93Si8zdMKo77acLyNii/ScCpmjF2u3126Gph6E2UNnxadWgN1Apr8zYKN
78bttXAQIRnTBFc3NiJBVCYW+UXGWOUQm4we1nTfGBo8YkjVTZuhZJ3ajWuR305WiNXM13PKPOmc
EaMMc4Uu9X+buDZRUWnKktGBOlSsQpqy/GvA2+rt9jiGNvCBtpIs5k1N6skA3UUshRUdA72cLy+1
tfWDd4kJEEajSL0Ge2BmL9lucltQ1GhoU9YAqhv94JTvqxpq3L+U0PpnnKoEiQMA3suPWRpoH6pS
9ppIbE5vurpwIo0WIlx+joxBCz+B60svZjD5XGWNLAyQTDQs3/SQxwKxLT7tIUHj+KeHEvhKbRxs
vyTd0fjuUsFG45a8b9sr42cyS66EnECor4XB/iwTk9GyBV8YT+4QUzWWyJH+smrjgmPxDbIk7EXt
yp1bm/wNr/vCG14PGL65v1wEb3/tUwsvHKrB6CbxK5PpseoXWT0h8/eOSkzIBVOt8uU7I+C0uoIK
Lt5ydSdDvowmtFnCHWS1pGedmaZJhHbMX3jwRBXb6ovD36sn/21Xqs9WGK6DPSbSKL+7XuiG+kaZ
cJaxiJAy/NvGVPPV7XpdNNA9FjLaYZpI1Pv08TWVIb02UZy0nh31SWUyNHC5glykodmIIIFakjV/
mZAZkLjOjg3KbUEke1xrWKQ7YbYvXyn+vAhMH9+YQeSKBmM/foJhrntM70PM/1U6xpgnD7bS3UIJ
HWfAfKuVSkHQYZv3Hbx+TtGdwIQo6FUgErcP8LV0EjDWY78Bj6xVHDz/JemK84VeVuMqZM6xfUWy
MQpdaAS3Fyj4SJYC2blVTHPq9tMgZ0+JxewaHHPghB/YVRpL5y04PU7HGapjFmx+voyZ6soWs89w
AdyqCMrIvO/OS4T1+upJWPV09mqbmtAafpzyA65jLmHRqIqseCUp1w+OWu4qVmNF2MoWTZofxqZ7
517EyH16Wdie5PftEuKczI4L1Vi92gY6JlrX8CQJUXe+AFoqWtCSR89E4SakrRsyz9XXB3RQ4KEN
Csj68YHm+SgCnnP7QI41bCRT7jfp7S/iJZ9C9P3NFqvlAChArAPF6Utj+VZU8ABvupFnPbsNcpdV
18rNXWZhfPqVh9aQazaewPZRr8p2qYRYBPsA8bagCT5p0k4vKW1HC/tqipZlVmI5P4FvyaTdYnZi
eS7Nf9NglbxKZjE+zdJg0POOoAZOlRzbk9nPUAzywUOmxprlQ79f4stpw8ox2whUTCtt6ngo8ej9
Eu9Rn9gw6Xv01ayBYP5/itftTAxSW62Z+Xd/oL87Owkhz+36JAIaZIrLEAdjfX6UxzY/oji6BoEG
50fgUiZp7DEdNiI1HzfiJE5yjOqkfWpzMpq8rk5UpZG7ydKZwaF/F+eKap7fVeExLc+MHjlMJibC
iC3MNzh++W5hnypG0lN1CgIkGy8hkhNGsC9/ooA7AX+Gs3pkBlrNgG2jLxLamy86lwsK82w1rNcq
ch7zEVg5M53f6BKBNzg3Auc3PaTpYfzvhgYXNibwwYzuXYS+o3WM6+7XKUJkDzlyx9L9CvuqUqci
hU8NfY4VZMo1ZbPv17QCv/xO5xQT9Px1zvnS6CMq8FYZ1qDBB2yHxqX27CAr14Q3NVdaromaEL/P
LOtq3YyvS+offEvr2pFFGGQnwDj5KsKVALNU5bPyKC37Xgf/eFaBv77Hxn9IrW3GmfvrItn4X6IC
YoZ35JJTJnDlu1UVcMeX8NyMPabNNxJSPG5yX6KUu9pH9Tue6wLCMXXV2a62s2UlknqHgipoHF8s
q3lgHxi09zv3pSSdtrvNeU7XrvXEyA1q0c9uRZ1pWseDzbEaxA9kFmnyGjaZ6ycFMSaFp4kuwfOe
WnFyNhebw9s85gGrij++d9H0Die9EdHIr5nF+LfPIr7scVn9lrlCv5z2AkxyNWmPgJpwNCTanFkS
pcXuEa7q4Q0A94itsyhcL52LHHhke+vgQMmA4E2B6qlMfv/DiVGC2mUi44UliCNE9eDRjiBBXOwk
or4gL12Fy4sBYG7swKM04kHZtO580bppd8/mpMvXig2D2SnnCoEFOHbuTgGp++jc7rENsXAawlXE
9nJHMI7vLNYrShmAp8w1Foae+QVK84jVD7T5RAMOaSBDRX50HMrkbiQh/z/6ZO70r9rm07jXl3C8
HNqaCISDY9NvpJLz/3ycoINiYNgVeViGvAN9ce2vLJolvk4483vH5sB+8ExYvjBFVIX9gC+4LfPb
hkeYBFC2lZpVXdchlNLK49ArlJaZ6zUv7KhDkfoZdNA9FL8B5pzt48HliENgriY1W/4jYg0qFvK3
za+BfyqXpURKGRSZy9Fo/vhlK1GW7dxGBTLyu5dXeXSyZRP4yLu1M3EnUqX42zFTM3A+GB5mKZCI
iAi85Nmi/srHdagk35nhopvFKXV6JfEorul+dyNw+ytx0ScBjpdbSrKk7gITRRwtij79xbCt68CP
8+7gZqlIqnAzcnsfgWABwjoDLUrLh4dnR7HhLcwxzR7WuUER4iwrfDNYxz/5uFXIvRrNmlbLOqFu
y+n0Ha6DjWCHkm182zhBeCJx7NvG/3gPKmxh35+xdU1UDxPBsner/WzniZCsC/BlSNItw61/bmkc
1rcT99U14jDwixblaUJ46BT0lixlxKJO2vjARJEHE47qShB60fCyFuPDmvjfCqfGbtEyP9XQdsma
+ARupZKNsiry6yB8XBpgYyqshw0X0W+E22KUrw6VCxfV7zZzfF8EOqjcvlq5JMk/PnBjqRZ7VGYQ
E9JF0DA75GAFRhPIA1Mv7KCy6UCmPLL4jJP1BteTO2fw8Gl8sIg6KO5zdA/R8PpkRu20mqZfrInj
1DDvirMTiBZGIjpgotlGGjQq6qIegmXWE5sAAN1r3V1BwudjPxz6L7g8KwBUEbrz4ameeNsuuzZr
VfNv0nPQek+9OqfY2ErMglyS9kXDPn0AREZNyC5scPB9+kv9QRGrDCy9fF0SKKb754KLCaj+KQHV
kwEO9ofLymYDn5QLZ3oC9Gfhfg9gPESzqu8wAR7UcrCNjuwIF+BmddQOpKq3BB1fLEnwiH4WXdk/
r7DdQMhhpan2ZEIpBpGpk/9Q6/7fRlb1klPdSl2wh9m277w/Guk+qg8I7W9SjZ81j+dgXKPlVV+n
OTAJvuXY9UDjKMjbMyadspjZovvWY9EAXAOIWnkth20OwgdHDjN/17FQpkHhZR/82fiR+dh/n+L/
U8bpR6tfN2ZdrIGRnaywhTbZidGnTGCdwsXPNfFDYBCIRRSz374Z91QgqFSXJpjCJidRRF8qr7+U
ujgqEktiIuUIE9JOEpp35UVrYMxYuFMUJKlZsjTohL9kApyZfX9TOnsQ0OgqGe7vstP0TJ1l3nji
dLE1YxqlMK51pOWXyy9f/G2jvCY+MQ1D06vAbfRJhgLxmozkqhqAjltwc5FJz+v7tMHlIv1MExQW
dMQJSxfePcJiq86pXEhclGzd5ZWLK34qc+ndOpDA8iqoDo0NLQ6d+Lrh5m4497MpeBPwqa9QCz8t
zVeDKzlXqeqPZMHPMfI8rzdrR9Orxfqax/YWZuCJ3rzX9FuXPMSuz/lg4W37G0uoWsO8CZrtZqoa
G6OWmWMFSPFq7MhgQv5Qu9Rmy+WF+unCQoAlM87oXU4Eli5/QM+VNzIuvJrldObr+lzQfTpOUvWe
RYa2gYJPkhjKG5vmLfYlq2L5C36tOOD8Ta9yEi5IPdFKn4lwZR/D9tK1FY66p4/jMQYGPiTi537f
rPjMgXzwOwyvL8qxoLFSSkLexN+AkEX7Wjmv4xMVEcL3e616AsQRw2XUTAd+m1b4OuyXgudclZa0
rY55ut3rKdcHOk1q8UE3DAkgSkGOa+6ULa18TV9k3Tla6ienTEGhbVRo+NdC5Oci2Tz4BjBXgx3a
cJpzui7EVdOy+aYdyLrGxTEBv69ZqRJ2bok3TAQeiowJX86gH3f0W+YVEdfWFiX0WGWI02pFSyXn
K+QjIBifu0DSTGURkT+zvYe11hrjf/1KIjvXe75s1tweMGu8S/XGFysbfDftHKa6w5KrZKNx2Sg/
6fVzs4RefAYYvRxkj3WcAVlBXvz6QrydwWmlomGx1zPAMOOdHauIwCzhn9lNto4JX6pTsvtUV3oL
A14yVY+C9EHZVFHAxtwH8IAQZLMsZkOX+j2dVWSaWjXfHGkIe+pF84i7ioOqOsLaqzqI4gdjoysd
0WzQhqBC5YRj9kNmt+CYmsoIOIkdU9ZI3M5QyJ0biCcBcnLPKL7QAJ2iNxPKZ0gAlOeANEj93+Vd
NaTnvntZh4NfYYjQuLsA3TQnS+nEko5OeqfVkR1enUBxCt5Cy89Psfn2dAuMizDGyQf69TvUoRIT
Z7qUqR6egwMtCsjBbSvfx4yg3ZnDtP/mqAglUrRdgb1hXyw6VYzyccQtHwXJW2ZvfNq8gYNTBZrl
ln5k5TejXKqUcetbyYxzM2I/Yc7TTzLuzzKe+loZL7dcpfw4PsH04QfHENDdoesiQEsvzbbhxfsu
YNsQup+Y4CM3QzRUZmOOif2qRYL5765jdxZSYG68Pay0tfABH45RxI3YUbyZEMFuuVvKb/zG43vZ
AIJ1rVsueSg5WFPR1vDroWDHXvxNXAV4gJM3GBbQmnpMmEVahUkxiI9AWYJ8FBYyVqHqYnZ9QBVb
vxTmk036ZEQ+56ow4hcWEA6yFwXGBxpLYxtPya5ICuQjRyKDbx1Z46mXl6a+8taRxmLtK2Z0Zk7n
jNmjp7vipKd0XsT8puTZ2G0ACaAmh76G9W4gfwmQ6YvhV2DyPgnp/NUMdMsuO+9zlgtsQw7VaaJV
YsBBByDdxz/obz3+N2mDSYRQDTGXyBnYLNvgyj4OEl4l21NGXxNOb302WLtEMawQpcJPr64YOdL+
WBy+DBlJP6W27tpMDBP2UxLebH32Fuiezlx7Ph7uzHiFV5gxr4imn3qy7EVYLd19W5tOiA7ZpZz4
f0UGthllXBbVjo7vZuo8eiJVp8bmqLV9bpe7lhJIPGFsGDhqerKUhUFrzTAoLPQAUc7Mde75WJLb
jpfJjEA2yP3WiSciO6OpJtNT8+YEfj0T6y4piMKJXYVak1tH2RGrSIzEY3R4mMtBKx81psyvT0WV
ZZJ3Kfpu+Xk/leCNMPpAmgocuxvTu/kkjB+D2Ru+WWcyM9k1IgdbMadqS+hA9hOa4BuSMthYDuIw
QENOiQIX6L4kgunEalMH3ol6ejk/Y0+7dXMYXgCPiT9V9aa1Ud4xzGyDZ5bqUwz15TfJf9fhvDSM
/KdWjhTuHI1VdyGRM7t5KQtJsMGhyEHKJ9FcwGCjDK6xtQxolYNO5KjfnBe2a7KvTbAXuhLFU1LH
IfyoKFqGlIjcfwn0Ov9SGD3U06+S45s1VtOm7wcWj/Y8Xri8XmitVFKWObzq7BKNZQ+D1cdI7Pxs
WEfSs3n1PYu+mC7aKCyUCXcgFqnzBnh0qY1Ub3Z3S/wrVbDxYDMVV1iNunYAfSwC/RvUbrvU9SLt
YKNIEAMgnv763qD5rHGgQixYaTMe3Cnv0ZgC43DKJNdoW31DuNLJcGyUJ2wWmG5cLjpPOYltlQ+W
H/ZdTLa+lg9JNwuq2q5vMS+j5caXZOw8KOeiiFG6qPa7vX+1BfmlO/y9pKqII7Cfm2ph8sHaW+gD
6e3vT/uMnQjKUw7XxKuiNlx7q43dAW1bXAs8k2ErnFPgV+YMkBzEPzYfpOyhp1cO41FffqA9o84i
fdn/SsKwGbvNaHndomZNGnzdrh4kc9UQ4t0OTEqNyui/IqYydTAbHmlvb9aqNyLVigeeBeLEMPV0
qX6TU5bIPmex3hF0GPObNeN396f6wboAvS/qoFexvPy49oFPxZnm8SbWfBu0ZZ9jeOhiSA1085ry
0XwSD3d+XyDZ6dHzWiWaD9DgpFwNrrS0jMux31IF1HexCLg6Xk7KYz0U++vIRsReSpu29Y2+1mRi
q52ebd2TB3afp6Mcb6NSP97wU1AtE7D/MAwYnUcwQEV8pbUMdQO+hLv+yZamijvcHIly9tZFAnkB
DNQW+0k6iDY/OfuKJuH9tza6sCARu8tK9ivD8rBWxbrLyeF20YzyRpNdcHuK+ma01mPMSlAnUjig
YWKTyvvU7mGZsZ/12O/ELQzOp1I31Soc0zYkOiUc6Zim2mwNKA2b0jOKAQJbXQe5Xm0NAfFeax72
eK08HTrXfxKSj+udCdZd0b7EYF3J9b0VgIj8vcbMGy+t4pLYTcIvxwv62WmR/6vcyqUUhFvqGab+
lmuYkqtvBnDY8Ku55DWE+jIRhllTOTGBK8JJEqcezyzjM/vUDPYGOq43xdroffbz/FWZFF0ozAzi
TshmGoSr+kn+g2Dzlp2+LkWeXT8bRrecyNogkolJaCIkLKM1BQbo+CYNXZIlOO06b86gXqHao0JE
ONAnkynShu8VU/UQdGS77blH4LvK4MM7i0gtiox1OcEAzsXsMox93IsVpfBLwqsl2TQsMr2Xvm/4
7jR2dxOcFdSg+xVBnorbVpKAeK2cYm0HAuqjxtU3q2LdL+Kn8AitcS2WTTdLDzdW/GPLyMIITAli
+HBv/5AvCgscVzmNcTDT76WA2sFlPxAQLImQ6Z3aLT/giI54Y+pntjV0769cXtRYNu4qZR6xf62D
DastG2d0VYXkA156Z27hfOYmlyIL+QYn8oir1bnFiA3VClj2qC0gjT3R77i1p4Iv9mEpKabkFFy/
QYEARCMi3rYw7eEQtEAttGdG8bgNMhaHUiHkBFT+ssqPYhmZIDLouoqRb/6uiFlbt19kQujrOBXY
dSfZ5G3jYPSC9sjFyLoeSp4GaX3Lzqwg97NiiVgn7BLk8zhePwH5K6cpPx5mWMrVTASGNe8GsyD+
cSe0RaO6th2C8kdDqXg0WluzkSCLfWmm+wAE6OWIBUHWj0dGEB1bmvk4sqOnPy/qOgOQFqOh/ukn
c6bgLhf54x/EJKLlpS4CHGr+26XbyqYxbY//XISBU9eow6JYA+L/FXa/gASAJRMnm9Ovaa0HJVJn
UwAGv+PTiIvcV9cfsh7ppCB6/9b4mqKMXA8cjFS2NvMRX1Lv0SaW7sEOCI2fQLtyLNW4f/VnjcW+
oOgZszbOtdf6Hqsm9kXOGXPQjtIF2C7ZmGDTJoNJpJZqN0rte8/lRJ2+aVeuDpvKmh2XZgXvyGYe
BHgP/X1N4CPajeU6k6latlndDRABreXDOO9FJFL8kYa7ZEq6wNuq5k42eVUge/EadGkGjCz2XW8R
gE0DTvCRBAKtPeqxxPZ98c/IP/arBuyF9CAwMiZ+C1SP7AXmn4dScW+N05L7dWA99Uym/XA8eO/f
6Wq/Bxkeqi/1O33NA0csu4EWygzBc4MVzLUFYkTtaBX2Fccnut5JVuXcoccozstY+R30w413DDSv
E17830754tUuoDygc4BIKfjr6sA05PlzTNvmwe7u0RE8ENH58iKNftYXCA4wZSi9g1XZ9f556tm5
lniFwUYb//NUJDZv+MsT0gx9gNnp0xzIy5eflyHw70PJpUsF31rkNe1GHT6Ygdr9bG1+bFCt6OMt
0JTsMKeL7J79OYPb9sWBgqvDRU1ok3I6LXcyfJ4ARyc6DvPeZzO42Qpv0wYAwS5F5CB30QOyvrfX
MkZXXe+/9hBIUG0KknDYDvwaOXgSiQDMkNoCEewbegf0DbwA1RyYgmjzbciL6MC5Bdv8/ix+Vag8
+VmKkJeNmQSekPXGOyMMrgEFqxaHrNQuY75P6e+t1RCcuKEDVqsc/TBqO1uChVP3uNHEdPqU2ZHX
GPmBbQe7yqnzBYoratqh68poadTTjAA5lvmiZvfYhb0CiWEIo294q29dUFIWI2VoFXudYpFjCYrF
o/V2BkQ99mPTtr1dfCDtKT1rR6IznqtUX9Slut43dGjKxuSyfYvAOg4QQAvgRVbtAgUWwJQLwrz3
fkotbEx1oJ6tHUF5EHNt4Ia75daylma0p/DST5S4J5rp4/rw1ARE0qGcBEtVN5hsc6dsxNeN9We6
lc8wxOOxmqJB15suf2X3Bqoc7657ZgG/4xGbL0P5FzXYOzEspfPJMC3j+ary4GLAYuH/n07YEoAY
M5I/dvEmW1wjxIPrusCEOfyWBuJXWGzeVPSmfa3J0v8dip5pEIWCOu+QiRqi+gLDSVqOH0i4H+09
VkbafwRbto7u/igncuy5HPUOdbzVmRfEJV9K+s7CFejj3S1DP6A1e8QLyi+J+3/LJEqjL7baPjaA
JReiqF3H+RJFkfERWqrzlevzHYVKxWByo8R/vZKXyxLfE2iMtq56Ehy+IlAFJI1z3rqPWZSrlvL3
xP9d4rZLwo7MLCqUb4yKu1DWfBd4JREZrZqxGWqdzD+XWnt57Y2JVKP6k7YhtpyV0lWJDyMEqg4Q
ZE8H+3/6rPOCyKSoPLE7Whew7vcyBGJ78UsFsd3etF7/cbB60f6O6xRfA/wmbve/RyLtvZ/K4Ul1
7de4o4tEOODxO276fdfJjoZbXVjWqljsu4BejIHdh4/PA1HvF12I8Yy8OeSY6fRbgiH877df7LI6
lviVnfSCJBfgIEyqq1L893Pqj5M2b/VIhIPLbfch7lQ3pk9aUsALrS3KWgwjuP0PT7aq4xwTrvLL
OVWWVzsuWoSV3y05umSoH/QsO1FU3/aDvYedUguy+/quT61SRy9Xgu4hw/DERZ6SgIsI46xuzq6U
l1LaxGfeMBZBJWdvtxWcnn3gN3C3wmZ5iU6d+3Cpllo6LbONgorzPdhqBaW/MCBXRBlL9+E2r7RX
4IzIx7Ov1SiFxo1Xmeb6pKtHo1k7rSfZqtxoNCm844ndxXQPp8OVt40D9UEsKoWioBvSQahgO1FU
7A7Hsr/MwFgSVvmWrrloz/WvbJ999cniSe2KqCL7W00v/Q+YfOsc7nLDE1pQY6zBe/U3TyAa9yoN
tZwAZZO3s2kFOqo/YG3yC47D+3l+q0XwghhNQPkse0fIzLXPw6ekdtM3QZ/w4oRrYWJyJuXbFp26
ef5/B6lt5Ee8QM9xhTtdOQIf1AlcKk3GHbYEnUOOLkxZ5NWq0hxpKj5fu7B/LVsf15cf/2pl/TSP
BORsUt0u5q1hygvT/6Mac6rsvA9nvOGJOjd4y99o03arkOk2qi9G5o7L3f+g3DVpudTL0pK5hvpi
a5x7dDQOfqFfkaQEJEHLK4jDVRP5ZeKCol97UiTtIbcefLVSrgb05V3X5FixeQmFh4Iy4L7zYla9
c1Nb0Vde3AZnwIA7TxTbSUUdbqfhdR6O+6MNS3jxg7VIIF/dmJ/Tdhz31W65cVGQeSe/tDVfb8zd
pWmsAG1tMPEO95ZKq6nUHvFDEos+7btZxrhYnt0DWGnPogF1hMHshVEKucJC0IflwEnJD+M1blwv
5MHx+ZTGHqPxOU9E64/+i+K/PC21OmSejDFnbh8LoSmZTeFWGoh9wbahNTgqrgvRBy3qokxG0a5k
70YkRNk9b5M3tEAc63P7pQnd3pa6dAcltYcoe6w2mIOh9YHs1gTAptdMtXDkHlk58bohA1qaVqWZ
whBu2xzslE3Buq7dN5I6noQ8fP9NdmdEB1LzA11xLTMqG71GU8wGBdGDbRxpHSQObGAXJuj2At8V
Unlvs2ACOkz+0cpSgS7/sJdziN5M6oqPZYpefIGkw0HMIMZEURX+orG+qR7FIzKXJppS5rO5UWhq
LWq9oRrGW35urjH2TdkgPSwTPShiRFHn0Mo5XNYswJnBpXp1PiXSJo3mu+Oe2dTIunYL5T6eG5G5
ljN4HHgIZNJV40DreAPAjTG7DHll+d70gbMaJo+lzO+R9gZOdmShzVb4Z3BahqRHkWH0MS7OG2vh
qEZZIlkWJW8ppv6IeLzOvw2RTUd6CK6dfv55l9t9qtrDtHC61rRKc5CMwTmO74knoroCtB2EiTIR
xNi8EAf+1pjQbIqx60bJEqegXfBpLFUArl1xXi7aIZQCMGHKmw8yshpJ6ecbVcOcKZ+rNB+2nG9D
z8H23M5Q4sTcsYj/E3E4IthqRF7pkhMbKZSFzKOmrqvXXmVDOh79wDQ6VKdU6mHB5wp+klvHmX0d
QgZw1bkaST1XbicITE4NBe88aWYudA9OiN54Gh7uGrdpD+T/2BuZy1rpwo63wLCLUu2GVYlHmmRy
fbuJeL5Gl2OaBhKpqIQaHGyP6e0AvD3XPK6N3zvvSZ5+7TDZ29PSqwRkqDb9775fMGugNVC8Rvin
2q1PWe6ai2R89ZzPFtNS/rWFVnqs2/6ZIfSkko5aU0XtUTmuYoGfvuTLtz4El+UUbllGYPlqqZch
NBGF93KuaClsMsQi8AeBVnha0X6NdTJ5p8MJ5wKBfaXYElckUoHrypXiOSdgBgQ03VGv0tByylRL
aMYCGATF0srZBbHZ5VIJigpkIuEhOneTKxaYsVbhdw8F1H+Jt9mrArqJFfU9Hu9ve9Hcbh6gbct5
+8NzQUq2VMPVzlqmPYVJ98m0TSP9j4PXhoTPnCPJlmMvH0E8hilDYIOIwN1FSXGUioLYXfcn8ewu
o26XsZNqV/G9aIB95NgyuQgAv6H2Eeqd+Jg4W5m0Bn0PsxU4rl2zBrB9WcycPYdc9tNGc+3WEFfm
ZJh85Ay3N1QDkPhj5tLFz2oalbXMdn+Y2l9WL7YCQRBbPyUDxxYHUQuZsecMQinLogk21hQBsFo6
xKxDYRCZC7zfZogJ8p+TsPXH3eAdb3kQNFHyTWuxwSxc1jG5eJ+FZfBjwS9u7xHud2joIDfCCmO/
Yo28TCOkwc+J5JdxaIx319BB12/6JvIRqMvO+LqCZ5rikWi8pcUELHI/kbg2xZ8KlSPfXPNa1ioQ
+ndehDOJFSrFrIP+AadYRsiEFGILJzcqHvgt9nZMPeMIpI890dui4XpfQ782+68FTrZY00Rik/wH
jKpBGxVEgObPymLxKF+tXKbSnwq2VtA8cdn69MlRpSYN2poIQmcRWk1eDApNU9hsq14ocmjb483K
p4bdhYBg0Qx6rTm5e1vkbpqcEdbiE5AfAijvLg7UFMiL2sfFP1Io6u8Ixv8c375OZd+bwyiXO9K/
QeGSA3NrgCvYefWMnZ7FWraQ/iWswIMaCsxTs8GpyL2TQDf7JMw6eOOfXpPrpx0CnJg3BUyAhViN
6U4elotorNuvBH4+r2bZYFek+YwjHhLie9U2k2KvOJJTZVEzkDfTOezG9jPfaqCq/PLGNF1/aM/U
GVFJOGDb9rVzj6og0ZDOvRZ2jCrQAjSrDkCFKOjC4yT2Ha4jqQJ7/8iQM+C/RKtqrX7f9C9IYpD9
PZU3RNGMvi5e+g89CQu/l6JkpC85raNmNEFwyLnNZhaSe+GPYb90YIyMsYf+VimBMXm5u4EwzZyu
4g4akOYR3t+XVHZESZFlH085uUvUu3G1uk9OO1r/lBujPYm2+wKnE6YdEyruZ7YCXTxFzHnD30ew
Oks69SbSZ/EIPN2OgDA/UrRS1SorC0RwLmJe93BXbENlA77we1DBIxf8CJmj7JO+UfXoKFHAdZ+7
nCZozyC1L00gWbucXXIezQilnlk5ERWIByThUBSAhoo/1a9zhxFNoeN3FfMSNW8DU9zmoL/l37QV
4P9VOJ6FO1jjuPUHXawbxF0aBBTxiHmGhVuun6FtYkdqoQVevsB0UBPYKXKITBsnMdzNEe6TeEqQ
C4IGjdxcKG6AQmL7E94tnnv1hifx42StxcirdAoXaOaeQjdhRu0lwDYmZwB8jDQ9GgGACWaRJIFo
b1YV/HCzBWjUpL4xWKBwlcsImwsU99ramZBYGulaLVqwN3EnBltGRTI8qSzRs8RUcjyxkPPZ01Ie
I0zotsXmMSeYC3ia8W+VmMfRFGECGybaAlEaysUVSq6bo+4GwuOYdSUVXkLzSEk7lhb4jCO9dOMY
xIhAyk0pHy8043Jpj3D8fU9/pqPnrdcrfZjHDc7ZNt7i2IaJ+6X9bi0bqlZHptAjOJoxwSPx8ef2
asBa8BdYFoV1j73PZ/T1zrpla8Ch7fdo+nKNjcha7/d/h914xYNXsUXELru0nbAJzuVw2+RN0iX1
ek/34NMu/IRs6oLaedP8CLckUfzgbppZXCduM07+gu8TPpdoF31dciptCGn2UbSYpDr9rUOrjRV/
E7YTydHPrXE1cwyPkVa6vSkum0OB9qiC8EQW0qk+cSxjHG0chr0mq6Gq02XsdiG5A8q0F20CBUgP
MFNrk0DYyoDW/HHCrIEoFkZk2tYo/mb45RP29xR+T7X9FAt0HwHmXCaJnBMryxmnkH0Z7quQbnrG
ba14aaiEs/QKE/2gYDpKv9G5j1aR6xifNn+GBxNxwaRh/5kqWtQeXGSEDm/ov5gP4zQZhFvco8P5
d75BDJmg8zbrvk52jzhaGUIA1gIuJgWsfiQ5UPRMkHUlPt8hzkcS3iZLx828vSJYGrFWkKocnkbw
GwfErz2f1B7sknMH+6Kdzs8Tp5sKt3/5uCuZ4fUGczvHU0vhkGxj+JD41ylXBsSW3YHHL0k6Uh3X
7fQruhrTQINwwOqt9XmEKm+n9XVlr8TMqrJcOLbvOcXc1qd6ZKZkh/YgLBLT49VcLuXRVE1rWuQu
fcj+bYHIBBaXpJF5yrRnn7H1fKlgn2MH9Lv6knmuhKC3ReLKXD1PgOOBbH6BAh0/InmxuzCwZptt
GNl89IVanNHnsH5gubhvCbv9HWpDS+2jgyY8VNYV1Xf7ShIF8NV2Khsoc7cCOwdOwUJzy8Bf7T1d
p5QgHNSDPYqcTvEsuRjgWqAuDoCEcQBoijfhhojTjD6FznU2Q10xnTEzOeh5vM60uR4eD+GvGuJT
jFqsE7IFHlCZztt3JQbuFM+h9avkZnnmBlCvJQKzY1psS10e2G8eHQcIB5dK+quz3GB1b8qOWiEb
+U7JYqVrGa5o5WeEr0J3Ne41O0YJToA4rQxtVghWbfhl23V2roZ++oNUjPSIc02i/HwNE+V5WCWj
WwBIC6x8FDKrbhJcmHB3w5X42cQjcAsaQm1es0urYM170Qf0rfwuw4CIksp+v8Low91B3G6DwYGz
wlgXJhNAk+TIz4N/Wb+7OzFI5U6SlVgllE7qpk4G6UzMYprCiDik5hc8seRdsTcY4jU49QhGQ567
tovD2dUCfd71kh5GJJMp659B66Zr0mOyw2v1im5AoULY/ANeSwcpuP3PQ7CKjj3XPeKR7/BkcFXA
oQvRVXIa8j77NJaj8B2TbjcK7HeSS104b+hHPhvOw5iayVn1g+5DF0sNqyCYPPktEquVGg/lVXmI
zevi9r7OPQvnFkwsBZVKT6Y2U81HBWyRe0nKT8qPuDYobg7iaztP+LUVQ4soQbAl8hyV8OmCyWqG
iSwXRf6GAYyLU3X0ubiBemljAClTPUgflhrtxYG0hZBU+55xrHzZYl3Z6WEAzCllEtXe9En45yQc
Wn733uES8oj/PSnIdfQ+ovy4D8XPQp2VkF9yT/rGEeChkkhoc15APLyPrCmFQD14mr2VodAOfwMc
2iMB0uzfxIeyMPwJ80CE1Vs2VC1h6O/BJKtqyTMF6Oj7ybCgM+hRmAMScoMD4tYVkTpPiSvgrmFi
nsaT3CNLs53aWTw58sXZAViFZcWYSyywPGK6eMhWL+FbtH32GlU6tnbEDBA5QZF7zV2L6c+4nxXS
n+X6GoUwleLe/HyW5wvVSDuk2OkU10YPXIOQ09PFmxraVk0+lqGZvO2iL1WPnSPnNuQLLEFmBoIR
6umpbTwORO7xFCDcTdcmERili0oWJDllS/KsbiqTrDIjoCkZt7BeaQ0qZRJaRvZdFnpNoHzxFULu
Xdr93ZlQLI49Wi53gq+jLWCAXqHsDc4D+5dxUrTnxfNoGLcdSNOioE26zLVa6eh7mDsN06NS1fOj
JkL6xsXch/vZxeO1llcyvB/A5x32bMe2a50zYe0cMvMz7AWaQriLwpJ61WZdeHqKu6gUT2LQlI9S
6ZKrInTBEaCZCSoI6wzfd2HpT3i+/txAkofqG7vdi35l7ULJCqNBEYRujhwWKFVwGoXB315+U9Ux
IU02PdD8OfOLWWKVRYZer77cs/GZrO8/eE9+Huj0p3uBEm4ahZzJiEh0nTTF0HTVUZWpKanxlZdz
QVWA51gwzxNC6hIWqMVlDBKo3+zpTxPDqpPQY7FD6dWWfMgKMRREosA42LA2KT29QESeVSMLzsFO
EIrlbjAqaW64kteSdmLEzqhBtPMLciXPR7EQQOL4s4CIaPSNLpjO7e4BGl/UQ7KA5MZs+Ev0ZWa+
DFClRrHucPTCqWg1D9fbKORjGCsBEkKvsrq0LBOTXj7MuCYVDxVFVcGdNqojqINoxVoknoQJn22V
ypw9A2d3CUwNjafCm1BO/DRrfqRESWS2sWdzDgSIW1DPQYloCBnrjhseww6inbtYsO12wsu7x4NM
xuWyUqMd+wYoXVnVUyZed/P+Dje8kTH5vunYn1UQU5yDuVy32RHf/NNert3L3HlMipg1ZJKtmBkf
Nq7P+3fhYxhFgUVACPECI1CugWS3gNDsp5eBDwNqmfNDzsNWUTbjCk4jJ7/rwmr35l+5FxQXVrcV
txSDrVOVOLrZSclTq656SvzHH1MbG1fRgJ1WODiacB3stmMp/lJ1PmprelaRXVdBRHRc4/XE+yo0
pT3SL2LRU8BNepbfCW+93SPzc9/L29TX25l/TRDVLo+LwkrUymmW2sgketcdQB513WHkniKF0xTK
MH7v4+cmnzR9duKNlCHLPiIZIr4Wa0U/klhdvC5QmpmyfnrcHlQ1SgiKYvYj0xNaepf2LZea/igW
md3YZhKMNjqu4oXSpLyzASHYrjS+TLj+bqCaAsm8wlD5dnGyezibY1bH+5QlVAxdagDTX3lv7Xp8
BagNt1H9qk37Pg9VLLJq48LDpGfIHmDwkXOLkQFSNLh7vJQ1c8wzV6vgcXnqNxhHKmcYWK3B2mXM
hcJEQwwRCf5qxT2jW+GhZRL+O+2FDGVdLka+m1z64vEHkm/XmxwZqw77Fb8TpdFwrBUEZoR4kfEb
X+a7OUunsVn+S9413Dem6FIJS9iy+Om1t35sqQh+yYumC+EToZAFoGxjHQzY/Ct5F89PbqzTLwgR
Z/yz7e30vCV+Z4Y9sG1KaTqqq5U5eN3k6D7fN40dKgyLEwZJ/+BMhxWro1XT/k/CoEpxXxVibHCn
uw0ln5hvwoY4jnDvghZY9twME3Tw0nAuS6EzkS+Qxyg9hxbjU8JggDZ5BfXl/+2c/ghLoPY88plO
r5Ars7JCjSykw1OZyFcYPMn5CFS6/KNoeS6YzTy2UTT0hMxDUpjytwAP+U332/wnRXETPgP8Fr5f
oqYNo1pq7xDv20LAHK0TdHvIyRvTAwHcWtnyVwy+3knoAOnAdDxauQjP+Z94ufUQk7UxWX5bqnJC
+0N+tLxleEKqO4ETrN9Pns01DTdD5wBFBfWVkXU2d+0dux+FLhCjI4KdobkupPBxLjVTgptqtZeV
pOguDcOVaJtpT23mMgPBGEvopeo3PVRX+J7OKF9Kaob4MDzrxm6cjUySm7YavWGMUrcPSIJ6qjp+
aQVlhfgyYh4JhmEEs+i9xdpPW4lzAU3m8xqTMWvT0LX/CRWvWHc8LVgV5HfsKT67COuZ4N4kZW9H
9CwAxa3qVrYv5Btzfk5nNQauuta0ujIGaEndgWBmEabzeCNCu1FestjnxT2uNRbCXC+0o5QwYfYx
EUf3xysSjl6K0F/V1Gb0DZczGcOLnY/GpDrXYy3bYIRO5GMRIF2rTIRQMnB94q3ZIVSvQsMv6/tA
stpIQNaLfDDLUSgecaUACMzov6kBWPa1+yTqvXKfczqr48zzvhiIPNE9VeY2/uibeQ7pL0r2qIqY
I4DvdfHq3r1HmmcTUJqTT4dTa+hIEgTGRIdOGYXimEXOqieiIkvtDP7AQk1Nzj4JP7HIskjVrxtK
K4MjfX+inEV5R5mlN74hnDxDLIodt4w8R1y7s3Rq82SRvgeUtpShqG/l9wZACYYfYjIu73MmRyqf
pEOLU+JpJrLH/hQHxqMsNC33yitQyUiCt/ioXwl/myvytfQWgx4gPwc8UWjHAO1d3wYDUYOdmDdu
rLouauWt87f9+WDuLrrFQgX7Ff/MJanCHGu40I7cpowt+PdWDl6STF3UyKzq9D/9RTF1Xi1c3ArA
TUvXIwa6hZ+5hKYrfZObEkxGTfe/g8bP/jCcB9cJVfk3JRuuMFSzT2NqWZypfgqkJLu47kPeYWXh
vep6iCvmE4rawDHBE6s4m3Eb7TEe2SmnoAgMZTkkkl+NGbSqRTuVv8tf6Ne59B+8/mvP/vRyMElb
4qR4w8CFQAjL44bwAY01kmRzVz7LGk0EgMME3hnpxM7oLnLQ5jeQt2etwGrK+cmScN4HfDrN5gjR
BBZCHb01EXd+mSVw2Ztg5j487xLroZDyU21fmSn2TKcDNnKgkvkfazeILKDtzCM2QHpltrtoQYFY
EN7cIwe8/v9WiMiRcvD6F7JotrsE8JDM9Mf3c5K5K2F42CSp7tJHJOevEUaGuCczk3E9BiQgBOfv
kDp/AMrIQWhCCWvs2oGQA4AQ+snN4wRzWt8LGpL1qsVL1seMvXOEsM71Cef7JPeCVMULmMEl/87R
B1/mQCK0Vf/shcDLaJOHkkmITrEy5pNamZrI0sJGGQU9Hcer3rjCc1R8A/jpF+95FPHvv92UhDh9
J83t0nrOkEzqsOEppAmaHOxljLMaYeNPBAqz3059bvngbsQjLINM9qv4WzFYHsLk4FD8/oC5ekW2
1tSthYxFhCp5DJYt312I0uNxk13si5KnXuclAz0sUNWUPh4O4R14hLQEQ/SK62Qt5dkUkK/uz5lx
48GcvBksA4KaFJ/NGxjkmiqjbaLl8ofu9aCydKN2SqtIKl6OBpf7j0xCJqj8NMShYt9k7fVRUn2h
0aeBRl2uSqZHoiIrQI4lJjzZUabmPDuCpo50ionMtHBOqU/RZv4xqa7Wu41cuVNyKTRwYns8HkbO
INkNJtQLLCqy1bCWtbD+cgQiBwvvlwrv/msHo0AAJDQl6uHu8jXW6Bju3b5yf/U5eo347Qungkbf
knG3Qh0nsGQdpxZfO3N9g8sZrmZie8+/Ovn//lkzvYg2Vk0o4WOilQyFjIo1q8Zch7JEPwxEoKea
BlHQzWq3MtRBl/l4R5UHPy6jXksjTkT0Z6Op5LDC0r4x0DJen/amGPtm5yQhehmmUElpUQKdRu4W
0xifms5re76q66s55ookGlnbv6FF6+s9EimmZw6kRxAquiRy0vwsyFLm0qmfFU2FmxvKMFs5ai+5
GNd+oYHEg9dfr9zXKmyiuGK89RpeEVLsGPT8Q8Jw5xayGz0lHiFVQnfHMX2zPkPuP4/6eSIH8ek7
1A9obZPlV5mKl55UsfKZpvjn6WKyyjMv6dZHoZvbupvslUA7AFSEjzvUXN+tYGBpJ8yi9iFqXikw
CPLxiIsIE/gAyMSSiqk+GiiSiow64wqHlugyQJbC/pQ18AU74cxBwhFSDo8vxbbLLU+KoEsb7y9+
9wq3jxtY1VZkIsxOrFso7p5f0215Hi73SPsDf8KGwMbHnjslI2wyJQAld5wC21NdJKYBBjEIR28X
QMn08xaqR7nPB3CqFCc1hZACkTDCXK4gunoZx+GuWrECxZ0/IVw0ncb/jBz9Ar+cyg/rrqkQjZhN
2VnAhIOQT7xcriZwf4jQF67l282JIhIALhllpuTtInB/YFbxF7hDG662N7tSZN91VjngSSErHLQ/
DQOqL6wWljIoxrxfkWs9W9BzuI1V9qdNwVqO/yVs5TfWl3uQepucpKEJegl65y9cB3A2s77j08QJ
G/f8MIFhV0rV88JHHDgFKYKLNiSPoPdI5dnzNESEV/aEwyVbSxQ6U56Hq5KFFbjRm1mZdGE5IC51
M6yD0NvhCcxSdybvJL2fbyKmAp0a4ScZp1x+WiVYi/RyxLPbSe4NUhN8QrxhLJj4AfDhtpTDMSTI
5R/4T5ww0T1/PRJHqCXqSiqP4ss4832KwNydU1HxNTpjOEjWcSVMrZMc1TgcPT5jVqI1klKyEYHX
BzBojhG0twcFlJ/hmiJ8a4MLI5dG1ceIWzwJMfPOvhtFKeZaHnxGt35w9awIfPh6+wEH8IJ6r7Lh
uSBv9VeZ1zWyLP1A2cGI5Za2YGF1elnYM6TtmjQHSdjJvL6M9LoclpeTbE4htHx1ZPGLxwI2b0r5
SurVKYNWP528yn0NOv/fDgtsz6J9QrkaZUMx/FUNtR+IShS+lQFuDyZNzxRoW+Qs8PG2J3a/ebxG
weJ0FFq0010gQkDAHvZmq5w9Zh3DNB6AVyzId8S7+WX+nwcht1EFVXR7+npdy+Oa7MUak5zPf8xT
7q5qc9aQmu9SAEMMRnwkiHI2GMwZkP5IuuEjrWNvVlTg9Pjh5L1pdAlwmy+oudoG4r2I9Xa3fcJg
H4mGnJj3IKUYtle6pmUo7TEjtEpW3wmDoJUVHu+stzvYyqkS0P06pPuIhZMAoU5fNrMwH/lyCwY3
IYyj0+TPN/sGBXAOA/QmJxTIyphBuI4IOYjBhqOwn5hNYTSKCfeYwvN5r95YcIsYR4+vDTXCx98E
ItvFouWQS1MVirWngtWBXixy/Df5H4/P3WITQ+L0YG3zX9uOMFDo3VjSbpLv2Aj7TMpqZfj5imsM
DZEAkOnq/311+1ZBEcLDpGRNO6gkzB+HcLyzIl0ZzSlDfZ1WlqWA0OLYqOcdl6ZiwFrmxMLWUHo3
IdErtov9bIyBUCKCfn50tbNkXDplEbbN/pX/gaiWI9JNjWLb2M5V44tk+nZSD/chC0ahjKhGBr53
FoSKel5XNJN9avgNK+NHXjWCPMFAsfAry7nreFLxHReD/td2gfT8C9ERp/bOqhRZfkWrnmez1IVr
mYIaPAfH8qyDy5ArApPhMltMLek355Be6BKoPeMJKFE0ZlqM1MOZ6xNy5vO9t5zepfOYmwvtNcmE
mXA/KTetbtGYUQHUaFaCVuvsWX1TbxUU2vuf6SriUIyZ3qooEyiN7FKEWKvSA6ySYT/enR3gNXcL
MegwI1eO994aFCNnqutb0eesdRZLLUmFCQ4jgpj/IOSS7CCznUw78154OFRf04aF5kuPhKiEOtMp
kXPEoz7ecZ6SigbDI21f6/+aqed/mxSWxIfJXG4waOW7k/EC0bK3Kd3jTmyf7P5nYcQO6g7ME8QB
GuNOZWcsrE1HYrU7Qp7l5XVFFMcKDIBGrBq66yR3uhYMUHrKAs2vtHgXmdLm7mEUkdoXpDBvstCV
MfxQualXHUUp2ZxULtuGxh/uOMAHR4vgk8MAXIRfjIgABGBVQRcLBLccJ9Pfwct/Gc2wNCr5G64b
H0M922zFN7T7tqn+GMQjH7FBvQ62MJAx5oJdmFffFg4wQ4Jxh5e57GYt/HHYzbBfvrfGsedeOIQX
hZ22zcSwuCcDDeNyiZM6jUEp5HCVwR83uz7ioe9zXKx6xzDQb2ersMPHedUV77VZBMFEvNhmWBWr
eiZK3bi64DldVMx6JBQzHTUE983HPwE0ZtZyeT0ZOCARTikCDODNiUlOenD6vuSWU7lumvzvCJv5
sK5xIZa4gT1U7VEi1P0PfoLRxNx2ADTTWCXgpfTAA0OFuPEjfo297AqMXi9jDaZxDeXMzU/mSu4+
2HNbuonKHZgjwCNetesDoiVgkN+Ztj5R4nqzJFS7EgGVuJtxEaQM0hTPC/W7jLg4OCJO6+RMMOsa
jj6pRVowy1Zir9rRkphj/7Gln94f2eCPnp+A86OVXfjkoEcmcK1v0hoWeT9SCpRkxpXWBG5cadgI
tTyUDYbbBDbWki8xAinKtbvXJPWm7I6pcpW2fKCJUxtVf1wtJEwQwifoG/G5GPKUdH7T8lGUmmQJ
1ieaj74dIBu9gv8sn2SDTwbelWdRj4h/vobwWScc9xTrF/jGbyfy1cEf637grmHMqhpg0liDuXIJ
RtnOpqgP8o8tp4vzpyZZ3XFJNJm5WAkEBFgHtSBlwMBMBbwkYE7gX93oXxvnRd5fMI8+FJfpr0uM
VpIFkJfZALHIiNtMl+pOPgIU42KGF8KEgD25XSjSBGkSRf4lxxbT8lXkESKoNknp3y/n47acjobo
WzjMuGg5wTYQK8LreojTLE+ftP4qtmWEXNmXfrY7ex5sR73YHy1mu7MHliXERu9lG8KpK/WHDKRE
IIgenxOTQlnNPgZCIiNWiEIuv1CUox99yPA1fDpZ3pTWoolhk6Wq6MM3xIdmceeSk6kWr0rLnMn+
OIAHbaZJt+mJmODzOWJR7XvTG4s4MMhM49ppBUQGxLXZmtca/Gvm7wr1b7cux6QBia606OyQamXZ
itZcdAxoGAIBxeVu3qGUa0UtPS3C2lq59BwFmUwCQjCzJ6Ce3QjaHvTXhPlwIloYUWHtxG36i/cV
/qF2dhvrsmFkC2K5JxpD/2icn/veAHxnRlLU9CFzEL9N8S/NKeQTM1MwAfdMcUIpUhjLoDq4e/33
KOJcn3f9Sz+IwSkIOO1Ykux5fEIuWoM5WcpsigajNb8RYT9f0PTrA80kA1ytWMHfeb+DeobH2URU
C/W12K21YJSFdRKs2CJ7skC1o5iVl/OIpjRVRTOvLG4jEwWU1B8Ss2EoNl3UQjR5Bm5f0S0KX+9k
tS3jSiYAipRxCc3lQcLxcay7TPKLJWZqnX3CQE2fG/xQ1tsHtnVvvY+OTGvthyqgj2r/ehbzbwnT
tRliAiXgynsN7+vCvbjMaRt+GOdiBIVRdmcsARn4+gNQPnZ9i7jkEUfOQJ1oMG/HRW4eUiHR8/Iv
cZdci25yWGmLr/GlYlp6+jmrIExw3r7wigyW9936Lz0xAH8IMGccFcBAAcxyxAmR0ztgTKT4hQNX
kAYYQU/OZ+J/QGivwrKklAXWnvu403y570JaSDcOUEKO/QVWBvgfk/sVLBNFaxTPoMM1+uKYBaw5
2kpLGIaDXsENRRvHtzZYVj1I8la/iL/Q+8KySP35wS4ZH1VRMbxbB8sej9b8oaphDH81U1NDBT3T
DXWgllkN8hAn6HvAxqlCimlbX3B3W1X5S3tdD+3neCEOCKrKcBlZFIt+qmqpnH0dbZXij4vPYFHd
OuIXXg5fmPF9LQHA7tWn4K3ez84CYPLViPJwUm2rhWbfgzW984H/7gxz1QzjgqDSlNffftqx1ZmB
ETCd/t/Ncrw0/+9A8297SlVyDzZV5Cf5cmg4yG/2060f5P0u6HrtUe/NWyPeqx+lZyw3EE0nlWlS
JCJbc3sJHhLIFqnVN+mpN0b6aNCsyGzeae4INEnMDU+OMZHbfkHIAtILD6UR5RNBAGxtNsQVwRzn
5KM0+ivf2DRVYD64pFONfMayz4Ud+XqbwtEmkV1COLLtByrghTKchK+8HfN15x6wPUVyoUbP/Cdq
7adgV5+MiNVxv/9y024rphX22hwVM0AA2FzVVJGztTgn16+XyTalPEadxCq31UkRKXnxB993j2fk
lpasa9Z3RzVxA9bWGUW/l8FF1BOtzKB64MNlLQly243bTla92rY2lRe3l7tMQbRE+bm38GKuAN0J
kcuhsKpWB0enr2j89cFfbqMRhILtQ7zE1RXNCkixR4Rmd4lrOwg4wfhdy5XP+3ITon/w1YhwEUED
DzvH+dxNPARX6Hkqv4rq8ogoDB5++gNlhmhJ4t9GiK+n8M7SyJpn0Y+O8AG3bkxuSfiT7mOBcP9Q
P1ucS5MV/OcB1hUsznk+Iik++VBZ3ZIY234PjGDAPlui8AVuM7lG+cHMglsv/W5Tp3FdypCpY/6X
ANG2r+/C6IwwXkov9CsfFj5yb/NkOvkbnjKHwMzz/9cwdcGQSQJcmCqcn7AKEtPf7W1yGoYhNW+n
AxHmXfJBCwD+jenkQoe9U/BcS8JPEmMFgQ5pxtZc9zDn5uXkVymk4GoRSJCb+kqXfqtnQfcYWvEp
xClvUD3wZNB0kZjcZQpmPy4zPjYB+kEIzcnRHPNv17rdWvP6NAUj2PNhShIxh8zEojkvuGsvE7l3
eZMXYsdMtpAQ3JNgTvEnCbV8lbaoiHa22ivsTj5lQURwQPAJf6GlReonwPgz83ajP1/nIYRDv5Vf
O/3ENa2knxCR9V4+cRCb6ujqItcW84iAAxW0iwOLA6N3VWYMCPFeOEF/mzEa/GPBLNUNo8zHXMxM
0/H6UA7xbdzdbxMKakx15CzJVimJHv2vqwCgQlR0Bi+/x5vLqRBvc+/65NHdIYrpjCA8i7UGQC+Z
CgKQS4+XsZxdtp0DUZ5nCrTarkMCTTaE7JGKJhbVqZwb0zPJcjQiI4/M8kKgS9XmnlEWVB/prqqj
ifZwHHjT2EU6s9kegoSeXr3bIa/Im0/xcFD0eHyp5PCJ9CpJ9H7Gkw6tU7BIpmxYcCw/Xs+ghbt7
01VsV2eE7cr6yOhLkegV3snKm9X/SIcFgOMpRjuqFymRsO3Xd8ov4PIgdPKUIboa7FqmLqOIUFmu
vVeZh58i0pz5DaIp0JJ4GU9YywZXUFARKDhdrp+Nlelq1sMeryiDCCNqIw/UHytqhqgojMZowvHh
u8ydAMxOY21kFe61oQmqLeoTjWyscuY5JeyCuyZdaYzZNrVEptsALTBO4+IWnJ4uN/teghJc52uT
MYI9QhL8oqLIf70UnYymmgeqdwAjtr2Ofirxj0sTaVZvkYu1wyMTstp/FdvngiEd5T/mipvQ+7r9
JYMadrXtxiDdppHvoE3WCBxVkI/U+VBn7etzo0Z8+RefI0Z6UaGmq6WSjJyUnakKFnuN6ifgg1Yf
ZIy7UVWeI9yb8B5leivtuwufAxrMmHyN0Mu0Z78LezyaLkGyFL6zI5jhOAy8oA/BVHgXzdJnI4xG
LhOW5cn5xsf74znhTn+/AlF0gYnvtDCxYFTisCT00nrJDk68weoRbV85NGCPhhQ0fwIDD5WrG5HI
9v1p5JTT+ndok/ipJyfJC4I1n2+jdaUOue02jFV5ZpJIS1rbhoJuZhT4KSTFnF5nzlMbU/xj2YeI
recxU5NClXpsPRTccglw3lX2lRqNjICj3vwmUmPXwukSHSG6fgP8HFTCwKGDXIYBHjWr+kxWWN2y
xvJ9k/fLxTzoK7N4s2d2ErpituDxjzoe9XlBWzzCcLO+UfMrehVW1NnGmUE3aShUEW0CCsvmOqoC
xC8NhrhFq82NC88XjTWd2pJamEwFWJjZ5khYKjnstgTwvqQKmBtZoVet5n33Ix5egUzCNNucKmOi
WFTLBZsBhxRjsz5BAGjhgba/oPo6Kj26QwL8hdK94eEpfgo1TXEGDXhMhjZsPzh5Cr4cA6cDgq9O
3Dq7OS5qMmVA6rQSd7NAJvg/jrNC/d2MXP6GA5uBjlTKi/OL6cJmwC3dNsUBRNhH5s548SoYzleK
bxPfrGy0vQm57DhU3ryXdwfW0gRNAiMXBz69ToQnTB3JhOpro5NjFq1RCcF6XRKw97OizdPMuQwe
u0V3QO7pqGv2oC2jKgH2dH+CYqol2fslgfzSzqVXEC91nvDa1NZPll2HYujuwOXiKmAu9HKCgbZY
8dIMCUVxYI3FFPzI/SH0b1qfV2tfYxjz1qT1fxJXFcMKSEmdut2ZsvgE+M/zbB/8rENkNXmrj7lc
X+TA2fY0l65o6vaWhXQo9UiadzwOwPh1spknZ9+CpTpanwEkXw0fYezfcskL3VtYIPJ5mr+R/87s
ajPFuglFHFdqdiBK3CZshP2m9j7NWBl6cx9zP51OOo3iFDoyiwA+ywLerPXxkQ1zkDuWET2neCbG
/J9/svndipBpHZVPE/Uz7FlwnVFdOUaKYe3JpIerB+oStMgtUluT4Kwv94R58JXpbCRVbfRHoezh
84YJ2XFeca/TpEKZBWA9YwDXuTVMiKxLbZoACY6VyDhqrIzD3+ymUk6cASz6canMnEcV2DMRIfLv
bv8ROnAi9gq4LIz4dUyKDKBlAfWnsvqdFQ2RAOaH1I7lJe2zwLuJj86hIlJRiMF2Hbqi43WlE49E
8PlZOswfxRPB6PL0/wJu3PKTWu8cGOEk8BGFq9zCLQFjASprWPxg828F4nPcA0lG6FLsqQd/ENl9
yTOoYTzqzmNbf7bsuCf7V1UcHgVVu1HaaKqKk6PfWNoBvJnm8cmI8rcGF4BfgENBeHFzf20Chh6N
IAzXm/3+sYrI1N3HXhxq2U/YvZ0Cb+b66dFSymNBNHv+XF0/nQPWkVhVTC2frv3QatJpf3bYy9LZ
vHvWGybR+LzWr0cqAXSRarWVRtk+WLB8Y+RuyHHkqiKGmU1y0jvhPxm+SxHPLelwX7AmGLnPaG9P
XE0FhPQvD8OgNsAdtdLonBg8kGAyu1cLly+4ydmaHEzz+eMX0jg4TYI66kyPq3S9oxEsPYuOoMGm
crL04OZLHIG3aeMxTuBTPzVbQddV1+6eSkrjbOKKnlktcAOPYGslUIIPBIYUmMRIc/tldQoRMNTO
zUWy9ImrQRYvysDbfFN9BhtPMwYCfzYcV6pWWbd/Andvi+1EOIJ+4Lq1xrSFXHiB5L22YmfD1U9s
xShdgvEk1reflibuoJ+0LeJ2hyPFotEZKDFUsA2U6MFIUbgXCyWUcl71esvS9xWL7qD8d3ey1SD+
gItSPte+aoDPE4gHPpSbrMQ9g/YW1IHbTevrW75uXrHdF39F1nIffiHdF6bCTYv9ELklLG0/v7nf
rkMm7qrtLCoq9g2TcWQKWzZ0vqOsMB49+1wGhF0CgEbVkI0QJVBOw9IjO7QR4hV7vjX60HCt+nUF
UHNlwBTAFvZBfRD/qWVQSSd3tbdweKv0NSfZHVkWEMlTebg2W0w9MrXth3iQNUaOfVQakfS0SthQ
A8WqgjFqYmhnSE4IvpnpMsya4sMCjrTBNTmOahdoDvKfG/3Nm68LxO5snzqmpEfGQg0jteyBaknu
XzLQSQ4flG/E2K+m1OuNtsYth0mheA8lk1il6y3KEmgHTBEd1HqpEs/AbxbAAD27tkhcsPcnN+bW
OKdAqqjZlHwnVonhqxwzdO6FKk1qPC67fP661XVT0Cj/fYpQmHsJIZ+dUh++GHavs4AKgBtHZOdV
DYo29PXNYWGlJo9AaHYDqZAAUsZrdgbSdQiaiOwnrjGUfbFK9zrqdxLcu7OCIW1iAwH5ydngOyGA
1OMC62yGu+11lrdzkiPJU1yoXsxti72x/seSgl1ERMWoLm5Jcwc0pVKdYRq+IkOOu2VGr7cc8SjH
5O+sxm6CWV8lrAyh6HprQU8MN+XWJZd1BT0lDfDdYBnI6sMS51bPYhZ76v9XbnwfirgsLC1Bv86m
ZxgNrHVb7HlL4kx2X54NKQQgjtyDOIcg1FC6Gl0pK9ozR3mUzL4guwCHei97IBP8xv6ZNDpooRf/
+tSul48IXuW23pHkTN4V1ow1LIHq5JHwfiPIpzpTAZ5oDcFontKox2JAruqO+2wtzHz0Mar/VkTO
eHLB+hn4AVP6nru3mATKIOhwCBHejjauoXFXvOpDn4WMpxPZx84Ye23uubarjPede8MSzUzaCbDo
DtINWxmB4iUowtpWZA4u5onhtUCZYimwzEOhB7fAvjXSDPUSkPQuFTd2vo7sVVISXAbaDEjvMpf2
x5hJ6rdT4LfLRLJKCBiAtaFVyA6kAIYWy+DocvgXXmIklGlNveRDwX4G8IhMo3mkSguyGyyr+JVt
gV4OMqtYyJh0YMVr3nsMqWoKnIpvWxvcI+fCNDoVoPgXnboMTAniSijDE3pMBji8EB6dRzKGJR0j
RIyBeUQnXLRCshzMaqcz1Lxv12VJzd6tfkin+dkVFeMPlqpjxQXlxuN4aYft/vT4+zWyXNVP2GOg
jHUpR5Rj6rjhM6pcF2k4k44FufxqplQgmpFT5WKE6Abeq8LXrxgcr4NJRbEKJFVLB4nkFSQfrMzV
HO6relIzrgYjlCfPegxkKOVCTDWtUBfb5RZjO0kxBLN2BCyyJidYQMX3ESx5cqYRfQI8jSWbVtov
q7IARq0qZxu/DeTTPksqrHfON2a4L8WaQi7qlgR0BteiZG00Ow1RlVMjo5T2Zkl+2HjkIwxM0jO2
43mAZXRgySXdyqTFzdVdOp6T7GYCZXkY0s1jiwgvo1RNAG74QNeLOZWQFad6TIqefa1eBf3PEKdu
7hEre3tf+rOrYfWt7dkw7It3QKjSBI7VoQ7kASEq3PeqJBbpT0xFEeCkrEevMeihaeHvhxlo0Oow
jWijXzBzrlK/vc+ijTVAPHgYFIaH5RkzEvU2XSZlXVh5E+XgXVPiFd560+w5spiN2OZ+fQVK4O0e
cllBA5v873YAZAgor+gVy8EKjUoziP7MAfsPWs/A8JW/4V/uUUaXBHT/l6+s+6t+A/hLrFZFIL5b
NkoMj/TWfxonWo27TD43TVa9oEkDCfU/TQRT3jJjdZdbdT5LQ99/LqLbj8jSZ84DQOmlYiWp7onh
spKcBiZZIX6nykCa3A+P9EZn2ATkdnQWUoc6e+pKsFK6xZ0VKH+04lc4QdtwKF9NbLtVUdoG1qrL
Pf9Cyx8wcFhZPMgLzpEiia0Fs8lYRzy50Zfz3O7SW6YmK1sI00PMSxYE/S9TIDza0HQCeQpNNMZW
BBy0PSOHCFFX3dpKZ1VVozHSB/n0fTjTS+8otUjzFSv1altScOfMO3RZw9X6dNA7t3+nWDjCJ6OD
zul+ltNRQyuzuQe0srrcUXeBjsSrv6eg1yMN0RCEr0ozyvUuqeb5uCWyYTka2CfInWEbW1kN6aQg
hj+LKvN+W+yno/xUNBFvEhQJAdJfhEN0rMVxGx1jD6kIklz+9m7NueAYMWMJ5TpUiBpfr1NktsOX
VS5Um7B0x+eEPUXIhtM76/CiF/0YPnHO3Hh5aamXNFhY/DyN46msiz6a10weo7Gh4mq7clzhBiEj
a85smAqhuHm7KjTQ0K0Nu7hR2tNJUVDDzaatHCXJMFUfgNAGvA90tm/VwWQpoqI/IDYz/2naTxI0
eUCHLObsHwvqbcCgWXbPLuRAWGiOsn5NT7/Cdi/X+6Hn8uZLXkOEuWTbMf6cavT9jLbEtux5jz96
1mfwkfowwEq/rUnzyyiQKmXehw0qNJVXiKEsXANeoGcDcQEU96BUHmx8d5UyY/qdQSsieh13Jhv/
zChdnAnylQ5XpGr5Qtrcc/FNXCQZcTthRI+LjgeEqPJni8OvfqYx41cCyCh/ptp2HHbxsWqQLf1e
awtctzSI/iT+Xc2BFVzC9k07n/SePJJiz6Fqz/i6OuJBv1ewRPhS6Ng4lFWu3rGw1OhokuLiytbi
htyXxJvmpID0ZTlTsNvTGaMyrE/tYSv19qTOwSWJqjg/lupomeiYhgAUjSBMrVkOpcyuxT0pDfeX
BD9O3PTEWRUhz19Xy7nQKaZDPMkNxoWCtD5tiDq8uwDz5fiBsYna8DWjVgZNlP3aboFh5vNesBri
u5fUgU7wA8d+ThiGnO8WD+nwDC6zrOxsy5A0F4+6INS1AH+kHehonXr7VcJAEiLTcyVkJJTdM86P
+k/UiT2m1E3j8kPlBcUGGp+GJA1p6/7f2AkZdpA1ZN0jJC5VMVpfrA9FO7sKCme0qfolNKUd8VuR
hrZyhnwi3IPvaj7DmdLCb/GzbKfgWHn51CaChJoH6cNob5RCGSwq3NcasZEAH32hka3y/GM/IwKK
uDyVXNhtMPPR/4E+UaJvE37nVhYiq6gCZmifPhZe/MsbIrli4wVHC6IQ7JoYhKc6t8x86nXLnK8C
11bXB2ew27agbbhfYF555S1jX7GpH/cltyoyhQL4pwT/KhTfVlmN8aZjbNjPHBh4lANQWvnADA1e
YShh7BWcLxTmRFvFkkTmzNjdbevzE6SfOu1+wmrGnEwKIGMepWvx/YE9TCHeEFsrTY5kBvCkXTf3
x9ju06wUJ1ADvsmUX8/k0hD+URGGZnwzHBRcBHhJb7piI81YGQgw1sIVkFyW2YVkI4PeSydVh/FX
MUqhJQadkKQZUNtqrVA8XE34Dv2GWmwP0q+4gHuPbObWscjutzQ7zUHXXtUNirMbnah8wxTPZR95
xQ+P4ZCPieeTRCcCZ5SVtOY9mP00If6l4xCNZb2NvZXkAsyETVctyrBOA56JodedDkF6ZNiX7MGB
F4N8he2FG3qUumQzZibCdoVH1W8pqjZdCcrggpifngzL7heewe0svALCobrsKrObRorx9H2FuK1v
ISfvyTzV9YNthjml404c4yoqbE1hYUW8DDOYNthTJ0wMMw4WrV6Up+3X7I9FhfQBrX2ha3+ciyw1
QyLxzsZwgRLpP7llU0ban9Co9kyqrP1Dnv7Qkq1su/HcuiJuRqubccwfIfJUhfdl+8dQ94FZmPE+
IXPwPe/dNxq1NLjwrNaQ1nZiS0DK/mumyR4WM6ynXodGrRUVOxWrE4avkQ2BjSFUy/u3jnt2FLXB
3j13Pk+TkdDbwjHfRnDnepCICWyBiprkfhNhESRE0Tw52TdO14meeftuGsnuGQzAckhdowxiICwH
32GDilqZGhEMyoeucAC6slqS/B4r/4FPy7WQiEqu+sJaxS3nWwjhg+9GO1J9dlnSvGfvnwj2SQzw
AP9rq2lEoxyO+YNftVRBDgbF/OGQGcaVVjpnCuWqmrikbss0PPssfRDxjhbZjSRDslOvHIgf95vf
dDNYrq0yOjSIJF6Pg2+26l42p9fBee4Q8WutGi39FhmvUhRQJOJ1hM1LprJuxpAxIYvHWB79J+0/
fRIxbjASR+/OFxPrezoan6/jOL9fbdWR3bGEUvCoYWWQY4ikjpKALR5lWcoNjqrKBFC+/S08C4XZ
okNjcnTaxCLOQDX1ngfBgU1oZXEYWxhA5StRmZmfG9XblqYCGEol0XUElgI/7DXBDKnt9oKDCvyj
G9uGTLNkGfcDjh44KLmo9DZUCK2HzzJjpuQvyQlKNHB5ewAwdJa4znnC9DuzPuMhV8TJb/3d2GVc
a74f/9bqBZ6gsYby3aadWlzLXkqgT6ImeVNd+bJn3nqFeHD1oPOySxgVp3VDsVGUjGJ40LaPRsq2
dAnJpfiN8tcEcUiyxB2yQGLI9Nh3FVv1//3e6Jgf6LOrcG0zfQi6eocF/yqPWpVwlP+0me73rmWv
g4DuObx/Cq/rGBISxEJ/+hJ9fLacUXmvdzvNDgt+jJptG1SaVL12liod783jjrm84sAeglW0C6bT
XYmlH8ZtKcyACaLSfgkeoNXq2nJvD0keYmqoL92cLDyNKqkE8T4rGtkCxL2IDCBqcngodzSV/lQf
tY/N09kAob6X2EZg+1cKVDdrCeGJxAZJM0PhKsIypvvOmBPGACDxboPxHhXPk53jbJv5ejqEeBsG
SsaziuGGbJtkvw3X7HAUcfV7MSUAQ2nyJp65+SkGsCIsMqKTFsopVS+EaZj24Bch73r3o1ebNnZQ
djNTiGOlAkU5JQ/rryuWLBXbNZRkv+IBgmALE7rTYK0cCjv/xe7SEh2oXkvBFxIteGJJyQ3v4Ghf
j2MzibhNLJ96MudmjTx+7PFyxqEuwh7C+nQaG/AnlJj+P+MIJ6uSzE5zq0r/Q/4cGDYEbsaDA+1Z
K3Ocj0oSGXkIo6dPbQr964JiIuA/YqBtzSXIE8bHkMrR++Tp+TyN4XG2JP9Zp9/CzSYLDI4T+nP6
3XFZK1SuGVUoiElnKp95PRRzgyX+NXb9ket793M/OQ0jd0g4dG0yNEjSan8if6zCKL/XmmDJbMLI
0Zu7JMJuQfClAKSbuk7YvV/C16cKUNAv33LpLGBwQASt/TOK21OC0D8phlm6IBLzWdh4dFWhUmQ1
X3kF7CgLnuJUeCdqdYdctDdk/s3SGlcOuHDoMpa6PPnmQ972qIacN4Hs7pGdO3Mg8z/ARtCuIsif
0veI630ie4B1cMGJFDudg0dA/EOW5HGefoMafVXyzcvvzHyOtTQTEFmhv9nqBtUAisexmZhoqQK5
5jgqLUTOdX1m7XXw1AiTJoabDj6gDtJRYmegvNAu8aX1yST62FnCQISdWaxxv12wB6RZ855J3oad
LOf6qoo6Z/rNV7ODUSrXMIgoYYGz8+xSBKQEWthc4MVTP3903ZtFnfA0rJawCmu7S6zAxUtUIAy5
8fxHAoEltOpk6060jLU7LSOsn93qCUdhrYdkBpSRPmmklWNzal6evM7R9WIG+mmqtXLaeyzcWZE5
Zz/RQnClD8Zf+nwIhP9268g3Wx3XiCBMFVZlvlWTspNbTATOak4mi4uhpNCiQ7VC/F6V3XDmgvmT
8Wo1v+VJJgzKeo/6DiEvFNqh33GLODcrJapgfVLc/F2/5EsVHjsEyu3o//NKnIBm2grwME+4YlcJ
68IUESkVPkITcl5KFdyrgHhKQZn18LkYX47lw9SGIVkPT7HLNZBmWzwyZqSTWnUShAhk4e3vJ3YI
xkwoLKofdlmVd5VyfD1Lc7ZrXLgD6qA1iUyFA9XfKYN8MrV/VOTADe6+2ye2JxRbH8YE8QHiT1DF
9SPpDFuHpBAqqt3U7QVCwsbd6mi4VZdrj3anruHYNugji/2A6r6lGGMp2xoJXnjGTNry1jdH5V6Y
4RiYFxxjqGzRkk8K4ET9WdILJ58J2W4vhbDgTxyAvhYcUyrkyihh1i15MocioRCcWF4NV15zHHEZ
1n40TDa/IcyP0Rl28VPKtazACcqU3SdPMwXmBOTtkDgOovSuPNNZ+Xwtdm0FXCIq5ol6TVaWINNu
VwzP0Jq8xTRR/YV7Y1iGueOEQNptWIw4dGo8swIR3ujcdW3k0269Vf0dZMegQ4o9OEsPpa1ocPDv
oSlS0//RPE0UyKy12p5dhNUPTDb2SFNNzJ5A87da4hw9ywVU5bNNSgJw2Q42iXKSE5qTCfa0bm3P
Zz+9ts/plRWQv71688dzvnjZpnMNYhKwV3aOQTNrNYHy0haiShPP5dB+BY/xiJ7lBoFNAPeAyoRB
zSGA8zO9yrLvGqzibpCxngzuxvjMy7P46vFNzUxP2OLsZYbEU+wCkNlIsPBYkSP/fvnbVDEM1sMM
q1F51o6cnMT0VPPsSOZWtTQkYZJIeHUA748oAjIMGlq3nXsr0ANfCabGlTp+E2rrqjNx7UqwrA9u
UdXOgcuCuH5LXzr7sR+Z/v5yHnbXRqoff932nkDW44UH90Sqdxns6CoMSJlv0uJ0Bsj6cUSMUwfN
ipGDaWf/vmwO1SZMq+jPBV5C1/zdLavT8c8bayh0yl1nq+rJCPofxPIXbbgHM4YWI9CPhVnr0AEO
jR51jdQ1QHBBFWIhZ7sq2mdrn8XDcruZTvMMc0K3gpExQUHOy83teCjEuHVhwaq+LMLzGhjIJ6HI
xVp7hyQlSTiIOFy41V9+JRaIfHGxT4wzRwFgDWlq9nM+fqb9LgMdjr/VX7JOmRhActYIHOS+QdSq
IzdAKHX1P+EajzIhksXHLAhvxrAKDrhiWvTEds+sm7fa2ZKir3Dj/Se44A0J9HrNDR2Pf9vhvGeR
zppN1C9+kBNYfxLz93ns7h3z8DGlhTKW9RFoIMlZiLP+W/udP3AXXPWVEXUqwNhEOUwMecsQGVxN
pnEbH7oTUrJp7sOjxTO2IV8GtRkhEVt+qogMY0sY/rCo8Nqfrr8a2aZLYsK98Cr/vKs0PauKHy5Q
ZMmMWn8uLop9AW/2BOIwlgYFFJMfRHX9IqJnloreeJbbmYVpg/rURIhWG/cbKiUz7zFBF4qfAaPh
SA9deNYftlN5J2yoYfwgtvhFuEedDYydYXvmlZYMb5nRhcTEDyk3K3bOUzsgLpvyzrZWP45jAKk1
zE8fpPgY0NRDx3j8VUeMRiLYdbWgh8EtjtA6RS03j5mLQoQu4pAjtwBPV9518+Of2CAKt12myoNq
cbkj3YSUek+2AgpdVmMAC4XTx8PUZQ7o+FIeJaBKnbiwLQ07CyFKl41BVitGw5W9xsi0EN1zY6Sp
Ixj7i4lVsXaihV5fCZh8BcNW6bh0EzmH+2VPUdl1JwGH8gUkx9TrKJN7DT4vk3sipgL86fxsMQCM
YDt1ITVotU0rNgOskIfqkEOhYOyb5WoyhBI10rzxCdh0eM/yR64czQ/GYW2g8rWyi4OrJBSJF1Hd
q8zD8/uffLyyphQ7u0xXaJ/ZFq0WsW22gVfGdvLTdPKYSm036vUAPfCpLDjtjY3sSJN3kGyi/iyy
ChzIKEecp0URn3vFYkfxVsF42P3xXq53DPKLD9MZCkjX0PKqY7jD+XPc7qrlKlYsaPAUbtQo0YoU
ljCbNDajViwEXOu4hb8BgXmnBcPIqo6Bf6Mk1L1r2JoLiSYfjWsbyMReEgEmwOM69H5GR4TDIXQn
Y9/p1mUgEAzlPQji4oHXUTIo7hiZjVuR52O3u5LFgZol+DvOy0pcqDBMbB+mCeyJQy9/77aDE+US
xJl/YrFejp9JYNSGToqEEGFwb55q5R5lqMlM5sN7v8vNLdG2HOs0gplAmJFiQpinpjFONpQpgiFe
w16wMzt0Uy9+3phdlVnxHa4Oi9aruXFS0ssBx741clMTCQHAgknBSQGaS9RmxVVPdT2JJ/ZtAvsk
DpJZRf89+AIm5g0xBtCmkYOUpqPuTRenzvwxVShWd+hXIu8B0yb3j2+V/27T4yKq1mvCGOzRH7lK
Sq6bpzegQRpLpa8QJfYQlssTe8lZCbRkSzn1COV3lA5GNQKpp4NBPUY4hFe30OYOXP4wawUrTX34
6DPLJYK3Ta40fYA5u2jjqiJ7y6ngRdAzxuHp6oSNwVu+MYyBB7ym6eK5SXMx5rxkD78l8OAGrQK7
+Qk87G6tzLvW1KMJeXIBKZT3QkTIPRN7P3a8W3LVtnTYSAjb4OJ/d+yL+M5uQVAtNO8dWAE2NR0F
BIjo94Zq2voy2DDqGB/3TDp7r+K9414F7baCIL8LmkP43iqugbD1wxH9tPwFnYfCtalzx5bu+OSQ
n/S61opUKibGEB9hNi4q45jm8iPerQfZ6GgLsuFt+ox5YG82ydZBAipADRxR7TQeom1OB/7DFW6q
Ry41LvlJTqSqMycil7izJToJ6S2RQLTUqxeJrKpGbXffY9nIOogRSXMfZsove7ZQdUN2ZQiq4+PM
cxJHF8V8+lj88hx386eT7Cgrv77c/VVX8qeyQjBd7jN7dmNUzjIJ/GWE18vwgayUiWF60JQQ1Dhj
8CFcvTH4FURw6L3XeJV0zvzRdy/xg+cPeS4/kitWvWyjBQgxmpU4CjECczK0gRSJRYiA8BmyaZBZ
SZs5DQPvTkxlE7kepWNr1xogc66hcpHBn2UIcLzGxNyGY4vAjgsaADaOR5n050vMgCxbt8wT9E7z
3/gPBVQtNd6QGV3qBK4hCIeNclagJSUAEObYft1FPDma+mPFfhFkhS6aSaQDwXfoaI+zap7tU+Cv
sSq54U38H59HnGokh9mfAT3MkZyUkkuxFzJRpa1gTDtg52LdQlrpttFo5bvXf+3mMnRxe3kI8WC0
1Xb5MHo1kxJsmsWTCiOSq0KdnMM8CkuE4AhmDHR+GXMj8g0UuEfMJZ5bgifDX2kvDsB/N7opcs7l
b9rJQN6mU4jJCTEb0OMUNLAwgrN/UZI6c/jsffoaBR1/IuiOEPepi2eVH6QwsGdo/i3f2m+WrnRm
cbdY9aCBd1tnv1+z3y3R3oFwUCu1MYnfbyle0UB8uRvxfnUqwnNnUv75nH/bBtaBMkTDbeWW0RPv
TmEncbt4A1MsuvzZ9w5Zenud0Xp265BQW8vVD4Efdkbvm5SWrB3dMaPx0WuQnWtUgJx5yNL3AbsG
cSoE1j9PU/XlV/FCd2ZFQSQqmfMrbsd33PrAh9gA3JT1wlrkn75Y0vEYDUsttQYYcUOposbznmbD
CF7XsPQyAUnEOhLTBlToA8bdvGi0builThxB6FJDk+crIAaQOkxn2etBhCBazNqiOsQHjERzzESf
+MCvUqf/Bhfm/AexcHjPf5UGJvEi0hbDf3qGl9sPulv5JOZPGChyNk10S/pWqy/AEzOL7sdJwWt1
5DnBl5x96NkigiBQ5iaAc9VkRV9SmppMN1KYtRCYCdQIZNtCNsEBYyn6LmPT74cqGJRVKzwOyF4r
g2gU/U3GLfaHV6AGIHYPsOZ6BIAJt5L5RxB+jIEd/d3SLeGURLehBC7oEg1Ma2AlD7jSycoR2H19
xP+0KNdFGxDWbMjBmjm2z+fMJkWjNkUZGgD/T2pCtgR/DeJ1NkiPVInSmUDpewHBcLb8ZuG1XLVX
45Wa00VNNtapVM3j5JZmWuV0hPHEgz+6RUruxlWjB86pKuFMj1KL+X+eG1nZ/+IuZzMdNVBbQWmI
DIoL9QgFpvuyx+U+G/Ur/XmTcm5Y/lU9LxIWnpc6M6StN5ntagBUn8veVeA2/FJG/r3zxE/K/gHk
nYuxnoyu6eV78CiXEDqWfgTe6xDnmdvJ2jU343zuZT0BFLuwbuLBnKOzmgTeFPrpvC4Zfhr20peA
FnRYTUxDeraBRk2mWCuzFVKBr+cRRCVxfGwVlq5hUuo+GgIeez+9GbcGBmy5kEN2ofNKcRWCQK+h
xrVgpWlm+2rn6mv0DhGEHjgG9s/I/akOUUwInyIxd1oRnaxrouoRUTvHXev2hiDjniHMAsj6RiyR
IbL9V6gYtiEBB23egIxShiqrFAn8SpVLSwH4qKs480z0BM+hiDHb8uc9ekaO0V98n0U6UZ+Yh707
3iY7VZESiHu3mBqQolMwM2v/RwCwHIqCIoAumoYiVgCrBOm0rYFEoKazMDRM9rOsyAWENh0CsYC+
5krtorHzFxpbMxOVdh1k2hnU4ugqIQAZVreumzFiN46J5iozUBXkW2b9O6H0eDRHKsemnaY6jtbz
MVVcm6e4jZEoyF6tBIvMlMN1qMjkG3rHiBEGCOLRO5XOUREjjOnTFhsg043Ksgs0DL/Uqnhw+tLC
rSKTYEoVVVGLhsHHwMX36ipB3SQ3m35LsTZzmzayy57Pv4/ztTPhhNLkwQBk2+/aBqyj6lNRwsu9
TdM8FhBNcPDbqhPf6d3qcOodn9ZYG1lx6drUmTLaSXFA8aKQ5/p3aA5ue2XsDGR3/I2YaYoAjyIC
f0KSAKKVsquG+E6/VvXUTS7X5p2nB+S3MNmXzIDEOZqsLtuaKl/Y21mAZHnzB/wMu26EQcwpndDB
V+dKYhC25tA8a+kIhVPPrpnkKOnrtFAohP7Jsmp1fTa6x9tRuZyD5D2ThHD3cVIb38BfUrzv7hFh
ui0RTwjvI92zvmLm+cHn2wMBeV17gx7UW7fnajPC+6VDVICKZSgZOUt0Hg3YR2DVKAMK4QuLYaX3
eoa5c191RXzHNPwYurDFPmYyYW1imjKAFY2KT5HzY/U4i2FoAzgLM9ygZmmMgbSMzh6Kr6zlWfxC
oA0OcyZl8GZ5/kyohLL9kAoq5lCg5X6fg+meQtP60QWUvZgrrX2jK7Wy4cljZSEJgnJhFdKqxOHR
aKMHRfjd5sAMdlTxdvl1g/S6G80QVX5qkJRKdJchh8layjRmUEkDTjcDWF2wA3IceFzZ7ZJTg2nB
yHrkGI6ddY1vtG8yxpWWJxMWzwQ9Ds09wNjg+Ejm9d57SpjvkybOY45SxTQZ4ouYlVXG6PFo+Fg/
HkNJn0yeb5JNdN8lsn7uWIvOC/WSP/c8yUIhEVVKhI4kduZEmOwTpz13eBl2CeuQ2DfPeNBBJMZh
HSDHi4vbUejgSo4NaRc/tKfmZYrrlGqKc1Mzu6/K5YiX+Oon3R9jmIrTmX+c1nfAQvENDCAa/4ca
clkS/GwVJqem/tq6QODUtFFQdrFYW0oPtvZMocjvOzM+YqvaqsibmdR9FuLz4Mvvg+OGmErDjEIF
olY9dqACTnJPlOHjes9zcBBmAA1UVROD9j9yQ4I9cY8ejmXFvPpEAGstSvMtt1tKi8zP0iAYonaA
HraRO8Ri7NrOqlGTHYcHS04WzEaf3AdZLx4PnaRsilH2HN2cfg6qyOvl0MHM8u6TRLa/YmbPdhny
Qy/Kw9fpHQtihflSShbtpSBLnGl+4EORaZmZUACDmFhiOKixeZlGhZN5QuVKWjfF3RGzYXfSWnNy
u8hxC2XMY3+XMI+se21G0f58F2dSQ1DUrprF3tlBxD3N3gmoi/CsOeHXBK3kqQk8c0xUbR64XZM0
i15uDwhtcfw2kWBTj0e665U3AKzA8SLU2Ax3IpiSFIyJYIZ771JV+3CVt9Od1HcJHJWTw/uMpjAa
hQb6zrd0JkjDYIYpgkgj8qJ83LXgg0S6zby2WwAgyXD0ljp+ulIBc/ISBRFFhWzS0wpPEcXg+w6f
RrAQMprzXq+qAaekF0nkC8p2DTLxBiz+xC/aXj1F0x6zEXryQgOWXcJUV/a8zPp9eZoHKlib/14s
4pCFIbhJmtDOTzx8nCDJGBmQJvupfKBdJufia/Urf+iV0rOIzlI5WMGz6/D9QkdUGz+e1ikPolhV
iCZRqOgWiUuKKYcx8plilX9fxpGK4XNd6Wh0n3sN4cvpsau9VwP7JeDAyOOlHYEt7PL7hGabOh6q
symE1zujoOTcDWjClN91DRkOH1bzx69+zAYa7jUp+HKN8ZXWGorMPjg7OtrB+9Tj0ICvJXjfbCFM
I2H+LE7RxtoIGhHCHqe1CD+RxF2JbJybJeMl+/qdmaEK2rGDqkzC4OTyiAeRsB3eg4Rr8Zy4fGrx
2RoNCwMASANeoQ/AcrZ6qns2Ah8roPQdV+s9PST8Ot68C01tsY0sWBAf6CRnkBBXyc3JblDjkXhK
lOKYwGV8b+rmm5yU1VAkRFOZbkPC8ncgb8H/nSayx4hRmt3m6fYrT7k6XcZ4BqmqGUzqNJ7DRHPI
n2BlZqjGaUJidPauRR8JJTZzM+jes7H+Fjms/yukPbfZK7VDAPmu7swVOsByKSARVjYlOTlVYiWL
3aX8un+lakNzdhYlzeyWP0IabpxUUTr1VWEXu0TFei3u0v0snNL6Rd12TZ/yIRhTo5g5PQkqcQF5
E4eUygf3N0ztlcqoR54wgEJvGC+kYUWLUjCrPu56hNlgMxXcKFO/6nFc5GFE7wbDA8umDZdVTAyZ
30bUGQJNRebU5Jz2DTRUMK5TLVU4zaUmCfiw667yk3G7h36F8ttpoRY3Qr60aflp6oySlVGvlxPb
uFpeyV4CRpAlK8Qav/pNXJ0mD+YqroVOsotXgaCc+jDKrk/+LGvuinshYP7jHH79XgIbgulKGdPq
U82L4sXurr+R9QMtFklPqN15LLUXvsPiF1ewGXmyn7hTjZ7w1Eo1O979mit7vHFWcYYy/lFn7vdV
IniXMXlYByvjnILQoONJe+1dg0jYJ2D/CdZDAgTi96vVHQ/bELoyb1j/ZAvtAity1DqSMkI4wOH7
/M/bkvntx/ubLMvGo0ACg2Gut46/6e3nlB7NBJ92uf5C64jjBa73wGSH+xJrDIP3H3z705gdf0KB
sWrS5xKtDGbUQPebN1oXvN0MWNUaID4hAG95WSQJ3QUcY5owdEnm1i0+UWAXaZz+rK4FEtJom1us
PliTdXNNO530faemYzgOxvbbd/LLhIH95UKHpW5iqZk7x6Qz1vfjwFS0a2ssAC8KaPyDo7TLM/i5
KG+INZWBJlIMxRoLrBeIPNUaM2jwK8wJlApIDfe+OIyhTPDOMQSbGV2loYvFLhLMRCjrIzxnxcfn
7TYNDHCIbl/nexiq+y1d1Y32LH1yz4VzB0akYyNuyILY7F6/IsHtbRCbV8bqnrHKZBm9PLQDTCC1
grAMFm5HYuvbYsqspUhHstBRwEyVLRpjLjzeVg5pOM8jrKiF8HK7+qdpCCkm2bGXMxrpmZRAHjEp
UR5JX71DKC+4DbEkCbpnf3zPeGZAWKK1kZOGF/nuiuM8Td8OGugbHwxexgvsfsJ6q6yew2CvcWHm
hEs8DuDxQIqkeoywdKvnLXkKHex/ZkQ3JC4G1ARcwwWwMERz5RVt+f3FarcWtLM7rmA3y3/71Qg1
9KXRCSgpbLRhnA/Y3cjeVW+9pT1mRCaCOgQSINmWc/XVNUmKbPg9Ju3dCgGVeXY+xzBBsVWt2m/E
EU3/pgkvcKzdWniYPVOQbdtmWnWza5YG7dNtYZBOfA7Gkv5E7GoCtYJTBHw63cLGSDKY7mK1tHrp
TO8TMSbhnNpvo5s3U0eL+y3SfDET9sOrLcaRsagKmmpj35bDynidYX9pcrDuVWs/oPO+51xfn7Fb
1cIXgsUdDq9KEfLQTsySpbkNycmXQ2eBdjn2CIImAftj5tWrWyUETNSDRX/8YCwhL8/9OPqMuBE0
fAEr/4Mm6qO4fht/PlVq5mQ795D8kvmVIQIscsVTX/BRt1EW4ZmWql8AAkmLbJThESLfc1kfKmUT
M2IrC/WBvsyIkAGeNeo88w70YbuXfYBnCNhcpTVq/YT9bIIC9I9gJJr+X1NFiZ4g5s13b1tYUq9j
jm6G9HCIwoikQfkWaXx+MpdO3x4pH+4iwjuloessUO/ZZAJcEcnjR2212Vds4fRcS+7x73OtJcSP
zaSn1+kEPLlQV7I0kF9iMwwfqdmSWbj6yn9v5LRN6lFtry1Xt7CNzAhccirVvPQLcB6tT2tbFwNf
4sIVAgAEEvViVXk4UGyFRfscZo67Ds463JIjnWw7jadTVYlQcWM9VH28C4ZrYhuDH12yiqodZlUw
ILliRCiuWkhiEUOfCnw44uIl0Vws+2CrXJVNbnkGIstJHVrfAtc0Yv5fwb41w3RMkUoDkaL/IwPb
0fSnvewVm7W5e2Wn3UL9k6K+dpOZpy8QilT/nt9evCXFcwhYPUw0JcOMOFbDIjbkA2nm6b2P+6iO
IWqBqss5uQ8AfgVpVHzcXZDi5a0XfqGnZtflUAlb/9T2oYNujS8GZIzBgddOorCUFcDfRHcDgPj8
C2kyk/J5E+xf2rzH9U/KMDIJW7dd3jPp/cZqJqaikyoVXafADcVYY4lGsPWAo3VDjZyhdNIGX7eh
+jaxc9vbgwzI8T/lGZ71uy87yVUU55lBJ2BITff9orDJEgnBLrWfUwiEXG+/sBc476ZsqnZ+AxsZ
olnQf4vaFVNpt4+TSvQh72fLkZnrPENZKecsk65yb/4z0pnVwaqQ5Ee44PpoScnBr2yWagI88iN7
h3j3zl2JCtghbk7lzYdg5xZCL3Wce5RLeBJK0wEvUYLNZXg6/47Xusx5X9k1PGQOTDmIdNnwmxU4
tszEKtTRQSu0pGqHrB2Ibwx95sXlKoHbfYyyS7LbsK+oZB8FuQhyzb+ifzdQfx6fpb+8xIR+we+D
JQFwMeaj6pkMwqJz3fsSAvq7kemoxNpSB19oZWoWUXhTeyqIwUr0ApnvWm8cZWpbY5/itnP4S18s
3acMyGLpsS1c5bQ0tQZQMu+coRMus67qhHpoAQiAzZzbd80IQz85dyh0nnV4sAvgYH4uJyjzU+AK
nLNZmbZaj9NGh/kGG+J3UDOviaXXJpgixwil9kgvBll9DnQ/uidLXWf4MpMMJc+r3LA3BdJfE3fH
AifsKHxuntfRzv1V++bGEfqMAl4KVd9HORmD4EX0pmmJxc6a9wEUnkUbEhC+PzXen52rpCQ7W89+
jdPvyVXdmuRk6MAUaWFxKypGa8fSrBQncthagN3o5mVf9lWNK4JRupMusMTQuNNJVzJ3ese4gcqD
kxawTEyANo56TMDr6OI/R9GfAkTi2BD7vZ+4fgMJu1QtGwoWY9zgJdGQDURHQBc1JnteK3arq1ki
rMii5v48KlyGMi+gDW5SJKQ823xCllXFvHpJbT/KOv/Vz5I08W4mllOwHm4F1uwjVTUYNook3zCg
bRmKSxFPwltFqYwYDuO1sNJclq8VCJkl5KvWoP9seymS6NDoJbUmf58HwgU5SpAFYRMycTbdOQEO
z3OD0aCbtPivW3ZF8gAymYKIcUawPM5GaTVWOXO6iguNkEtjHsvouDcnUFRt9/hDhukQYrbQ4hBD
vv1GwKormn8JmzEjnxdXZKPD9nPrXZOfWgC44Y7OICZLnwmtCnhArqg+A7Pbq5yWETmjqYlPLO7I
g9eIIBHMt1/Rv8ICcKeFHjeMeJECgCh5dsqtq18CH+EN6wVcYrVkYmsWe48zvliSzqKucY7HME7R
i461ASKGZD5J6fr/Z69T2N77ZiZJMKB5+liF0kNqXgIDzHvwiDNN2xYyMpw7EI7++qKTCy0kv6c6
mP2OphrMf9YC58Y4EqtVvd4k319cRtPUhNT9JuI/EIPKrnRwDQ/aVYheUN4cuv3n2rWY0AFaZd3A
w77aLRWIs1GVazfajltJwbqZg0MbgmW06c+R8AUsLFBvjhAEAb/J3Qrvc9Ghg9xLtV01HPHWwpky
B1F2VSOHOif+pHE+9R6e3Y0KO+3zj/DodKe2o1sVvgZ2VvvI6/C44RiXY56ul27TMFAoDkVyY/8l
JEN3Lh3DOZ2hAjyyVMKWmpsH/L5nn6YHGvZYgj2A2nk62fgpH0WLFS8O3JAKF38jvvyZIsS6mjkY
sivhPS4k4gkXqgkVbgLo8zzi1P/dJ80gxXiLcgL+RPbODil6OFDHrs0fQAN2XGO5McF6yQdwtnFV
x3Rv1kDkKfBzr8jaF/g8m3x81931gJMicDMnwvYEI+7MaF8om4QJNPGWSZ5jbmvUKtt8mtrX5Xr0
9RyGrpqmBQXKRTrd1+87Z+wcGFvGd23hTzn1/bGwaAjl+0NQXTuykh3GbNJaTv5ogOuEDfI4jJJZ
8p3VgMl5OZH3kv6fGHazvYVKfFVNVpS/hg0vw0sa6W9aTXrvfunvduorlrrPGPnUNzfj77n3M89S
5uPcYBsvPZd2erGIrN1mNFfEE/ib+MiywzSMuGtc1SDBL9YV1iuwRuIkLzjOComXenyuOsy6nE0N
jVgp3i7RM1oYmjAOJEWvhLqcDlP1ye8LcxeYjWvJykQSanprJGzyuNsUtb6yH5KmlB1I3Hd0HN1B
ObhjaZExZ5X8QXZ/t9RE3YaVbg7/Gt72tqiX/wz/v6Q+1CLlOBjyMWWJZDveqEeKj2ZGXV4/4LEN
fdwgk1c5Qs7wVa/1ySZP0zryJDM3xRHk6U0ENVQoC4sMj5wK7fIm+ixUH+nq6TmYKy3IE0w2v5r9
D5FSjnFruVvObyh3e9tiyFeDlUoyisCOxzOmi4rYYGKPu0CHHJmauDvKuaRP8AT0zZqsXhJKBcKV
rHmsDQFaGne0xA87r/ho8l0XQOjsKCpcX6OLzX/iqVXxkXTzCQ+5rGdO12HLJtPWofBEJ+60VVrX
26YH1vATqDQyG1uMggEYeOunZp0E+WBoS7l+8E0XGk5tXiGR7kO1hqT6BxWs33uhI2Td3zP1IcTh
I9lkXAp9svLL1zufuecU3wCKzH+s5qtmmmPb/dXIWBrxBI0VC75Gu2PuYP2bimco7nPjVvwbk7qP
Arob4awGOnpVCe5dgNRQplXbBUt8Pf80Q4o1WH7cO3dBlrCa/zlB8jBP6Xfyq7XFiApmBBjX4fvr
yAWEAsw3e89B0yow2qJC6TlhMLgX2E4PpF/YhQmVR2u50DyGZyqIK+a/jpx9Y6eQPTw3gMThmJXE
w4K/R4d4D59iWL4pPAPlb3EqZm6TPYtTD0SzidFpfewisFYKUMJ0dUWT6J7SvaErdtYvGbsX21CI
eYpgMJxX7Pj1enoK8u70jr9ucpVHx58IbqFrQzTB5pr1v4sLzBV62v/kToXuowNxapQXPWsPoGOd
c9abar5IPJ9x/k66uCrxC7c1Kpd8Ydmc0SXhuNaMI7IhIpqLh6RUMfZ3ydPkWHA0qt98Muv3QnYM
NV695O3uikx8MhEPx7IVyROZPp9eRlkQ71wwvbNt6W/olbd/fNGOZCN/Vra2WYyi4DVm5KsHO2x2
ERtLgXR20uq+t5QO8YyqjYg2fNapBdoOT8HeSnCIQKvVy38MOEXlFNEKSuciay1EXdNrnkAGuJJb
JRVe1DvZM7tdsj4kyqVCbbaGhxIzks/CxAD+7RhRITxBgYI0ymW2y+G7sRiZst00ODCj2i+oheu0
hc2ldTQC1KI07Pguq47k0DKAD2IWp/HJE1R7dBl6M2jp8pUAkGS8I1ljrd9IDxLxcvc/8TpTD+gX
L/J3uG6qCN5TzYvVcRhfP8BtKCXxbTKeJIWhRoaOmRtEt0xIjKryF6dC60R7QmPEKWxnmslMjEdM
e/kITnDagI8lVzeeHdpLnf3kyfgFu3lpgD44hl+XGvN8us1MunTvVPQER6MYFUFjP8ER0J5sfBTg
dEh69uzch+Gzx8bX+vw/tfJZXXoOPaoe1yjTlILY4PbCHtHp4WaKqm7FgZo4r5UYtZvSBPq3wyyz
8RuM7mUWlFdErdcnmI1ogg4UWxBi6JB79anKwSU+y2HO2ebMJSyMrXkpJw1IlZAEu66d+yKzvGPz
+1/0uxmEdKrZOPtWfTxMdqmqZbqzlh5gHHm63l2uURQsGPcuWuQrHgPOzdM2J9hXLkt5t0Hc0MFE
3bL0ASVK0aONca+IwPAqpRLPp6BfSZMruReY4B0uEhsfQbeibrQgJO8ayVLSvEm6DRnGoC1tu0NX
gbIiS+ibXePAWJ9b/tGE/G+aSkHkg7Gr2k86hSHHZig0oKtOuiM/dTrEUKY67gWI/LUxCsRZmgKH
BaU3pxXzgnEOl/ASmgi3RRiCnAQamnZ6zLasb8RMToOUnOKQEmdKB3fEd6k8V7+lcXMeUch120Hi
tX/hpbnMF7rYXUOh0zRLAsL66c9CreKIOJcajlslC/GHbnOLt2PMIn6nerapGv9fM6QL8sLo3Hqe
Fme9LJJNHWorQEZNKHAh1LHMVfcM99l2Tk76pW+h82Sywq5d1vOCzYlk/J/mFGgtnLcgNB40MS4B
gcxYuztJ03gGS5SG/l6VXFZZ/lHpMN37Rk0VZERp6idRGiv8yduRdWoaIVAIfjrG+a0PlEFGgqHI
nZHKOhHLeor66bbFghFfRSRhf7+8g8AEp4TyHILjBm7/Fxyk3uIkBgGdlEO6IBdLZfAZUc+WYPqL
VuAejV3HTav+iqOlBPSiF3xjmb8scW530+drGnSnbQb2bHM+EOytxC6cvaLa0jQuCmm/2Npp+gYs
r27NNLY5s3163NRPSQRcu3Ejs8spTmr0Owp/n7cEcHXL+PB6FuTZG3/svGED/IYMm3m/CUk3Ehjl
fFhgl6sup7QNcFljlzseiIFuVMCq+DzAKdyw9Rq7yrTISzmyNTxxje2a17RBP3luvzShQmZVt6M9
pZDPI5hpdODWQAyQPVuXta6Z7cFkBov5SqiIAWsJ6PYTaQXCRidw3rzTISLPaUFtEtxF56N0nNaY
Caa1rtdv3I7dAnZqs7ZxsWZYVxCCrvXxs/V7XV8rwVV6GtlSJUFxDgdRfYm9YGt5OmpByQ3dNXLp
feHBlM5KD6UpOjtUlyLGsF3FlR7Oe/r9ACr9BOhJc6QNI35b+WgAG4vIvpd9NzsN9aizfClBAUg+
83BjANG/UKvRqI1GmeVMlG2Q1rHRckSdhYqPmxPBXqqnew+41Nf8aO0ulRoty93k4k7w6QggaIOA
C1PqZSOLSzIGoQAj7IuOulBt6Ak5f5Ml/bs3dHGbutgK6QqFy+2crUd3Fi2nbAMW67PzO5ZI8epZ
elpOsceFyE4FZFiIZauw1vBjKYRg9mPjboZ8QeJ3Z9GeTEG6YvB8COMSLnSpJ8a9q2XEFmP2gnxN
BoG+ctBAvzeIwreCc11sQV2vTxJ+UCp3OvZkNJy+z2QhA7CnQvmHDpkFX6xLFJVo5Bj6u7qwBLBJ
lR9VrcBAv2AkQyV7UgzwqSRI5nzG9Bm25Jvb3EYBBhi2RkCSmmMbmJXN+I6FeCv/rsBvLOwenXw9
Oc9s6ZDzwQm2MOGCUTkwEVnb3vhIiZGyOv/bv/wCb82duj5R4TBXpaOj2M1byCZXSqcDJpqo/jbC
L0ORx/mDaXJsJQRJp7TuAGI53ZEnclJwSAvOZoF1D92btLsVx2C5zQfgb/gufHOsnCapWuLWHuu6
6BiuE8HgHaOqSBOyC2/vccxb/ZwjqwDwGuC1HLPOWXBLj2n/4qmjg8yEn0+WorfEzK8E1qq98spq
sa+xbmfNcXxNfwJwUt7LGTKBoW0bEFW1bdXqHaS1bHpf7EneUxSb/axl79vgKGx43pY/xPZfb9ZK
WYzYJk+saUktFXLSs+qC0BSHRQNlLR5fMmDNLUnXf/XEi+wJybDm1bXdkn1Ulxru7DQlO7BKE/HW
IYgzLUE33+xQLPVRoE2w1AOwGvraUhNr7gY8Z6l4e/ZAeq6jzNVNCSEe3OFVBiNz0q4fymtJm+lM
sGUWdxcKJCb33HeM3SPzqirqEraTeNlyGO1VIlbBRzgoStG4u5L0FuznXl6agjqQppCCuj3tuM7T
GkZKhImOhOd4R4Ti+481TuaaO8npLphlEv/IDwFK0UrB34v8ogwj8Esu+Cne6vRhT4CqqmUmFHN+
v7I5L0SmInZ0rJW7R9AEhZnCsIPkf9pJNSLSrfh0p1bNvpGOwwM+SRIqr5OAxGbgS+KlgRnbn/w2
ZA8yD+FIQCObZiy0NOzukiRCKrRBqs2tpEDg4NOGXZK8XmNud5MJ0UPzTRsZbi/MOnJBu/4KAqZq
aZUkWk7RxE90yD88kv/yFWoNzsKR8dBE9HkqqTMaP/PhfVkhKNthJcGGd8tuBL/vYkTA2+3Tc/uI
tPOEpa/vpe89pjyUHMEGsq6VzEqJ5DqQrGAo9zQxEwxnj3mb8JNORjfkpkhV4IAtSIOhL9uJVCuL
DsPJcz8Ye6QbDmn/9duhiZvDFI28/LxX6v6Q33aQw+M/4oirz4YoqaXodVmu/d0Wd4c/n1Z8bqoE
WmTDrt3pDLqEKStTMg1AneJ/e8TeYjYMnyCIVxkoYJNZ0IDNaJEFOeWhjqcF51NNG1PeHk5/H0YM
kJdRVajK/xlXN21dEzA5wBRlm6XraVonYiAsv3Aa3qloWwbWpLoAFqxXdqX5DaJnoWn3rNAgLIc3
kSeAqxCu4LJyrWQ890mCBH/aZMdKRAiJf7mwvO1oLQUwyQtnItkqG7ZtSMEiYGgj2twFsU6IFRCK
zJOJYrOBg6nw1qXa6rA2tMQxG5aylDFuKRG8siar6Loj43jiA2HWLbrE/80TZyZpPXpXuDbObhEH
KpVY7jqCN5KUUhRWkHkfjZ4peOyISxjsDmmOemF1TWPbxvpCzUDrliMNihDBec2/eoxQhk1ZH92C
Asl5HOTBBSEnAPtSKrvYa0XOJEL6V6KKFGQPnrbm3BuK9xu3FjRicTMUVWx/L8ZCE9Dja43rrgba
kf9NXgg1ii3HlJsEZgRdN50pQOBiGJbfckIrK728A8hTKiaj7oGJ6DlMQbXRrVxN6BSCybrxsmlx
WFL83K9JxQpojyfVyq1xZrJydm/0EZHGlkReIBPUGpaq2/ntscyDvdTeTNzCHqZ/Txk86p8Lz8fW
7gYScgEBXUEeON8qo7pVx3y2wUxp/PAbh/aLdXRr7n1ER5CXuK1pwsLFax76FnFv+zcyBEH1RKfF
QMvPdw+nsp0QyW8A1UEcFktz6DRjFfNHg1Asdp6XGujsPxjK7EqjMM4QNurKeY1hcrRrQjlJF6XG
VYtka38ACaaMexrWPzuxbEwHRXtO48yy+a5xZvwex4pzICYNF+zRF4oFa9WORnsznnf6n3c29dbq
np20jG7YmS0dBZolgaSYbHfYfrloNjoGJBzSu5X5mdIODve8Xujg+j8i9QKzJCMqS763SLxCJooE
KCTCpmYxyLd6VPkXaTFChzBFjV5k5NgnGb01r5f9+HjyShZvBKwEvddZoNxr/zY+s06Su9cjsaeL
uvXyDMufz+++5x7waoOxxB9lHrX2tCA25ndK73ZeOK9YCtPO29kNXrUNPcEbpCDBDW5pm7TGEnOk
1eMUm5R8Y5nlpCvL6Ss23Ox/xKN13CX0LA61dZkh6neMWWaRh5x4RuMWBL3JONlMS6VjuX9idaxo
iCUor04QAcYsrkt3+hWOsD2p/RhGzVM2+05LnzKJkbePGjwPiAcyLmQR8BznOiNJjp/lyT13P8wB
q9PEUbbEWIxnCV9g9xjj6ydBbB9YnLT0IYjmVCDQhlS3lD9PBkesuukc+kRHniUG5sZFW5Uk5srg
r116AiHvoytYIaArSkcyeotyb4itsQZKPAfuMtE6s+n0yCYUFPkjH/LSDcicJSLkyj+09Z+JQjg2
2+J1uTi46MSHBLTIt+sXJxn4ArYOASIpff4dRm6pWuDkN5Z5OToYw2biEP9XuE4NybFgoQZ2+ozb
JgyvXvvHVJopvNyey8ndpRRjnvLHxs9cbqmsrSoG+BmwB5vFFK2964QrvVtQCKqsgj9fnmfvGsRJ
hFD+TkU0O2WVvSuU3Rp7sddf1bJ/IanpPdwHaClYtZIEe0onPe/mwfKtZ4Do+K1DCm/X8XIsBRsY
hACra5tnuG3mjOe9+/f3pwqLgUWtSUhjXTDtlUtAxp3ht+s0P6JfXwM5whpD+ZeVVXxt2OqStVrV
VelP7qiUkhtzS/+vddiJ+rNw2Y4ZwN/d+fxi36mEafKk3LIRbHkDpQLCChs0Yvl/wI/aYXsapvo7
E50RQgE0CONzlvHyHQ823Z99XWlFKtiaQ7KB6tLN6rD5MgOUOsligpbAxZesN0wISrKRgEGyby41
onZqo5ftShasT0WH/X0O90Jy0IJa+jP/iEetcBgwTg3yO+sD8hODmWMKIvnUM0SgDTI03e04n74q
PWSNn6nOu2UvXR7djXnjx/6e6tL2mEnAuNXqA/77xTCDsuyjEt9jLfQqEX8sc380bI9aFpbsbW2K
SJaRGasvi1ATd2LwBlZMS19f070tRQrk0GHG8RkojLHA+LH1VKKQKJs6z9ziPmVhvxqPwEIQIOmS
m1meY844Wc72KNCwaBcsYvQMZRw1UpGSdp1GCQl+eK5xYg5ijsy3fI5PNo7aY/o2eDIyL2i1Pgcf
UgFX1zxjN9RFwh4YHbFJme5yAOTnKE6GsRv1Ijkb3FbFfnQ4lvkuLkxMo+zLnRyoMvromIjYF+Io
hT2XYOC3uUlZa8XAsoYghpwXd9rjQKPevjC7kO3kARp6MUR0dJFf0EftlzEANcR/BVn+bSG+DWQk
scsqYIIQFz8tB2txKJ81xcRGKbGEh1Yd2scKAUscWY4xy94rn5W6Stp7FdAJE9sMHBILnMlwBgpw
vPercP5KTo9d3c6PIfvIhi0WZVuPoJoe/r0ui+OLjX/ey9iqf++a0F9MjxwywXSOoDDAsB6ZI+xh
f8AU4iiBR7vyUbzBQN16nMr+fbeFjTgv1xVdfG8x8xwt75sllF4ztx60viXlIJSsldFq3cqR191U
hK4gUORCEPBVD5k+FY4+DcA5cQgkpd1GUjf9DzeG9i6Cos+0pwvgNHBgqwua3Mw8D0IPpLaX3YFx
p6uxwq1gofIyNMXYk69wlJRL942PH11YGRvhHhz5IW6n0xtagVyb8ULspq52kIuMRPwMxN7AP4Ur
YE4Zk9rLTyT9Y09fw8Ie/lG/W1SfA3bnFvqmPp982JZewVJWInUPOtv4cPPQj7ihPSRyRiGn0KnS
YeFodRTRSQMD0ma94O9EmUyGLdnSPhOYFVPHmWmDfz0HFbaSlMfPKn4UYfk5XPA5X94bEjBxTdpy
rOg0ULGQo2m/T+Idczry0BT74yy8FSf4cD5D/WRqYXHd0Sps632B0NbmBE6EDdVsB7sZKKWv+Nir
hTC+NkqlpoSjwfD8Rw6wlN2jFX3MA2Y7UDVppc7wRDTvD5nLb4cu/K2gOQwZHhLyHEdJXKkk9L0M
6+cSLQytcV+N9IxYX+NYXwe1RkDFhKHx/Vi/QXYlPpkckA17yT9h9fbybvsSXE5V/B6SQZzvIyJi
O3PTptQPQz84VfKD3h0+uzoutgnmeeyRjbPjsyn+St2lkwv/Ijz5Nvx+VDQlZ0jwU3w4woPUArXd
IdEkKFIY7yDrttd2XidyCWhX36o14PJEBi2e4IY96cMuUWBHnB+CLd+Ij/R9dtxBveS0VFwuSLxC
Et+SohqgPHTOTFUTgMn705aq6s9UrEh6IuvVsBwxBaL/uGuyRBErWpaA2kvncDbesDjiA3pIN1S2
9und3tH337jMrdgF8bmvJAG7ifG62D9+E7q/zMk8EEn0jrtWxuryYOPwYFd+d3jzzvhm8JtUXnE+
rFg02lFqOJG7xAIwyzdCih5/CXo8mjQ+UCLcrS0Pg01IxAwC/No+KuVBmVdO1w11mJUHrhRUzrep
tkdGDuZHWieMRhNcE5XepgSGfqbswydjVHEN1LPiZaoHVyuGw88OMGlzCQQ7gXIYA4W7rGS7NIPK
xc+5VaSpjhYgWylCL2kKdKkYzsbvshvKVnK3Kgs7yb0Dn6SSk3+yseLKNpE/ywMAKcSatq7pwPiQ
GSwk+OG6bM68TYoJQqQIHdkxcCLzVG5arLQ36GIc3l9A24QcRdRU0vxhgl0DNHmWM/WxItA4gKkF
SdlSlZAlDYcQfR+o845UNxo8gKUULjoqqhg4XdhHr2+j9p7CDcNYJB/rHJ7Eqt2LVi8JE4uFpNpv
oc7DXGqtaw92KSxYgf18eiCFZKHEHqeeZBWmRmrqzjELxmIknQSWzr3Ep0acrVScJIV8gKUH0eid
FfHYHcvFzXvqFT95aAjYXp9ALYy/aCJnlh3dsM5hr7zR+ngWDh/o6KSuXp4RFcpFfnzMGuRq4b4x
lAI+kjg3546zJ+kk+qqFnmdu9dBF1/BHtGgAG+8k9Bcs7lz+88zJqbZMo0TGEMpK0F1Abn3GAOhO
vNVJ/KXGbKzuNK14QkGN7mD9Opyru+W7xTUfDBCdB6nHTo3wS9XckRFVK9DmAC+QzpFr0Vl7Pf8V
JPeAzlgDXeFy4eBIehMbw5y63UZEwuWq1T7pLgm30JJvWI1ywTqEZXuKFB134bT+ICPmDkUkMD7s
1l/tWgs0+DBDVrn/GI+m5g70AoJVL30Bk0ogI1dP9ROpxWi5CvBxXISHIcvN/Kolc5rgpFoFNZ/+
bbJxTkKrIhC89APcqqL+syjGFYz9izerlVWKkm/2+wlZYX6c3HzFVEaHR2+GM2nrjUEVd5jYd8xn
cC/Wnk+QQQmz3cirA6GLugKYWFPm8gnn2+tVx3J1AKbEO0ZG/68BDXcY5S5mRiNGyMqwVCzkKTVj
5jFTO+7qD6I8SxHIFyBV/9moXtdll1orP6GCBUuBeYbu7zqV9+y2jGIvmc00T9n0knDjes2pq+WQ
hLe3EB0yovNd/agHmGqKodbdpH0UBDBJTfj32rvxC+bkyy5Fe/LQbxvFTqbw9fiVkbwpLZK22Vwk
4onarEoIK3H75A5dtSzAuZ+ul+nCJjSaVyBILHxJCUPBEwgeORnzEPMcpaOQQyKGYK338KzAgNcF
BGJxeytoKnTEyN9lkC4zWF4mLa4HkBtj4kv5I8Jve9Te5eVl1m3TZKZr6QaxK5VBCkSaKZDux0aY
5K9p6Mev8tYtmITtSa6DfL3IM2bfKVzNaBH+lpfAEYUr7ET54scXljZGX4UgdGgfqZGJSmGj1YvI
HAsc8XLXThRG7XlFgxoXvnBHAIKKC9W5GqgRetyYkemDt4cttfou679VjDJBl8Bsazj2mmtIqStI
0wxi8buNPFCwVv4cTmeURFeOyF+UDZZrJBYXm7fIQcWapRDg+3csicLr6DF0QEbvARYAskHwCeUL
FwaPeATvgpWW0j24+I5cO+FrljX0xiA3RY42emIlgEJy4r37hoS2SpHxTKQRH/9qFTaHD0kdPR0i
NzidpIkANhPoFGYXwHMP17xCb3k52XgDCBWNZuqXTPxOiyAXdRli4/2bxDe5lT6qv0fRakfKEX/r
eNRWTpql0+Wg5tP5kbbZWMJrSgjStmSLI2r0wFWNn7ru3yNqhcO/Sd0+Y+2VFGiqij7D3ZvTc6CD
EqSkYXfpjHDK4e61jilJvr6yBeMJN+SsoGDYkmt72/5oih+GVSBu26H+fkhL4djQLcDdFLWm8DaN
jYHguzPdbzp/XBgj4+cqlDNNH60rqtQxuOnH6q2aYDfXRtUZZS9s6mIF4Cpig7bd+HxisOjhxBdT
H9bhucI4S4e0gsnEBsaJzP4XZaRoGkGgYfVOCVN+R6l8bezWXGtbfXu/daBEWFK+F+ghC1p7CdvA
uEtITDa3RP6AAm2kW9hz8GcFmT0C882kZu39KJNrsPQdKHl2q6PBVIjsqPvvTZwbnM7M3a/M7Eea
7levp9g9hJdj1pqihzFMxnaZfiMhsbdjVRbo0DZkorx5/QTEKh3EsnM5vaFDaP7Xulw/vD3aXCFS
Olvom4WHbzovd7Mi3lZBvkUJ4UcQ0ZLz06J6gKR8BwqUUhFskVWcB+V0WTYM1/8LLg4fPTRZU/vf
OGTsMaUBBxitfzmIrYowb7uEV29ccDeTgMTN21oKqmnrLKpGGeD6F/EhUaAYQ6ZeBFvL1Fz46chT
+SZZUBwHziUiwM9Y/+4+Fb2SAlcrcvLu3wh+8gy8w5PFWNXcrtsBO37KCLROhDH40qoH4KQTfey/
V6/hIk6NizUlLmBk7kOpjPGK26lse3KMLyLejI6Nd9Nw/D25BG8LHA7lMboK8g4qdbg3gJdckuQX
eEp0PHID1h4GUSaABjxCwXm4LWiryeelpTDta4yHe9MYIaRDsjfjBH2/jFOlUgpB/ZwCJrfu627v
r3SSyJOqt7VYl6Z28mGW50+Tze4srSvHx9tmbL67cNvBHZwWA1utVctgi3DQUx1lb41yBtjI3SaK
JGBuXWCPkM4K9TiCPO0/pHRX15/BJup7quLEcVh8F93ayU7135ZexGsFxXCHNe7PCD8hyGX110vT
Js3SxR/RFnsqnvWXEjP6NKu898F+ux2cmwzWdLtarllqhLI2RJgfKnUeLoX6KAMmrs1am4nZS9to
y1FEjo8N4etsMpPJOok19+cn12WsWZu3jLO2EVukNrr83htB3AIkhUQcNB7lqsoTy9/5WpErLqgX
xZvDUpr/CU2hIMiS/SgmVpBWf8SaeMbCsQljFdlRnEV+bevZ7Jlr7OMVCjFYrPKJpWxK6W6Ztl2V
pe5VTdlpCNhFqGIcLW0hZMeUH5wrmXilYm5cYR8YsmGGMDzqyJbpuF23zF4rrLp6mAM6VOEhVhPG
OgclUFPnKVkek9JzOek5LJJObTWpZ+LO6YfuvXPTCe7Bj6TFqZf2ZG+JuJTFelSazt3psja2xLJY
/dTjoGo1rQK5FT73gmo6Ueke7XqQEPpm+YIfNRP3cjMhoaekeYnV/RzgshmsEAMLkg4rmHHRzdp/
RgivrOtoxDyTN+VkMZ6W4ru4nFK3kmJpSvfW6Ht7T6QuSGNxbjaZX7bD15mDvaF6avQBMwqYGJ7P
4dLyHQ0Xpy/Ix5Za6A+hvzgQO0fLlBesoptUlRLuJyfjuX36y68mgvSUxx9D3fu4aqLrJ8QdvmO8
cVyzlpzUjbpZMxsTdfHkhiwQLZL8GT9d5PUwmywhmZBgI6DHMPDKvPi63Dmptb6YhVvdEBlMqUM2
fn+4E7LblCpvh1MqTMUKsR2jdfQjKBGbe8p5oSOi/A69vu9KgfhPvWm3PmcRidvNi0gn6QD/uwS4
1Jsv3n9/7oHpsQknz0sQ185xJfyZL064T4WtMCr4JspzlVeScrxcNfHEVpYBWuO0+UftTfVkb6E1
Edw7VG3MlwVMUkCKQRXB4AxtZObinKoVUYQ3mVsUx9qb/INVsPkZDR1Y51o4PM35SVBYyEUAF46s
vOmVTaE0VjM1iqwI1Wty3IhIU9a7T3ChCbDKCht648Z9iBnUrgyHFUMnjdbJ+e3jKGpS26UglN1M
POYhdilxrm+oi+4bCbZT34dWgKVd5DPrFUErqE0UgyR524YnZxLHEOou9PKNncqAKPDvotN88ht9
I0UONUEislpeI4WxnZKjVKmno6fk0QhqgriQrZ27Ypb/eWkJ4846buCOFJeuVV/4y/0ahcDb6Tsg
YZeIIu+ceWaWjk9TvItaLhsUBQ+dCdKL7j9mUqwoF36Rvj3VRq+Vhrj6noq0vow7GEY0x4SPF7Bq
MPuItXl6z/cFLGhkKLh7U0vLpV3fVK3yN39KUgNuG7CFQ8FgOgbuVxQOcjWVyMJfGy3VLzGEbV6N
/2BerrQsDMWJjC0nKnd+5oVIF89MJfVOQwZnQvyXWseOLXrNmXU9e6GmdVZSI6FT3k20b2U6RA81
fnrj82shdYyRr4Xtg8AovZtbBQo6iO2zJJEblHYWB3lZYtjzwXMPIh8MgkgSCHG6Bav1RbR2R529
IgmTAP2W6aR3S9ZKUDIGAvz59fT7WrSMyzM0JwQxf5k9l4ENs9on9wbUgHVKXELpwAEC6cACedm4
S2y7y2N6wRIPHvXIN/I3ArPzYvB5pAgbB08bJybSwvXxIUTZEFyFX1uS346GSpW3gMmh2TwxZUIs
jOUPBN74pxtnmK6R0ZTo+q2Q4/4/5q8pHGCCCxJTYX+YlWo2fWU3EcNxgpOUGYP7XMkKb1R48L3P
W/IrCSeKjjVHhA9a9EYHZAdbyi+xSF45fXk+ufsVJxMdhnMd1kLxC9TKaIAl/A+cpCLMoO5QOAWA
izKamx7hVmjPpqbUMaTVp+TQL+gQawonbuoSQq5j07e8wEWVOkvDwx4MxwjcqE0v169o9mryBf0N
e+8hQZRUSP0aMw3jCCytB9k4JWHCuUOIQySp/FUG01aWuLVqqFrcs9vw8rrTCfiv8taR9zgzFuhR
PeCc/kG0sELUN+2M2191jq58zbUI1zP7iyEs9r4eaX2CiAakik4O3e2Jb1xSW3PfagNx8/pE1xW4
qFCDAYaEA623DX/7ZtSsTxwKoyyLxXwHyx06hOr3z5+6XnW/7yK/GTW5MyL3DEZs0iASk22GzLur
iBRxub42B72uipvzRKuhmJIzO+ruEfJg+0FvXfAGSWKJ04dkZpLNGnnIpWxBgovGYzAesdfjBeIS
+AR/p07crtq4y+nneleqdSrfIMqgwkgm4XgwV+ug75Q/VWOnCwGwUrKiCDwu/dTUb4TKv4B8b2Jh
5ZjDD+LolpDJtUHJOBRt/V08XkEBtuxwP7P4mrdjl8dGUKM17s9wS61w6tL27vWpf8i6fBS3mfUZ
34b2Siax0cu+S6Z7CFOHP6MLR+62KZf4TmCtTtK+h1K48nFQ5bHFHDDeU8PMIXmpKDTlb5kzUUO+
hYUKfZp8QGCP5hdgLrR3n/SpxKBj5riFt2lwWWd0wdsQ4693yPtJwdGGjBrZOYmBFcOPxwjkz95A
/axtf6yCtRVc90IbC5aU9NzLIux85h7TsKJvT6ewZT1HMmNP8Cho7+irVDH5h/VPaBAjWBp8LIX6
v/QVmTo/v5eY/3YXjkKHoAnkSSdTXleUSz6UAjj9UXQAiL3d1XlLXeYCtTaHO1dDX00FOqxdcTpT
LeEcbjnKSjeHG/adUa27IPFMuSDK3TDiT0cLgMGY4mglA8TNF3e50T11qxY8oY/7Ow2Cahp/Tus/
YfgYTzVXO7YmGCLaGJcq88piz3NHe/X8DQjnCV+0fhwinMy8au45PlMXY3mTe+TR/g+xTyDWClGf
xsp+zvinroIIoMTAAaXrCFTeNVtmBiSvk9FZpkEnlIIv2O/AOtJbkXgpM748IBJ/W8HxVJtCF48G
Im8oQW6UWrPV+yWnIu5z1VVo+IHVaqTiEe61A8n37a3wr8FHQcU+cNDuqLLy9eSTCzigJcSMIlwc
JZo79lYi90P6vDIT/5eWkAIaTjMyOuMuDR5aRbmq4Rzh0ykQDBmancbK5mUS6x6p2unI7hymHbCW
m0vtFhnOcndi+w8gdwvaHzLQb+uQdJBf1vn+nnI+M1qc6JPY535XTd7QHTMHWzHubtIfADZaCCOT
noJ8maUgDOpt3DhHkWaBlZmFsORWRaMLWgHuxTzH9dGWpMohBSjwZ646bNbsRDxx8XWQ1vecEHut
aYgIyhjr3pUJJknE2Gv5/yNrPtP57pP+4iTW2gJecvTjvfdRvYUiuH8OF8Uqnu/JCpcq0cM0QUeq
WelkqHe1ci2c3TxgWnq6wXtfxeLMR7grNZe11Mdsv+Xf66xtfj1kT/IKzZkPDgYURu3ugfAgDSXr
A76uHrOJdtJu+iBGJIGmuf8Vazrp2iZ3NX9lpKDIz4wNMQ/dWEWGjIenvENsztPLJh6YlBfbqRAx
5JqbgjH/qZaLKiVNRu2b9qzakEDu2OHxhm8IUAlKW4NizjJFprVWIvKymqZ0wHi4QAlOAjTVDuAQ
XAlUq5hO4J8El0t+5yMyN3lQhmnOUEGX4tjs1wNdXJmo6Vdhyl6vAPxJlLnP1E//Rg56pehi/5fQ
Ok+Pe5x+Tv3q3yoafGCn24wbSu8ECFNudzJL2ZZMAqhqH4UzSLuv6G1aF8gNn3jO2F05Ka5nejJx
DdOVd2FBF4mVi/av30Aue6dqNinCl46hroRAzzZbFR+DPK0sud4y1yJjhaofC8fWw8U91cfrkn4S
fYNVMnFqoA/xfecDHEFAd61ChIG0KhZpN8KR8hDwqZ5xJwuPl/Qg3ZWzJzKEdgPQPpr/8Mrxq9We
XLFDNEUCEaO52uzWfr8kxvGluz2IGm929hEudDv3nOWWtJ7cS4EOr5cFZWIMfzN7pznmcZcpiqGc
I+RNJReR5g6ehVkc1nXs9YRM0rElz+x7QynaWcWLLxLPd1tI1pxjc4pSqhk5r68EcyIOuk10w9eb
aclEGKBFk0qxCptOUwQY/T/1bzBWmseqI9znidYEAm5fvJ8uKd6LQi7agfMQy4OVbP6L2D5vJWjF
nWyL3zecs9Ehrp2MJXi/zGGITZFVjpXRmlmEI5voZnKyfcz/Ch5Px7ENuHYSruzm9L+vE+Ip2V3l
bSPCtO4eRYMTk7mgL5KORQGp72myHIW1RX5R2Ahhrmc/1N4oGDNJ/bKfb/2D0d7u+040ZJJPOf9a
VHiKEasrMp30ORC+bjkgkXMGrGHQYYbnpxbeiHWLajTwXD0X3sfx6mSXWXgxCsqcqMuTZLVipJOg
CsUWhjm46SlcwwLnaWQFb3FxVsdkE8m6TTjeakwIUQTdLKdkUSJ7/xXOEUyeW1SPtUgXIKcMc4aj
mHyVt18apRAwCOnxH6AmMFf58V1L20KTUI8x+N82rm7OSjoa4eyhSH2TTav2e038OQUMgLQneiXj
R8GlxUgncx5D61Q2DNm/04yxeGuqgxKl5dOwCVnzL+C5SEP1A/89WDSAnyNRlZMnh3lW0/Q0rbxI
Ifn425LrAsGTG0bc/yIIDIcMAhcw1YYSK/TQuYDlts6GNMI2TU/jP/X5wk1CZGQ7jRAW43zVnZA1
EaURXdcwLJDvPXmA+nUf6YYx2mgRQgheoX6K3W+sPkEwZG+Sk5oK7ZoMw/dQipSfMJi1zNZ1p07+
aZOUFpCloHlB2Onvgu+kUA4WUO+PgV5XUEujGPqYTMkwgCqgVeQ66aAxm1tbufqgYrkt0u4t5SUF
4UL0UmjT0cGnDRe+xk8+V04Gy/dpM3i0C9Kpkgddw0MUGsOqFnERa8EQDOhwv0iUw9Po09pODeuh
XT4xHSQwtx5J2mayXC1HPwc1NZZJaaYyOrGqE1fPHV0BiU6Dd7flRqCGqKXnbLPy9D5dY0KvewjE
7QYhO0LEwfPyZEk+FCrHtZ2phoef5LFVX3+7PbJUR51oYZwRSTaRN/B0VTePW2KuosOWvLdUGjwZ
DLcM3lTDLCf/UvkNewjfJFyZNLsol3hCf8HBJbUvUNLvjqR8o/gMnx60oR8eTxp8TC92W6JjE8GH
c9n2KcQQTyqVr8lCVfo0yIXTe5FxQcT4eXrdrTasKAwt+dusuAasvg6NSVI/ujlgdXyp1IGoK8Kc
iZFSq4UuIrfK27jVz9Tu/g1RGFIlSC7Y9/v760B52TONOLmUJOeNMpb3AK8h3LoWI/HnBYwCvYyc
kmM3mIG85X1UtEn0yfM82QvMPf+m9SYKUYFRTyeOtrL/GOnC5piliJMQIrAHh94ASHdyfgyqOhSl
mcAcqnWzjsiRDjcvJWNiO+fOBKFplJlkPgVd0D+E0etXK9pzZgpM/cJsxrCO2ONoSQ2yFvcVm876
rVcfcKGsQY6RHDC1jgROeMd8hPlxixWIpUeE2y7Fo0v6To43O0xllaNSzhZ273UU/jBMqQ9twxAX
xsC+/png4ehPisgbC5X8ctJHJk/8NC84OPwAjcriuKd1hVrTBzZvVpWT6uOJXZnfu1gWhBV8EwI6
h9qlZULKBRjxpZm/bCxhoZHe3FkhwH1X96THREKNqZemyHMS/N+jycIx7PURHzZZHnhCC26lOpoj
ogo/YREV1jxHxs7wMkbmMySStsVjwyz3qUJIB/eC+xb3xmPq/tr0IUJeah2iRMoIei2UJJpB7XEg
/puFToJ49XhMoMdtnbGnmXipAG31WzN3uckThy6/Iv0AsW6zlCr1MV4oijigXjnMUzxWfTvKV0kl
1Gfj6JVpYxGMQiY/Kb/Vq1UmuHTxqYspsKecNTLEZgXlNN/uG/0ibaXMTWNN7/w3gWb7nQRTBB/w
ciNaxEu1tkVRjEi8mXei6civowwF/6kaChWSAl5WbPJoLz6Mn12/5bRADtSZ3W/J/tAYbuXXJ5lm
NqwGO8aZVRBCxTfTRpTqLG0/QdOZT3q2ewknZZjmilYcoyhXwpOPuEb7CrQuL/qQ+NsvC0CIihMg
L1DrrM4Ww09uMxGmc99Qu//l3CqTxr7E4w5lIkn24LC/Q5dYCw+2+iWaWGtmcNMyx9qhEGGZ0XjI
OphOuE2VBaFOXfZCnB311/3iQGEtjIy0PAUoOtC5Wkg2+EDK8ZzQwGw/I/kfIbzPD+mdtuQz8EqY
8pSd76ezL6Xk/ETvR34FykVCL0eH+lZF3AWMrmFCO6zFgdOZOMUwtUuzk//C9wRWoOHsP1Yj3+5G
8Lw9nksN+dEf9RqbBkHVnHzWLVx9TlnWAC0b5EoEtj6NQIiL0iToofX3NLx5zAgmEgKg0oNNOK9+
a0NWysJ0/mZBjmYt3R8GqBh0kQ1riEiDmBV1Pd10L+WwCC2wePNZoqa9zcmwgxL6+yBpDEZAcOms
UagnsOhgHOPWdMztZ1uDWzqVNdRUNt66dLpwFW0B//NgE4U14J/5gYBy98i+JGbLeQU85RBwXxLn
t5VAx2rb0gnptgNPm1ObTuy3PEITcq3aqjlqRZlJC3splDXaak82C4jCebZVl3k24kEqsVuSqvK0
pXe0URoKkNAybrNZIHrrczerR9UFelUBhii6o9FA+oH3joJWTOq241iDzBSts+P9TG18ymvPcHtQ
ETH7e6stj5VCLfZpNG+PqhfYR0mv3VmIbWq/rW/eqj/uSwH+9A+xHslF6txOlnkBHwpRpIEw4k/L
nCNpFgy3qUhhEn5b7DVKI7By3JADulVrPk8BB95OwGFMuRpc82DTlQYlRogKg8URBxrOWDiKAI7m
RUP+xAzFtbtE6UYeBQTZDzu1NzMawkDU+0zDJA4iL/UXOHVeW/ZZYn5oaCB1qGU7WXq0O+Mn+6dQ
Btn+PpXsRDU2hjP++JwyXWmjdAlD1006G7L6tNr7ZWyQAhRl23S9O/o72sNzrXnTfjp0jqDmcj+r
OEMQ1/yJdib+tFv5QcMR8thn6AFYho3/2PtVq2grwl+Ib3RvINp5jHnbz/0Y9sW+7DO5wju8sPFZ
jYxWp+fTxfq52JzZd5oo0wnhICvTcYTDC2qGepU8xQIVZK0y622FRvgXdlxVedoIng9F/+fSQMj0
xCVWqVzJMN36dbMZHtVzxdnM/xknMTblBhglUqs/GhPKc1MYy5YzIzQ7sZ1dIDaMooz+DsWIkCZ1
tliQNSQGw4CUBp05rpDxcGO6G4zJFtIqE+emndq9H7+NIf4SPh53BBlvmWVnAZO2FlL8Nb2YvBlV
F8aCHNd4uFbUsWLfc6u4dVvoaDa8JdNtjg+0k099zXgUZe3ozErV4nuf48HpytElF5u3QQfQDlmm
sp8xcMe1p31mcAoQlZszligJYxY6j/5AUdy0WT/T+fPQY0HHEjpuVKAOyvWIApfyxrF4ONxv0ccP
tXrImuqs/CbTfzENG+xgX1RIqykQpCRRFaeUT92BN4r8Z3uFwYSgwOON5bDvh0Wzqzgh2vVEpjTK
+ll4vUcuHoNtAKaLMaLdLyuZiLzT5gk/4byCksgEeolqCBFxo8B+CGVL4qX/iXFNcHpHcibHaNQT
UGB5zKs3ca0SQIqGikeLjnM5QhqnnBE6DVVT49muMY3bHoz4aKA1LA+ESVOOfrTARmzaOd9fIsey
E57JqzQX9jg/39MhaRQhkRurM81G8iD1sTjazTVXlJ4juUyoV8PL3a8JJmyULvW9CcQeAFwD+CR/
wpfsZU03wjmrcZpbcg2BRwW2RSbnpCyT697y0E78v6KyvmT4IxoNtHIW6mz8YMEs/Hwti9xtw4DF
VkWXu5vooD86BRt/keD1Bym6GBLRsn3pIPR/GoBh4/S002aRnJxcDF0s9sETEQ1zGQWYdqej72pF
KRgPQEyIYvYvOj+e3D+qr1clPUH92kAo5iWd+ilgWIl8BgsDdAv51J8/8VsZK5veooE98wXGB9+b
Zm7FwIYLBPDWWVDygTkkQVHjNxlwnBPN7fykzrH2sl5+UE6gU8C7WWo97X6/TKuRQcp/uhd6YKL9
XLg0uGS/jBK3kubB0ry1rkUSbNuT6Y5aoxU+WoHiCqfNVlAkMbFRw9e84K02Ar7onGN7dVhYkQa5
3PQyHMPMX3rN9zIfN/3whAq0V8PbCF4K6UHCjeb80sWZqRteIPUgJaJolMEFJE90kc54Qp35N5Hj
hYLpL4Rsuk8SnvRwG2DYTrSZfVBzbPrMzShwJX4K7ukadqpvxWj4/pHRv3k6f5SaieKnAQCV0W9V
c53+LcaUcq4qOL09pAtIDElHIbc0Xh2vqdZdmuJG6Xhmh3tOT1iV8ieNNRjyBFop+l2xgBbxlP8Z
b9qmbe6UvuoZjUtpcid0ISOOlxWZ6twRjZ9PEIx7edchIz5EC0j0PoFBQNY8nbzEkV/3HkHFfRe3
K4ErlMaFMZTXvwEURaEs6EB+HL3IiTjmfqrxW89TIMQWBjHvxSJkZKFB+MLF7U1lE64ugJdyicch
4u7TOjJawoV75E/MdKWYo1dv5X4a7HKb8vP9wD7ErW1ZAHF8rHoC1nAgwU33f3rpElPJHy7JVqHV
mPDUUm9cdBCTtkqo8JUCxyez6mq7WZMR7XnVJ5pJYHpqXdFqVGctVcjsngibvypgeb/ilrX5VI3c
cOXXf2teDNCQSOsXbj6eRbVVvYM1BtUmjUMLIwHE5/obZ2FSEqwANNysQ71NIOSKN5RWVb6KglU/
VAlnn670b0w753Tser68imx+j51JrE3nWHCWT2D2PZw5uapakZMTPfZ8TabFMpWw1PCBs3y8RagE
V2YE1/SONZvm8rcZZvJKHb+rhG0qbliv7KVXDFvFi2LtcWCqJvIaXzR+ebEQwaCF1phwBTP8HpCA
Gbk+uSHz9uZ5L13ihZ1se0Buhmfqc5Htj15FSFv5s2Tyw1YYcQ1UNlaevRnhW+ovQ2C1d3f7snbO
mNSIcGY5x3K1ZZhoJ9KuqvGtayXQLGYS/XBLp/I5Xg6L0gDXMSTsJtvtmRTUd+FFpfuZiqr+OSGA
4KKG/blo+YIwDcflINOCbYwL+xmN5VAB3ex6/5qMgWTSQDoTRBGr5mrw5dwZPt0mVeQAzHuOUPZW
yycBRI5IxGmZWZVbaOOfTRa8Zlj1wVUd1ollKLvR+9+JlK193ADBRFqN8Fp2eFIV+hCtECiwGsJn
pqBXwJJFmXL/ziSs2skWfXtp8xF8dTtzk62ixcXMINpbvWqDu6/BfwqHRjitAro2bQooMuNhpHgB
KAxLDNenu7LB9iP7aRWQm0oVQQFglX1CLihW3E4H7tAFylwoENj7/k0tkprJbNVWca8NLpgtyqYj
D0mFAP42F4EMXAInY7P8k5u5tVgZOF6p5heYmN/WGyk/LuQLb3YzX6OXE6G31moFwn7LVvZfTVHu
uc+RFVV+uPIlhXYiJdNs09I28JZTLUjU9HGy4AI/KpGPxb/1MeM2XEHf6B2QZtRYOigtQhnOv1z+
cRE7RWz9mSzkqH3DCJZuXJT896L7a4zGcK4+z9jKK+AyySlbDSQI2D1VluRcalLc6U8lQAmGMunb
FwOYMVUV0cqbmA1v8zAqwgfJyCf5kkAnM5KlwEYHs0nb1fpIKDOIXG1hUnK0huYZrmbDQKz8OO0o
RjkCgYdL1LFMmD73x7LuzoQQpdiD8pzoKdtFOvIauZn0tYUr1NdTQpmvl/DCOAaK0k/EssuF1uCh
Vc89CoBPxzCOdBDeeSKMNzN+sBmifN44XwPMvenXRkYYmN566aVx7n8JintTLpRWsgY80KLNTEQr
jKaEWSQ/9K3tB85eFBheK9VBqoJx36ayLew46Jc9hKAPhzFZQ8ok9fUWEINRU+kxVG5WoOkkq9s3
5JbX9t42HHJIVt6D+Sphodf3w5zBpxnpEDUbgm1JGEZedfjJ7lrCvlP5YFeBgW8JKSi/LsAB7JQf
LZ0QCjtKxuquMdytuJCSfX0Ohui4Rr9ru4Mqmqs8w+hc+0ef0KFddgnFlRYhvI+ilbkHwoQo8dd5
xmUbwHNCdDfnrbJJ9x2tn7acv7n0d4vXHFmJYXykHCAIbNIKm4LloT41ReS1gR2LXuEWcfS3NXKc
N1kWHsV4rze4TjpvBhA3nOyoClwOhq/EZXykgf+7wtEI3zWkT26RJaPw+Ndf76nSax4NOrSnlTNT
3AH1ducgNH5SHhCls2vGnM42ph3viIpeV41WOG8c6LydT0BpbVNf0E/IWWpCE+Ev3lXn+R+M9eel
dlAgT+wdFdYYC7IpI4lnmI/mTzZOS3MgO/SKMXWo0dStjdDAO/R7AIOihH9t9I9912Q4L6hplCEn
5bm5WgTVr7MVEitIm/4y8O/QpJENX9wPC6kVRARefAROA+LnrbC8Z6LTv9dzAE00dj0s4/gtGFhR
/qVQixf1nf45isac2Q7vrVi7taKQ1/WX9Q78MJHDzxmdCDAUCdfBC20Srrk97vA5HTUo+9A2DWxU
UdFq+HjiCKC8MAMgj7y9WI4Qdap2/WcEf58x0HjB48hFRYHtQlNadLaK0SrywlC4EWukCO++/WMv
9/Nl3M+J0QLmmoUuNzWeLrZzs7WcdeAxIm8TqkMQa0KJYh3YIHiY8kfzViMHtpnAoEks5nRQEtiv
9j30XcvmMBl6fnnZGONm6K75G7RvRmv+QcgzHNjYvfr/69H7ubHCybFiard+zacMAr3rmSup+BnJ
71MgTJohHuRjJKngSPaYFexp+qBmwqTSIS6jsq1DCZ0GhSU5vL778xuKjVg3Lp8maAiC344VVEc5
D6B2v0Hovl1FbRkBhTOxW8JQ/uwMkMYbqLw7xrb42itgy0dbtwlcZqrrBN8RsCRiOeB/kXA6LvGV
3ewx19ctO2N/6K5ieFlKa6ThyOkafY/fF01xAKc9y9nYZcglRrBs8sL3BWLdQ2HXpl0cveWfw4Ct
cGVR/3oqY2QOghcQKpNSOwM9XxKbE+eRfgkoV+7O/IhuNXbKih/627bM0RcyEEX3bMtYDudYlIN0
v1DE5qLV3llmmR7pRW8GvZu7YwN2nuu71WeVj+OPKyncCAoeyeT6qR3rmts/NenpN8u9u/U3svsp
nCupkE4lhu7Dhf0X0ZvlhGyfPxUS9ExclYZIFN++fXEdhfayDYOO4jX0orqBOm8RbDxG5P38ep6s
ibIBQ1BQFZxTfnWcKOlDGsyEZTnmsCOMaAe9ZcxmednFfGrTOADynMwxpZeJk17KE2Uzbloy58h7
uR7T46P7I0Xrh0qXeii5lR3GRyCtiZYK1v/cj/cU4AGXdAl0ekAbG7BnggyoxAL/w4sSPvGyv5Ed
Tw9mu1vmUWPdwIo90G5XyVoLaNkEwTSyETNjKPNVLJr/qN1WIIocrk7ylUcsMeAPkgVsN0dnRLtW
7iC5gH1AK3jv5fW8ABo+HQQcFEphhhA1Zs+W+ip33wHWAQLKwG0clsWLBcQ5sCpIfQhivLMMYhB5
Gvtukiu629UITzBh9dXpoFIdYVBHKbwGGcv/kHiT1v7hKuFFctCjbl2iGirmkO3obj5mg5aNCWc+
Hdn/RwIhJ7ggir1uiS+Ms+0r/owLlE/37u4c/jj7ALwJpOnvDIBka8HIf7a5tN1hAG1i17JMoFVC
uMQRijWFIWh1P23iLMLB0sdX5IpJb4O76cNXp0pEfWxJWmcugabXjMit5SS6bwws1oz47AzPrqfS
Q73qCguKeHj81DrD7j7imByevCbP/pZk9Tg1w0G6452sTkHPfatDZyOwAe8AtVsnR3PEtnzRyL/Z
Oa7ujW07PP1CiRKZWWGM/xVvwwh0AHGpZYcStSqLlr2/EbtRYi+j0+Fpl7m+gTv68MnasNeQbiez
G2SEGU2UUTtCyADLDUK0yH5Eerdk3HyWKs4ZeBkWRBkZRrlWuem76uFmCBo61IDa3OcS6nOE9rYP
A9iQYm54h9w3Oo8k2G9ITJ352KLypqyMAd5ZRLUSoM66qUKHVrpeicvT2Yf/GWT+MTicCKJIwPtI
EVCJazZVmK0bto5DppMT+SDZhQxPena51ZTUlWopNy5Am/P9gtxGVWAYsFqbEyC/VI6lKKuKLuFU
3/zbcutWztZ7lNXBVaJq4QxgFrrQFwlHCyCRm/AMo8NqCnAXnDLMXnvJ7VMDZjFUj58pbr18XiUl
0rz1Pa4JBEmMUgdlyq59I5nOT609lDeeTl71VvizpuO2CETvN4QTC2UWi321jnLqmrR2xUSP6LXP
UHCrn8Ew0J6+bp4g5hESYiN1KSSxmVywigrhRqH8UH/4ccqaytvJKQaV3rcej48CdD8fJeoISw4N
0ehRLkhlQwctqm6Ro/BrY/pgQ0ADMxKkcAV6ToKKh2vYP1GRsltzgbWo5qnHMHDOlkLngnhdKzkf
rjp+6tNgqcG+v+zHOKaW1HSNGf7qvdfxm+HAXkd4Ts/ewagZWghi0bjzNxVb1Y6zf8DRtrF7nVi3
EJdzYl7+IoR/IoNYpFcyfwIkst9TFiQmXuurKgaHEL8cqfE07rn6hNdDUyOASRBsCZ4A23QDMlD4
nE7p/uay2fWv25CWgP3RVfL3p3jQIPJdKAVb7zoveOhb//pGEXOi7DIKo+7FTsOYF8Fwyzfig9hN
TqIWi0cZj50eDfyGvTd4uDjcM/i9+hODZiOxLUvA9FWADDF667ffKxX0iFst4WUC9yG+VtU4x1YL
Bs+Dn9/1oakOobaChKJrbK7156vEabkmzdpUngACxDr8w6j91wvUD1szDnrCqAlDbYSmgo1qKuTM
wYSy/OY5Q7mlndwSKT6rx9NVR0w7ZPRXmiLLKg4X2WxLdf0iTQ7NwaI3PAn72mlYRx5ua+1xUEzv
YT+fZNH0w01PURiiMpXLOOlSqtrvAwcYpFqA0nHl3V/oP7FNCUDOe9a6A3IBCasrBfBOk5zarwxK
LGBrSNFdZOX+IMOJdfQ+hmGDOo+EeMRR4mXGFV3WaHzVqLoNuUh27LhFwOjoQupr/vLLf1Q3XNuW
xwptf4IQEUVGEkWRomofhpKo+WiLYpu76QuuDcCyAe8EG2yMjuBQ5Rrxx/r4etk2q/9d6E0ESfqz
S7+0xY9hkoMMNJAGgsHYpx1KLS1/uFq5P/qqNE6tFxUJO+GrLkeN1QsFjmXzwJ3znCbIZyJQ7uGP
p1gtdwbEjBbPTjsNdSk0SwEbHDfcEqlFO/55Nd9yDYzkgVLhEOcL+0ViMhmWNEMtuLdcgxE3ybHm
eWsY6B77vFQdHC0YBvKyRy0qF8ONowoV19VeNIjgnfpYbOVdec3ctvXxXhberOrTt2yEbvcf3Eiv
fNfM71MiUvq7PjplByMz2v4wzVni/AUm73dALTf+9rXVdLKV+dcxQ78NpdGjo1xaE8CmfBgcQJYM
uvJClGIyYerHNo/+Uc84Z80nUAClQNfwu9F2u561b/REtLTA/gLxLl3ihzXl18T+7z34UBVqdzTn
dyIMbdyZ2rIFxnNo3/Am9DaaRvPVkcIHrt/C1SqleHnKR5Lj/Ego9tJ2oQFNtIoeJijz01PDi9f3
eg0DwIdmdQBxx3FSbn2l2pNCknMBC94xFR4Nhd5OpKuwu2S3wifOt4HidoKN1hMrxD2VTgM5Nbsx
VKMQwgy7fSldOB5QWQN3h0vtb8QHImV9meGfOTVghO1Lrx3OJvkmF90jtKSTeeNCg/liZaAILb34
VoUfjYL//+XngaCfNR6pZnz1mpiCYbhlg8hzIgCvXdijNDShwxhxRL/QQxJ/8/VD3Mkfht66UZtv
OqX7JE0NpfrO7pi6SAj5nvlZWVv+fHcnL+cjuFkf3wUMss6xOckTNr9TBsXZBY5GvQRUtX0s20l1
RVhOIT21QyDbd23m9HcVDvhS2qEqJjcHAbKsppwyPwfYFBUqz4DGihEM9xdnz8wlsvWsuAcnFB3W
noLgLX/2YS/FuUCXY7HxqVHnEfgMXHVaQ6xN0XVWa2fEkg15BNJjL7P/lZNgEEPUIhokHOO2cTb/
VQ0JZm1hCyM8KyXGZJYwIQNNztdnoKWPWP/qUWG0umjVct17jte1tKY8vdfHK4xj/TWu4XRqhTa0
RKcJpqR3+QEpZGo4bVkIugM4McbzaUMnh1ksuXOIpOKEDVK23a4ZTc6qJNe3gBG6xT6Q6BAGmn+Q
idZ/q0ELefQA6ZJ3E6skqSgNIlpeEJbO70x0FtcCjLCnnhmukwZVcRplXOozJXKKmrTpn7wRoBCc
4LfBGioDXzE4X6VlmovjgtzRdoGpiqSfiGa5yf1wdQQKAuKgQ98+wxPMuFQbrl/YKxTZ2r+nQKh5
yEw/+1RUec1nAST2EW/ch939InMjLiNRK2bNcV4FSmQ+Mb2RVmCJa0eS0DGj3+doC7v5vE3Dzs99
wiN02VwG5hgA/aks1OSlgO+7USMAM/UzYQhbdG6GqN+IEwF65IByjzX2NRcY601Uh5ZFnuKyCmem
S75FAfcMm7okX0TfEPKGjK5R3MkKGW5qlvuJ53QoGue+aPgfbrBOsVzVVrDE45p6xdwJFdVoCd5m
l7DNzBjOSez+Me2Co6vHmkU5pMuTwNyFVyDgtqbqj5SPsu7XVm5+SG7qqlN5yQWJJGuNBBEVbzWd
BqKBPUdcmZiAet1wgVFqVHEoDKeDr6F63WRJzSRe8NJUVLQXpRw6XiuHyBtc5pOLu2IsnmzFqqth
bRHa0D2ytBawLl+tB21yNRfklNBZDXC1NI7OBpL0NgSKXTSsh8D3CJBAqLLFYIpAAAzUSiTMYLO0
OTN3Up7lYdZK6p75gVmGjaPB39nAUNcpY7JnXik0ydPoihbJP2an3SVrp8kRaGQDSuyoDF5LiGZS
i0LbCfuQyEH2p7X8OrbNL2vWEus3kzDaAW60wV0sVEMqG1dPwQpzjCG0tN2qiWG1ikrfs3T3wIhq
Tm/GjHYAUt9f8QtyyBFZYzXbQZpoB+pCvZgCfkM01Cd9AOOWlvsdbikb9w/vJTykBP/9HAXYWpym
/R78WaaJp/NEBJr6aCtrnW7T0GrUuYvgANWJs7GnWpLx4M37e+igGSvCn4VkeFDstZCUuWtkBBQ4
pz8kxEeoQpZffJW3kHUi5ePaQ9YaqJjPBzIP6am8xdQK6IghdO121/JCfywb8oueyss2rdC8s7kN
vWXfXZHLxR6VieHOldVbAc8UqKWNc9CM0NL0W6h+63xHS2Hyz+JKNJNzDUN4RNMtZheX1vh++7yI
s7Hre0XbSP4tW/sEn/QP0u9mE37RVQWEvosuZqzSdT9u2W3uajVk9eP2GqDkbpLecuW26PaX1Oqb
PgbtFXICxPOZC8N9ZuUQjxkF5QHJS7heZQHRj81oWZUU3WMpxsE3t0ZzREczgDzm5+Pfv2AyRgEr
r9HiCFfDEUDDokfPZ/QuD+8AJUQcZ9OrrxFsZeEfmMoNGCogXpFly0gPNhYbW8h0RM5SNT+Rj4qa
M0AIA/aTXEwXDKGoJDcHtCFn0a85KNb9LS5qm0fIZq9pe4uYDAjODD9lp+7u0KmSPPv7Ftpqv5FT
m/m6AYZZfj4O0YWW7k0pOnxTu2mRNh1SYxthpzwGBZvodkOwfpleAVvZLUefULe/tIV73o63VWtS
Dtyfe41EVJPlCsKOIREl2vBWlxroSXOEEbB3PkVYkS9p3b1SnQpDDAJBC5noHBryyXX1UWkYVV2r
YqtetU5eitA4SNT7GAYw2Pk0blYU5y+iM32/uvc71EeXJxZDdSDROHz0WcySws5jEW6YL/JoSRR6
uEACyOm6EofhFykWvT5uB4eQgSJTOIbcW199xr9sKoPpwB/kpzICLUvsa5P4MEfWbQ0dMs5Uixix
VibKtpg2zYBKlOsHdQwtHSZnCypkfNTzehMno99RjVdV3I4tc32TMUpPNbhc1zlxQdwZqmqsmfTm
HJr0G9gu/EnOVg4EYZYSypZ9E62yqu00HY8lvaQoGYco1qOy3xXQ8XrlI1frgTIcXZvjREK4Wo26
zCjv90DZqI89VHHrz16vmbX8kLV3Pn3Gp6rZjKUNUkarvyOhtrEOYiQoyHQ/uOwtcbR12FyJJvze
5OLMcrLj4MiLIyghsX4mLjhZ2GdG4kKekxeSLaLY15nZcoG+zzd+quF2CbUClsPmNNVFDA46Ezua
OTKerbCSJVB7W4Lv+FX2aWu8rFJhcp1PlRJ/YWVqn+57IjOya4KRQg8AZYFqlXazuPpy7DeDJvtN
Ft/Sf1DTRnFbwhOckWPi2X1u+WWCJABLgprzIUECbUjmGW7InZr2/Hg/W/YchEHxIy4lHFoIXaIs
bIDjhSkHi983AZdMmacClnqFnT7kzvCaES9wrIEcHrHKsm1Gi66PAcvkznKimq4t2mNPEcGxtvAI
4Up6nd4a4r4g3+nmDb9L4iD+NqK+3wSrvVvWfEhT0H1VIh2cL1qRKZF55tbamLQJIc3WMYhHxUwp
kyTos77K8Siu8nzkgMXIaFNOIlP+idMXJerzg5fu6ZntzV0PCO8kMLDkBJMAGI0/KeUDeT9WY1iM
6jggwNLKQb6FZei/CmS7jfeEchQNbGM8czNZ4zUBbx8tWQuFPu48EcbGhGYAvXehcQlAiqayioKl
Gqnbv30wsbme2MCY5J1w0jdGhAOdNwbapoOevnfw0nz2Lia7sCwWU9Av39uun//doz5b1buOaqaw
LtJ35MeN+1CHXwNwl+ft0ZoDVgum4GOtY0Z0z1rZfr+3R76h+Bek7mJiCxjJzszyvSNQ/cTqT4mv
rSAVCfrNopbfl9nhnNVvYODZheEbmN2yN11+KZIDSqyRnEiDIkgTN7WwMn0FQk7pgUvsA/GGE+7Y
3Rvx/TlStTMSM1yY41/+ZzGpTdKmgB0rvG83Yn2gxN4Rip4NPuEc28r2N1IN6T1lcEIec36tsm9N
2hoZ7igevhD80jKm2c4wCw70rOVoBT8I7+mBSpLtMgM1Lj57oHRYiyhrbFv3nb3Rr4r/raNfhh6Y
1hGQArAcdp5aLqlr/aKheHcdtCVQtbSXUz/QxGFwwsZcSovRdfpY3IU01chtxXXdPenewtgy9R5N
8GqrtylWkIeCEaH/cw7stCtnJ06SdqbEPwnLldUyem/h4vi5IEObisKynhUSFlAbamzsQ0X/NLv9
ECv2cxJE9YyY0l+WdsyCb4bFSVbMiln/S4v+QQUajhmsGqqq9dr5jQOuEXOzm0iURXWNS5UfzhrL
VnKbtkwwqQrdQzq79yGtkKPV3LKyco87disR6rupfKT3tBiLN1TzStt6oW8kwkTcaUnEjq3iqWdW
yqyhI62qQMKisd9hxj8TS2CNg3+GKrQhD1H7PdlzOqBHj1R/vxCxBr4QFBxsqH9ZjdFdkVWBsl6a
owQnUULIjlufn0pyPSUvpKVwXSt3SfeiC4S4IWfRzWY1WwKMgcgZA6IrEWHvKAPEogG+mkAdinyZ
RCNI15kuz5GY7aArb3TJvpuAP/gA5RmoWM70EUf/BFZ0QfasoEPmLXUwthGJkzFB0I/Y7SCoOcd+
PFuBy6b7aSzhkyQRdH+P/ttJO8nR6a2xuTgDY+sZxXN/uBqC0z2shj1yMGZehLmg9cliA7SLSpr0
fRFYbbkQ0gV49iNfI35/jWVqreQhX0C3/2aasCjYV7tJ3oZO86j97aOcjA1D7bIDPI6gccm/FPed
QqKYqEujRn3hwp5O2iPq5Vxj+at75GTYbtaoDJobv3ZShtXllSvCdhX7yxMpT6h8QoJAQedgeY9q
trk6LSqBeO3h2l7eAzdmuQNSotoHWuvoUfNcTX3zldu+q8cw6VRaAM6QOJ7eg1uQnoRCOPMhbkH6
zC93RAPkle3cJcG3Gm0hgS3S++fV1m3cPCIDfvguQBzwQG0HdRsb+sL7K6qgVe6QS9gpC4kY6TEc
SU4doDC+gNIagJCFjudFHSMWTGAFeDtWJcjeffbfgz68o/KvG/q5vtr4DyXcSg4vw9fRlQFCE8rQ
SY5Oc62qyr0ff2bfuKrOh7vT4KrkD+JljYYQXBRdyPgmRKgVvl+SYmg6AqR2mDyKHce0Qn3W4LrG
/g2Zgtm24E40pzSSdI65VYhocY74OM9XuuA2kdbcfWFWAnL8by4sqq0wMkqp/fcJSXn0LFYpbRbY
7T3yHK7pNgQNnaFzsXcbqUog+pvUiTje1n+ThIQwaaJHVUkCCAeMEyMt/Ad7EHDFHmpuJxmTLqU9
RVZ7MstSu0SljNGk7WAROvOYLf0NUsBpTj401jbbtIKTonVhEANowMyLJeS7z1Y3DWFQMzjU9pwX
9sCXZdf5R17R4mDFzZbDGB93l9Y2+MCOxl6P+cgjNpKJwIqswYzO+uKBy3iTbQKL1ILSVsWdzEYw
pCPGCFWL/2bDibaR8qiAmPqi92DsF+7ql6xQWpcsx4S4wEqrjbxes1syczWFBlWxYUrdxnmzKQuq
+Mrt5t8IIY6WrfeAPP+Iv3Y2qOLONMltRG/lMrtSocEK+4enU2N7vpzswLQBkcrgypDaYZffT5ww
fKePuTObehCQIJYH6nBHGol2b2qbPg3iUyPn9k5Q9ZOzlcqkt6ywbTKhg5KA55IH4Ac0GHCaNkEs
h6KLo4DpUBHeBHlSHRGaBkSIfc45XClwjrk6QwzhcPgujNhmGcsFrvzP8DnvFebYFDaJ/KMFfCZG
dKaSJHWE63/S9jrNQtsI0sVxzjn0O9cO0tZTLEWvxOq0oZn0AbWZY+X5T75KLAReD+4D8J/dB3UY
3NhDgzzFOf/2ZwIZh/xNRaP1+SRRRebDiYq2Ef+YE4YoYxe6BF/fvpb2gEiDN9wgJz5zCzXoVune
XhIR3LlG9OFkDhWNDbRFbDw76YAHKckTouD877yZNt1oQxomx4hcSGF72oIyzwcM2kYgTrYki6EO
FaZawxp2fl507TYdgRN5hpbbSAz4T2o3g5BcE2bQZsG08pELKeVRpE7MGg1rE3dS2pjNoB1Yc7m9
QWQFs5ULInPcj3ZwLu721UcEpFRM37VESKUn9WDoVucolk+Ob+cVnw8duDbyE7r8ysE/Rkt3Fmg9
dQW3O/XpmBaCXzgGD/3gtAd4fxpALLws6Km7G8FDx7Od1MCmxo3tFTjOSYIA1qnWFR8fwPwSRMaZ
2bHaqKR1mAfb8kCbrjMk+CCiw1aGU21uaYB53EobhkVzjaKvARZ4b4cwvZdjfBrdD9BfhXSITsW3
h9tyhWrPmowCHie5XHXCqsF1q/CETrZFovKAn/Z4lACI0XkJ+qU0ma/5j3dm1d2PFWVSrQxKjH6P
4Y5OM6Xwg46Vs1oMb9zC+OjInVlO/ZEQYDsr0h4vwohGi5sAqkLUUIR70bWJo4xrWgEe9ZxKvKg2
+oAhVcF6z0B/8mvjSjVAmm92vQHeqK3mdTlTrW+Xz/ooxJTg6kwCcN2zbV/YVHswqstjqh5EXCJ8
b+6RH3M5qjmoHkw7bm/bILRyX2Xymz1CgNGbRDkY66GB8MzyfQn8kvZ+3Hx2Vhak1wsvdX2h6N6I
3rvYsJMz9i+tByi3ZAxklcvMrUkG1xbCWsMD4q5OGPihgvZClV06FGTYaMeKFXs8k4a3Eq7o9LxQ
iy27VpbDnU2FAKE22fm+SM5RftnDubMB1DZZDu5nTsyWxnkszafjPy1NgKF/cCFjSxfnGFrod9eV
3JpykDflxd6nAQnYilRA4P55HA16rCHV2iPHddghw2oFbpDH2DJNl065t+4NJVmux8OR4FCDDAos
fEcPJ5Qj12zqmx1OhmzLUHSTB6AD0cS9YjIkSVcobNLdZB91kQ2x2dwAj05Hr6UoXsuJCfPGgCru
s13kv2PFVvkLmbGo6OX7/rAlQl3C7ntAw6hBuUyFdU3oIpu59uuF53dfPMs05BmEu9wo5qyYAoKR
DU6LJd+hQUbJSuaY2/QRm8H/rHVfNtykcUdHeIK4KAgjIgWJY57SjIl+TEpWx2iymWBMQ3Hl7KAQ
iOqzzLXTkTd78ezQkh8rgq+lOs1JOOr3vQnXZbaEojMBg/tILQbVktDM5cAL/m7sMXIch7VK5e0t
mZDJNQCpWvv/LbqxFA3xRypgDBCf108s4R1TJYhgeNv0KMNSisSN9K6cxQv6MzqNe906JPPXbdjB
96VPJMd6th+mUju5tyaDz5NZXywuDiBROxk837stnyzSaw76NYzS9KJCo9/IxxvF1fEcVdxsTh9N
QfkcoMWsKgECKfD33jg/VruhoEyiPcFImgGuR0dzwJVb0rUTTLssWi674e/Uhyo7I6vAtbQ2ykc1
R/tdTzy5PwX+Qs0JMl7lwwqbKIb3AEmP1LNaiCc5oHi0SSO1hsx8/Ng2tG8vPRtMuPWhM4U8mhS3
8hzqs6186tipzGrm9MRyGENEBvrSs9nu8/IJcV8gUFLp6i+uDeNSWAdQwNVisIx1zx1oYLtKqdlR
s/aT90mPGCdDuFzbDq76nTeh6TxfC0+qnS0PIq3wcphSGov/Q8ADlmirPmSmlnuZA4MQoWlOVYrG
cqYjjYsjHw3YRF/K5EioKUVsSIutkx1qFonv1xUH1bTMk9tPWbXxmftpaNzcd0NyjyFAi8vHeBJd
R6RiJhS+ZhUDiD0+cpElGCCEqCDNqcaOG5vsBcbi155T6MXxAhpca32IuwxFAyogCIHVuOW92vFT
VTFqho+4wbYgyx6fsc2wZKwSIjCv88KUeZRYGdHJS/92fTMuFRNPrfFA6w6ne75ssEZsH6WS/4Sk
LPkP1KOwChhdS17dKsS9QxAguo/yPESMX640H+mflzaEyg4Ng3hieNhMl0zeNZKNnTj7ndx5Anek
4qHjvi709zJzVb6zAv9BGt31pwjldj6pQDmj8reEbTtCrDtK3lGfv3rsqQ2dyemk3j7d9sj9ROfU
b2x1TSQSMgNtCBuesUUwPx5AtY1KARHYW80b1wybZSre3eAuhrfO15SZ/cIOfbgBbdYuofWPW/pp
eU/ATxNQ5K2bQZpDvEEVPQXBHia0xTlDsxg1quhD+zBtBgQIcBUYNdJZvJZXC1XS3AZ3cM8JJL8C
HPgZq0D0wK2uDYTnIEufmvExBsfqY+kK5WfZUyvf2O/b0GMLlfb8k80CXS/NWdmWvsyq1x0KANRR
DS7YiEnRZv/zJ8PZXFi4Zqm18fUxCeMYIIE9gW6w5ec7eY7UPKbnlgIJZORlmgDvQ8chTngMzWmQ
WZThV+DOlpDBaenmSo82cR3DagoR9dGjs8oIaFSi2Mqm7L1y54yx6qT4noUhB4LI+ChC5QKKnJNs
keHn+HNqGj8DOXb1OG4ISDgj0i5PAHRKXKbvSKGpGodRlzjQb2Czncdjw9hIwkk1+TK3L/ibJ7pd
bSIZF9Sooch8jv/r6Tgcp1KjqXMskignECOJuz2JCH9wE0ZWL/b3R9hAqcbltsbqvOApQYHo61uk
naYj6ag+ZrYjHop68gggiWAvFlN+Z0KHzxs3di2QP57fxug/RG65lGOkGQtD8Gmu2e+m64dlhrua
pBYeVhu7L5qX41IXIbxAg5uWLVP8FALm6RR6AunQzv0yORAXEObLMNZwQGj7l4oijroFAYwXC1OB
FyiCS1IYuqSr/pDulFmYioTvjFE35+rdyGK/GVjcSPVCDwparN1JI0BkqDO9CDQUm9Fn3OujTPhJ
WKpgFiRRz3NOldO8upZ+KmUsquXAMXZFcrI8qfJX2FhUog2DjQubKgu2E5iBuavtrQ5J2NqiAAyc
oc8DkWzgs67K57uQ4t1w1pOY5OY5pC7qp9u/Bsowe5uVdoYejXkushigpc9l2S40G5nLnt3stkS4
42IOggz/6zpyPxuZUMNjQz1umTwFWTMvTLs9wjBhG+f8SIqvgJAFCLAhIt7zSkrKbOsmHu2BY91+
6MJRLQC3Gypm0ur/rXycnb6MX05ovX7iv8DBfVB2oGyrdwFrd92zIqycS0b1xnfJoi1JPI0Gm7VU
0SLVphjabt47EuOFOK4cCVMlyf5ZmOCYH1ivoqX+1LXnzKMgXgIlh8ATcedBBqtdowIewa406/pj
B0qP8OhUs5d2vkX2HY8PIGx+0gt01ut2hyr8xuG3l+3hILssSqr86IY+rWkzKg43CS3SWAx9lDJi
TVjsCwfO0SxSsWlsyPiEQy8k4vRbVUc3MQTJilaNazskRq2AUlNfhoJYoOwd1t5D7e/p7o97jHAi
H43gZxvt/2+laF12vJbmVVBZshl2fHhldXhMKerKywucgURWhMW5e5powHlLZBeh+6qm52Xb1sW5
oXsbSlWgTKHvoIJhHlXnLWTCsVPLu/r0hoSU/A8G6wFBAcJ7wmXLjBs80qtn0p73PL0Eh6Fp+S4d
2QMXelySJ1ofbkEr6eVMLJSyb+R/J8RunjHPdf3D98A3hW2C7+xEBNeTuQBkRxI+Q3JJzmBIk4s6
us/ChLUGMNebdKRMVI6c0cgvs3fNQJlES/KzcNNFIYtBEl586fKn5dkakGpUYDADWzETJsC7mx6V
hlVqpdSAjK3QJc0w/kTMgMD9NdP8xG1W4aggEZFX3O+4xd3kOolnE+81JwqjR7cM5UsWSBWAd1X3
k2tg8hG7MQADz0nIuY/gOgC6owKKANDgIg7NaFJwF1Mk7ox3x+DUMwfGYB+t3GGP9Yb9NwQLRtDc
/sprozXGUtOwdVgrnT7/QFpPX7cEksSKJHfrkka3OGJ8KlMJ2752HtDjzOudQo4B0cCd618NXGxs
4ybV2V8P5hbfJqYgVM4ub9cpdm3iqFr4XWbAJr7XUggvzFsnv2ghLA+oXxnD33vsdxXHq6qpIAlK
4XweY+7+5w/m4p1xde+QptMU5c//b0F+HejCR4wkG6Tkbt0KtschY+7gyGxAioTaFZ2rsTqPV6uH
1cQpJN2zCU+RQqptT02Kntx5m82T7pgTydgNdTUBp+E8EvdbU9cEC90owQs/8YZOLADnQ6a1p4k6
WjsB+CbIK5ncjz6B6VmU4eyWz87n0m9glfiQ9T1z0dCxRBkQTly2pJxns9BZiFtacxMsJlE9sroy
/CcHMXUuhovN0JAnsOw5gCvotswoQiEtNsGuTVwPLlJhMb0M3QFfTBWPDcqnRcNatNXnTYSGvdRG
3Yr3Ok22RyGBehxBAVTkc/ZddR96S/FG3QOLuoDuzzuMplxcfh8YxkYn57uuNzXXGs6rhXkp1xbS
DOgmZSXdK/4Bm1RXWQfOlhnm6ylRmilz7sZM47zD4TUq/NWga4jAvvE+CRy4o8Inw3NszNL9MQlk
Sf2wwe4QD6PcrYjdwm/rHnaFH5jqLNWuXy+gQFQQblxuIOCGpTL3xzPMavKMFhTI1+DExDQZZO7h
E7iVlIElcGjQlggygTc9whChSALLUIfLXCygDiMAPc27rD+hqPXphcn5YjdWmAqrRd4ueukUFd+P
ik7RndQJ7e1c81PHHZZML92RgQKqV+lEWdV5P9mJ8VQw8Ti8IDSeK7wuovXRd89+1OCnc5WtxU7q
JBI9blQC/q5f9qKnDabCCvDZ97hJjcNjJxFyke7L5QIdci4NTBFBtUntVgP76OMAOS3V0Jt9ybx3
7BVKRJQVF9qDMeVS+RMnjTub5o0p9jG45ZHA0/dAvlMFY2lbZLaMqon2Gvrb++MTyM0aXm+tQS/A
2rd9jgXb4p+/tPnLzUyQ6aLEootFCivMv7J5ybV/AS1YD/vNTVptpwn0pzHgoED/XS3BiEKa06J6
vXXxYKaWWYxU2SdRFUV3Cl7Apyg1gr6NZRq59c+O4QT9suOCNRS4s2A8NU2hwQ+4IoAxIG8Bcjtb
04+dVH3GhrwXY8zGamlT5duJces5+Pyc8tsl2vrGtKN1VH7/EwrBrR0DwzXEdbJgUb01q3HYAN6Z
HUrNXfSaz0fmHvPoqp4Dfc2v2vJ16TmoBLNQRHqHPW9hYXuhA5O2SSFQnFTYh+oudN0x3fQ5T0Y/
ubFQzggYvWtTZwKMVQITw2uxRV6Sxaatg6apXwz1NHTu4zBGbbcHuQU7huFzZqnt5BPY8VImzn6H
4tAhA7CKf91YcMe6G4YzVJdEk/glfdTLd1OGY6J7Uoj+lG4JbSD/asMdgi8A2RXZBBC2Qv5K5qq/
8jEzcG6+wTerM+z6Yt+/Px4HLPI83/+loEAhWsr22pOGm5Kd1NJ+An7aGnb4VJKf6PdO+QmcN4Ws
9/ICz/R6/v2a4namH22tH6q4Oy6nBrUV4ekmSRfMCK9fyq1bJ7T14eCDC8H7PJX/gRPB0wpa85+n
Ejz3ideoJIWj4d7kqMPBIm47PECln18vPyAPBmjbMagyqZW6Pqn+VyhoiewjI9SoKaV5AQ4zxZ77
Q2iNhNyUThjFUIbxVZWxrMou0edlr0ioSssZNUW+ZVtVX5PWIYDSDN9h+X/6hp65hRj0RODUb3NL
BxAkU9PEF+TzsaBniTzrvU3OjW7uPaAPy0RmIoaXfFBXf2lSBmA1FvtpXswqu7O1pO7+n2162/mY
mV/SZ2T7NPUnRZao/nDPyGmqGLQH08V3azmXdKr0AGaTFt+tzMrBIG8tCGxv0dSxaZH9xNHwkeaz
9Bvh1Ri8MPDFWtzL43pSNHHdtAvshs3/t+UmQmu2gOicusFCHWQKDj3LBbkGrBzVFC33VB/YfhcN
BlAii+Cv24FXzXU908aqxj54zISSNPr5C8RZVfbCZqB2SzK65nZcBdjeXJ8Ro15vzIsaHuM7I5yS
InEuEE85Wg3eh1IjR9mb468E98yVQHffB1hPh18g8LzchBC4rax8atsqmIkkIfAcIr+XQQo2rGIF
dr7W2VWWHTC7E3RDKo9Axz7uWY8IAVDshcnFO86Khtb5fpqlfct+WTqY1SyND6GsBU+ctxrWldBZ
hfpT4KR8JNlnh4vyw6uBIHGbo4e+DhnT0fLA5dGmuQ2XWbB8trOGfv6SnyniWx+ndN+cnL5HmF3h
PzN1ueeA6JwQhy/vRITAllnnf29JJnVpC3CQDXiSBmV+JMrlZ2yWhD8ThgMg+V1NFkQfxwOcsZPT
RJiYmwT21j5U51624VFU7Z0865Q7ivcwxnB0j078tk/23SUbnZ0wvRw5yjc4MxsRdSnvUjC8tXj7
pVcGU812uSq4PANP3t56ukQDIHdE7OPk4sr33tnrfIEaQJoDe8Eqki/mu3I9CWQE/YEo7XSFmhWE
diPg7NYjWth6pD1q4Zi9tkV+cngnwBft9MPEm+iDjSw6QWWK9tEKvAIhz+TpHGDfQ2ephiZLlWK2
Su5sbrBZ1AHnLkXgxxzHEJFrEpE+0llMhizRYJbiXdhR21G7eH9ljDq/wfQgA4HIuddHlKKfWULV
ca223aSSPGMikwJpjpiKYSrFIaIpXF/Bvs+fIBPTlXOhFhwB/+uHZqb4q1KQ9W4G2WYwEnWdWhYo
avu/lG9GEa6WECbMxR7cJVCW3YcVmVRRunhTDDUdB4kEDiGlGKoAlYlML+5pG2Gy/AgzVkFKAahW
IVSz5opGw8DoWNJWq/3KWKhQojVu02JtFc0RPTq6y7fGH6dZkWK0oAK/syDwEYAOwgwXgR9uEceo
9uR29gS0omD51lWHkNUABz+zFXDVq2YgidtmrTyPMfiUSj+dyaUCDGBz02hPqhiG38B6csdgSUCk
iUOxFRroCXRLLkLkeGnrlEdZaJy7jFoGBu0A8AcfVD+wMak+GT34xc6Gah7g6FK1WF0vC2beAP25
gv3ERsqJYlAx0Y3Gb1JPcyhdXlEHu+oUzMI8Vofc+F5V9qzd1c51zd6iQNrXSTCPt7PICK45Q2jk
TVyK+QVRZNEwQRxYBqJxSvGBvVK4xrRoHiAda2QG6X4uUlBblGs7ZiVewmvYymJmD6dEvWVFqW8w
+B3AwUW3Xt2EgNcupt8cVg4xY8gsE3DeUS5O0coJfX5WGaQfwcIJ8d4VYV6fZdvyxCRXXRyUfxZg
Wmg+GlsZO2OyiVl8BpLQQueEN24RcwSuHyj81+C/goG9OPJ0fyMdQyay8LY2vnAbOD7dRmoeEHEo
N4toxlBqXgTxvgYdv2tzUkgpRooEx4rEz9RaNvGu9gocYdIlwBKZWqUKollKSCYIYXkzOpz+ZcxS
7uPNuBnVpfj/Q2TAm/riW4tfsiLN4MRSp1qoDZgFAXIQVIt5E+DUGBOMMf5phcbHl095NHkTEVYV
z1QAqccjl4k89qGRtu0VicmAv3BJQo8bGa200CFZpI85hhxB6B7VFYwRKh5ez7/P0NzjLHE3QTYY
99U19vNY7KeOk/QZrd3e6d5b2gs0phSojOcKHMzLQSl5KmXUiJl1UIUHspQc6oJ3uUzH6ZNd1odZ
apGlMyh7dyj6/avvl8ePVjEo5H1KLOiuCiQ9G8XlbKP1FKRUzYidm9ZvgFZdgzpgPB6ItbdjLHRY
AyIUaTx6B/+Qx+Pp6o/i+KzxcvXQWxCjA0jmyxzKryVxp0flOExWRyo89Orn3995Uz31e30Z6Jh1
O/Pvf8ggZzpgfChiD1M3oyzRpHkbrh6hswNAiWpCfhSjSrJSG+LEsgPHMzaq4MRH+SFNzrWIENxP
bu+pLEOLcgHCfITXZk7Xx2HOokLp5RrSkRA2VPdVhUFrJDCCCHUHfo/WR6KOmYuyy7p0lRQpfBnL
6kaehn0oIwCk3WCpB7pA5s3sgu7Q3Or9NPoaABilloJw/yeZtBVSu1PiN4cmItcPhO8ozn2lYH4k
vxbZu7gyW0fTx8yMczvBnmC7QkIIl/5vRyBZVPf2nHPJdOpN5T2tsvF2dKmVHR9QKjRaSeqbKJEo
eYR6uvb2dt4M2eueTpmtBmX7QXHXIcToomzdVJAqjSDOPsImiur5h+I11oiM8zELFqjbZeKmXHJ8
XHg4Vl7Nc5eUKEdkCvBEyFZqD/VqKFuJgIakEHfG7CabZIVFRJRrZQKX3i4opeetjwSyIJYSFEV2
fJGyie93cStlThokegQMnKyjKsqiLUOBUG7UdZ6WlkUGWurGawaQxrsKVyHp9P4i8s/2oaiPg3m8
fJ7gc+6qbXHx/0pAOabkFMdgKPf+yG8o/U5Mul+0TSJvqh+Zmzi2CXpatLUy2sepkVWGElKYn8fC
e4DUvhhTjEsMT1RATtFe83sLqMDQfDd4ZPce44jT17t7qXk7cyu+gPxdG6/Z7j9PxDrjWQdylS0z
EgBgFQ/MRAG4qO+rr8+IPYa2A2FRrZVAc8JgSipKXxiWqcZtDQH5v8Ry/p1krzQ1Z7r9E1OGYRuh
VkdFFKsPsRJ6/FTupa3wrJNpvSTOXfKXmiFT8PdHAA4HwCYhCx0XFAJkk4o0rh2f+gVs/oLZg1mQ
gZ26WlTqnNDky8KCCr2h/myiRhtmkmzSSvLSwcvat6aQFn9Ah19YxfD3o20nB/6sjvZgOrOYGZen
51AoKMoqxF5Lsa9yMzCUEBSd7D4QiB/GILgu8Bvc5LjhjFnWW62qDMh8mn3SD3VHeUmy0d6G8UQW
ONEr/OWrpdBMbycYOckMTjcBXbTC1uJR+HbPJiBuTfOI73MtRKpI4YtwC70CVDEl8XQ8trdW/RaQ
kFn6xl/lE7QhNMKRF8P3C/UFRoOLz2WfotJhuKd/GgcgnFb8YeW0cIy+10VSvDR0czFs7Qyt9qPa
eUbgZeUMNy+U0zThdquAG0jaUbbgwmIh8qxMYqz2gslPrSnkN0zJOwUSS/wk2iz3dTgerSULE3c5
zx+rJQdfMQFWbNJzC5AvUeBg+iUVM0o5Vl1sY6oS6Al0o6HcArkkLYYzs6O83bsUDYKlW05g08g7
wQUlpqLcWwqDkwE+GRUjHQZ82u1T7SkwPPb8dCD8EzwoYm6h2Y2MlHkttmS05zTDdrzDiHWFtlHe
HGSX/e0A0moZJ88uqU1XT+FqPrtJv3Q37xwO537LrHC3zsAAE15huWce8ZFMCPROsDLi3LXpgeNz
sGu06htxmdFvLRWBtbXZ1gZ6I34TcaOY+1cCrEFQjm9QlZBATvruTl11RBRDB5zJ056XOSNAAoB1
FNwRKxhGsknJqpskJbwtvrpjFWvDa66LgYb7hLCrS0PpXm94QQqQK/POWQ62Rpqq+r0plyTkquX7
lS7TQin5Q/mKy2u7K13tEd8SaHiJqePBU705EMAB3rZbN63AajxPrQMx7iI2Iu5mGEuuJhTg83LH
ehaT16KN1ik0fD60+aXyP0ihYyKYF6e6lXATnb3P/SIS0NNECMQH3/xZN4CdkQsEVZ3Zxkev90Xx
iQ5Bpw22OJPPTfDvxoTv9s6VK/x+fJ72xxo6pr8v6BeqKcWVV8GzlSF4dgDCo73I6pZGWPZBewYw
4M0XJdtHQTSZDJqywRcmUBTAWW80bSMK+3Y8I827eJ5tXNKAp4Ib0CKbzqgl0ZMNyl3QR1FC+wbL
wDD7cJzuK8PCUBtIs0LEl6WZe9CzdQNiKrysnISZawSPcHukby1oKzlDQ4msFIAaZZDM2Zd6J3MM
D2F2X29XKNTU7odXpji14HBMGx5ndFTPTWBnQwpRbw6PMS15rSKGuAI1WNQ/Jg9hrxoF1EpTNsk/
YgeGPBW1SGs9ayrA5KEe3f2v7nZZ6JhT8GhTHzyuY7MaofiXMO3QSf+uEDEOJaY2gQ+dTyPx4cCZ
FjdUB2XQgJGS2ZXCWEj/MRWC1NngvdqeKnacEGSN9gdr0/64lV9rEGAb0vJEDpmmp2eYqjBnEzc/
aKDfdY/lkiT2MEJU6bJtnlz1Fbfd4zuctDU9Lr/rstcu4nMDq5/4XCLowtio9tU5MxBpQ/b2o29R
UAtEJa7vKAAvvGLeubq7IdgFr9R+LHo3glswYbwGZDbBuPn0+oaibYlL09pZoNWe7hQ6vj4lucB7
Mo/tlZwnlzFNuXKb2qDM3kedDe1khFKE7ojMEZQUtqHB2fY3ix67h4zuy9WpFjCS48OgQcxphOdW
hn1/L8Xi9LcazMn/94XAQT9MYzK5kNFevYxGxji+bpAuA5oYHiPREs2DMTTN48Bvob59prYSCxoM
MMSzQY49cyZ3ghWPzLgIJU/y2kDAjMCEkpBzbY7M6jKSoaU5tYw9465cRbPBH3LDOTJm3WAV+e9J
fZqyFLi50LNrRNJOtCEFJnuDN1itqGwLscHU/xWX4bxDYAL4GCtqN7fjMu39XK9GLTjiYpZd/1MI
nxRQCfQC0vA11lUcyj/rmAxdQGSlTI3wvvc3gwiz0Hnu/KRJRXsY5t/tQs7wA6Zg8tySj44TASp/
LgbAw8W0Mv6wHANEYGrNDTuJ0kbISUR6aFbEqR4ReD5+TrJYQIkcG278TZZS0R7Jf1SBj8mWbeS/
zm2RRGtTYruRuq6Uq9oUD4QLrASumV0oo7LgpckylSla+56PYwpdTpMveeM6a4bQckl9RvroatfO
HzOf1X+aUR05ukPwPeOAzDwkJ1kc8jhzbbLaqZm70EXXn+iP3CRT49JB0mXotCzsufqKnSCzUR7T
iEOIGAzvl3y/ZNHkQ/tnEtVsvCS9XABi4S2XCN1Ba+xAcS+ezDAVAlNx+a745gCocu2YhYwA3sYI
3Sz3rfE6rwHknGYTntMUfF73DbpDWms6Z5kgRg8IVGvloCY/2kbQuGp1ZuIDPM0laPczSGLLF8N3
6IOClfCrR3Sf6heD0GcJKzk3O7l1BZxfpb9ejExMAXu0t929YgKocuVsfuaAlocwGz7gQnLpuzxk
ZZSF5F7uYfI+7cCrnB5WoZj2N4pVIOACK2qr2SIy5tqU/d8RtMRrJwDuVshTC6CIu6rO7gZ4TLgd
ecdph0gOjJigJvAqI0SgNE9t/j4WDHzB+ueKEsfrlaNRO/K+UxGi80ev2QClLN4ajkjEN7lbW9o3
66g1MhxO0BzTtSoN8ELV/CdanSOJ1FAeBdxxhcq2TQ5O2o8HgKzXBdw/KlgG5vPlXt3JRQx4btE3
3PMLgmJxbMQcFgLWj6VDeTJw1by/AjhVxTKfvTDACRVtyCxCuiK/bKuLy8O0e1575hR/yVDIRNk8
kj83lYTNUqGMdrYb73vwZH5vLsF/xtOyTspWNhreGoaYFMx9r+9mTDz5yoiI+J5dRqYTvEzLHiH7
OZXg66pCEHPIUFfmUComPaoHWzVijW/kpvXdtl3GoiX+Q5CJjnDk/KgAo0O3F8FtGTHdmyxQVzmR
7ggJfLraQiwtlKIMd+c+Dd5SYRqK0RplwIfnBlowkKP30gKte7guemd1PYFkLHG+XVs8ucYYzSlE
mKPzOoo6lp29CBGyY/Qwyz3FjTV8DXcZPduR9yk5ztnaiGFOSiIYOjB4Acsj8mFF1ZXqF+sDsNUF
f2SanQIUCMymchFp0eUJyGxIouBHbIjEGgsj97FG+gDkqk1o01yIwuHwX+0G1fUEzcWSP7gi26ja
rhJlKQQYn7vMEhhkJbndr/jpiuZ2hhmWTedpcV1zhBLuL9m6UDigVEqYQfZumLCf9sc+iJyobJkw
s8Dx/kBE8d5mMG/9s2gkkqo1CDnOX1VO1iM6WSaMC/zuCw/Cp9/wUnsO/ETqAPw0/ObjoN1nPxUB
2A1BNo6jakh8G1cBh/fFCr8JAh+/98550FlOVF/KWHhFkVCqZAcIG6JOAzcySJQgUDCZF6dNt3WX
XhlACL8Z0qrBjDcpYD08r/c5Yml8p4sDqOSlMWN3bqG3blcGTcCh1d+XaKVvbjR6/slF+N1QXRJ7
NceEUUnoPfi7lRD61pVezfsx581mL6HXfSIIix0R+hKynGnGoL2sVAvZuRv5x70eoNTAbd1bDWwp
eHSy3ITNY7i+lgD8KcFVTgRpHoBHqVqTn1CdszdWopfN/mtsBF+9jvt/+vrlJVIuYksRvlQLhhNS
x6ik1g2t127IAyk+pT4lujcoK4KTBG2VImgQ/FWQpM4GRVr5ut8hGJ55ns2kOUTpTwei4mr+CnBi
wEfewjYs9dtuCD6j1HdQHXUa1BpCxfOPiNFfdlh+CooPGIrNJNCdh9VdGXCK5VUvAaaOHyo0NPqZ
uumAotAJRLvOf2vNxIlKzh02NnQ+hxW91kLzutEido06yvOq8D7o86PjSuwa4DukiOqMLX1zitM/
rqt8+uiF7AQ07Q9Z4hk+EwWe0xcgD4QqjF1hemm6eM0lCin39X1XfYD5tI5jKjxCq2+YXOAIL+vw
KEpV6VIY1T5t5aF8nn9+vzAkmEG++n68WEkEiPrZ18OdLq5XHU4toLJKww3O8jIV52Svq1sAvzQ9
3OPXM7giVm3akRBDuSNjg7NPbwnw5xR/VCHo7A0lHaBSpPOb/cltr9dx18gOk4Uz3zHCIYhUArhp
izXn5hl73lLNynAzfcC7VQcttZfDNyF+PErLO2GgUsH/Jkr9QshhF6J5NeVjFka0UdJ5R0IL4NWj
jLwnGEKLPdnB7aWicTbRJ6C45tck18ZjnFzQ11D5HeVSflhO8/nVpfT/IKgp2QnIo9K0C/0K5A5T
zphXZebMXGyXOv/jZBtX5gq3BSHBC5P6lavDDY/C9S78w8eBuAfKGI6dq9U9+yRgrHg66rstOlBg
YEhv7aNkw8Qiv1WxbnkVmfnht8n7kVCCw84iFyr8uU9roh0AQLH1JPRcHdxa0j3NewqXXgiuB8gw
ZsfTZZaaksx+OA4wbb/29VOM8j23o6C3QBxnrSke4WKRbZHS//iHQ/8nYSG2iEarkAXDw2szEY6W
rQ524UUXzuNrtOh5lFl6iJp5weh9cxny0Ks8PweKNNrtaXMk8Spi5YELkR4z9zlF9xxpL5X3bg/E
EH0Wu9awkWVLMMJEm0blSzlb44JNLe9WzIHF86UzBj5cKkmDXxUOq1IoHSqGEPXUggACTaFvdAp7
RtUZUU78Vb9mCC6Zq3Ul5xLXKBPFcU5Xp11188qC6jdbRukQnUJKeo/W58m2+qHg72cXplj+DGn4
iqrURCmbOsDMg7rj/lwrLuJ5mbZLNphEctGtx5pHqj4Ab/Ttzb9f61IjMl6Da71lg4dg/Sw8rclZ
34r+yzKtyx5MvGF+rIFRx7g2fbbCbIf7Q9e5WiDqRqt+9Dtn7yQWIE45QaRZe3ig2icemcCwu6Mb
JCOgckZ79ReTUWGAc9RXNJjk0LcvQv5zC9xeJ3ye3IuayLZhuvmHZSFU9zYYvG8KLCcP8utYs/QC
H7G5cLak2nRCrxUTUoA+jMFB8MMJOFYpWJ/leJUBV6b5bLhF+skEIrMqgVf46BQWeThRghe1mE1w
pgQWD8uZtc1cLurfW1WiZBdj3gpYgQYDwtAiuLKFVEETWSKc/fh3l3lWDdwAtIRB/KHq46jE8IfR
X7e3qgM63OqKSJc08A3YsFNg9YcJyK7xPAXTHyi48s12KQ5GgazddF/Tqv/t+4MCwL3Qbs1yeY75
fUwx9s+K5HFvQMqkxkCf7gSMwdvZXyoW06aFU9XTRankEi9FCZFe9k2aj9Y5Xu85ZKngifbEQIhT
mTy3Z5ab4FKF+nf2UVem25M4vVnBn0xxUPURo8bDQqcX2rEBT5Cd1S8oQRZdqwCYlFJkSn2lx6Nn
aco++oS1qtTjq50SvZBWgGAWcDuzD6z9eR/Cb2nXDvLkdeg3zKcFVI4RMJUpSzW8v2yTO5kDZO7q
dT9i3ZK5a8tZDfSzzsP4nBxA2EJMOmkePj/g/oPpvX6iF1gc7t/JnAU+08zhwTgw3V/xpzsOEAJW
IOQPdzh6VSHPql0fSkZdRdfP5bON0m6bZlO7k9SGmgCixRsEep8pHxrhJBIVHRaf2tM3q1ylwCjb
5+Yg8qvuxzC7JzhVUtZUWlIivxH/y2/tzxW869DUz1LO6E2VDpUAjgLFcIcziF1ag9V8iMRw96T+
aJjFRbnVmx9R/wA9JuPnxmyuKqdhPBegL+D9eQo4mJuS5Ilm/izRRxKewtNBLskcyeY28ai2sBJB
lEidHvEj796TdYvi1Tg3TYRp/UUoHllU6XcX7AY9UcaCyA2gs+izQfMQM9PSBWS1KC2jFPZl+iD5
MB+Jm3v4KWH3D8d+o87U8onsESN9wV/0UlBB8amlX3ScDq1r93CrXNBuEjLCd6p7Z+ncjVKEs0Bj
P3gzL4RNI9kyCQ5mUIgX0D5uGA9eOBgp3Qebtk4DMOvwOvn4EgVBqcItid32nwVp7HUFQNkxIa4q
s3+fhixzsvEQjtxGHpVTb/ijukTdlY6+3fwFrub37/zq/0m5VOs5YPZjmIdKZ+9jchuQ7AEtZ9qg
UclOwJgIrCBNfFa2uypctnbzWwrrTvoM0BebwxSMlO6ZSFm3kgsHNfKG7yef3KwsdAVzAWkUzaNR
DSrwaeAMH35HUB5X97AVz+04/5B4bHYIy1iKpPrBbqbiqMz0GQeTkKBMRx+3u4N4L8VxJF84SvcH
/KrIs9H1PWDmhdVWalF5TOESfjBsy8AuyfA5EWfKM/uc2n1K3XDN6OyR9Ei4FyB5VjKd4z+8L06y
fJPrEnyctNDoVzGKwMKP1a1bfGszRig4joRq9qUT6JRZ1Bu5M8866NNgWKDXOTEgvg8pWQ7V3BBj
tVR+zpaQ4Dke7yoii3aIhs+hw3JKy8E7wUlJvNULW39B428sPqh32rayZLtFCVtKAn/k2wetTLZT
MzhECr5MkSA/GgCgGcAfvuLhNMWpZIkBrUtsEJnPEw9Drnvy9hsW64FRTJQOK0rSEGS/6OITfeYC
PAss2Ov5CAgU5wZu/2U1N/0HPbt7NksNEnpplPdDRmDHR7d9gYu1xT0yW+MAcOz0iVQp04w8BCYR
GDDtrS7K5bPpHaCsmJPmgPtZLI5h0Rna0bs9yD03Ed0mxM6/1QlV8iC8nDFeP2zYULZDmPCHRdau
+F0P/FotHSeiYa+Q6rsISF+B9mdkcIIPoxxHdDqbd1yjoLfQ6LvfFtT+W7V5DpMS6gdFLpSpu6dE
QVmagL5S1tKy0QRkdtf/LiUkV4/tapHUR1f3d7gv9Uwg3PKQ1sVHKt5kw6j0XV5LY/dPomO3kQmw
5j1mlbJbInPnxq/CrgIwXlyUXJyAduCTavZcOsBPmXArgPJBtLcNKXTcGLuxnFT0adanBt/+nXdT
Fzbq8xZ+wgWdzrw4S5v2ApwExcd64YcTRvU5qV6ysgoTBqg+rG7/KlQQcLXCJtTIejf6CQryhdfj
We+ybJs0dzdwvLWXXn/XcNfnFpIw+H4cYdm2qSUQT4upOd520DY8Kcl7NBWHPKAGzdI0srg+uvmg
enThAbOeJQo49xAuApHu1eUeiXqBJaXYX5GIgzK/7lNJYtWpaepUlutUNbliWhH7rrXR0CJlZDE7
be5vStGzv9V/bWw5svoY7FSZ3DfSIS8jiGzQFsY2hXOQDfs7YuICbq95E6YvvcnPxvTibxTrB2FJ
ge9i3XJCVJMph7bZxZwidcserwxQhC0G74eEc5+k8TwLVipy5BUy64Nxv72QFdvWSaNATfzfXrb/
+1a1KUX8wiKpssl94PTagmZlukfUoEy/RPTi1uSNVoBh9gBCP/x9wGHfl/UFmdwpPaYSRR0ekq18
NylZaxNPlDTMxu0fiQZeCq+qSAeTLHj9Kzkb9Ov+WIwBme1pBHVpTyZ2VcoWRldm267PZgZz9+pD
MOegIHZMcEL6X6whLxIVkKOpI5vwSDKm+xytiR7eC+pWIeqVSD5puaTOnIf+NDRbq8OpI0pWQaSi
h6qmW/TUCP1PEjsYaMYwjWK3m+ZxD+hziybbrwQxkF6ToWsll3FLtMok//eKBGzT8hiaOZF21imK
XMrU7/jNgkDxvLeuqtrdjLYGOtAnx/Rqra18y4vXjrosaU4lXTwzehbXF+fsIBEKPgePlN9WlG1N
LKeEjSIwSEdJH9CFPUEFXVTqmMnczVgam65TCHrmCBVI4H9w5BKwPF/4OCYD25BwzxdWxhR+M5uH
OINPlIdc0xqxXgEjfiTRdVellyzRjwgHQkE3o6A0OHP9NfJo0bUE/ZLLG4mCCQTC359ckHWuEsJr
dG4CKoPJgg2t76WXeB8aco3XWUgJ24O+E9AvZsac6v1eKvTRDbdxikkHtQ+sEkQIiWTAvdCd2K1b
4+5GdGwSaenjXCM2JO3XI6Ow2wFcIN9dhxlTlMuqNhkcrNPFP2lmL0KO6YaLuA3pLIIByAvyw9P6
7VEXZ3NylZUBvunDRQeDaZYF1BTC0xjVtKGBf/L5wqw6qM6LDIq1YkLXaXLI9cyyeKY+pc1tLlP3
qlrUT58Uhhmy8Lps2jm/vGA+TZyyG+qDalbZqGVl/GKpoaBYSMnsmQEpR9XfsJ/LzIg8ZlLuqEDo
9FEi+A7lt2k5vpkLTWxtXtm69kIHd+L+XsETrWv5PR5BYF8bds3D/jbcug00TWfS+207dKqlqxaG
1YF8DES04RUZNkzsqrxOgtthzo/qKY+2fyc0awaFrKfc/B8MCusI07bawBkkAevWBH8yHzPjdEC3
5M72EmNnQHWWipsqlHdyAeRKiNNUzKuQ3ecrRXs+2G5wi8qs3nPQvlnXY2mHDFYs2iTINvh7j3OJ
VJueJu/88hjWbD1YC/bnK9BhbRTpuR+B1uGXyKaO7u/W1AUAXlq2toWXWnVQFvn1dfc6OiROVHXU
n81oIDJYAqNh654x+pxLZl5yFPtcnCUC9njxItupGXwPHs6cwa0+NHInsHMdYTMbK5oSIYXqc2LQ
wFjSAwabK1IcipOJ5wkozaRhF8fs8KjkBKLLaei+LiDKSBdnu2NfNW3WuqQrI+9+IqKbj/MqQn/o
SSX13y7Zf/7TszRJ8iHst5VBmuYG2mWeiGMQiBEHCDOT/SabURATDPUtPoxFI19gsGOKqKUKXMp6
TaCpgAOjtH1oDRU6P9/yTo2uAeGs8D/yLAYb+cReCcDeVE8LNwOm5aNTeYlY/kiy1T6Yl2617Ozr
ToJ+dw2PUiR2HgOONhAJF5e7wpsq+i/llIew1zIOKl4ND38CW9mzM0X0/wrnMXanTDIwA1vb9Qie
xH2S5WqhvXnhYshhf6VwMl9V6BOcwuUrZ5ywgaJx7SNlS0+MA0+j2g2xJoTxtlcYeBAKjrpI/bFY
8fRQJlB6l6XWLGywQA1RS6J4o/s5JoCH/gmv7jyOnfMPuiESk3j0hMOcYIMtGl9M0hNDwcRdEyGW
Rb6OMiebKew7hSJwjPfvXnSJvy9J/vu7kD3aN4iO62cjdi5kNJEqlaBDn5pNwbo36ULacKEPMRaw
Y6NMuKQesZ/4aPbNknXHsWZDdBhwGTghhefoOG5ZXVJ1ABSXuBZ9421ZYyzZE9HEByN1wyhhSxPC
lYFn2KVYTH5ihiepdGOeCocVRBmCYow3EkiX0iJS3Q472heGPwX4K+D5nuNt6tQgdrw4NgP0beFo
Qc6uCrpjXf40EKPwiZxeYMPTF0/V+nuv+Hey062oZ7iJ+0Q60COLV3Khhi+Iw+7Z3iTuXTf4Pt2z
wX3AmsEjOI73+Rq2hJEY84kXc9gkziDLsJ5sUOwtHa6hbOhkRihbD6csR++nwIx5t0To7lPbqubZ
fiA7FFpu5ABOBGohY0rieh59szGc9RNd4iQa/eM02eSbL2zoPd89Z57yTh0XLjWmpCgwfShCT9KQ
was+g/Lsxe++B0qtBCaTqZanGa+2kFOF6xR72mVivAsy1KfiQ0DfTzcAMFKFG53Qtb4zCuI1M6m2
mjPpKpprhPQyHusYE7W72tQXXJazVNOMKrnGPNntErT6MXkXQO59GfGdTWD9tjnskO9RX+0MYBXm
hP7Ss6olzzbNoSwiaLacKmm9DVkZQMfVU4dSrPk86NQdUB/zV81I3US3uK8RcEgekluLGnSSjhIq
LhhpCS3uOQoeIZV/L8iV/tAuiW/ey1WHfjheCa+U/is4J/qrTOX57y6b+a8onoR3OjMtTFj6tPzD
cUZOJ8G1525HRvNUQPJ/rJllr7xB39kZ5Kg4QXBruF0o3cGk7T7N5QaEVe6bSecWeSvuiv/PnAmw
OFCQGsXEwjmoUAZJpxlXdspLo131NqVaBMblxBIhzmnV3SN/3CJ54hf8inh6cv9ifFc6WkYqJS5L
dFmoqcoZ8NvgxWYl/2w72WEO9j5CMuwrWZIuTScJ/fTNEXOQUNJeYsFvVRfMZTv2t0zo5ltRVEWK
mCjoxeJqOvWAV1oqU5SYIoLgGVMpREJreHK4DJdQBrE/iTco9GuGBS1RMH4o6ghVf8izx2UTOjKi
9lz93fGeMarSjA5nf9zNQ74bKoTxbikpVc4Ehie2+Ol7TcvxhVj8krFA0OeN8A7hkIsimibbKllh
2io492fVf6JPEUw5vn1huvXbmibJvbEbV8R9GYlSIBChtvLHfYynhqrfuwALxGPhzfQfmv/zVDwd
CPqXnZBe9CJ4J9Ym6Wg2Eaqhc0dxOMbyq74jJR01j+Z2nVBw4PLbmHTd9VdG5hiMrIYxNOEbwl/e
lgDqB1IgtTrZGiRbsOQoMwx5YPZ97LAFo/WtMY6gCdohRqgu46NSo/dl9UGzLLjWq47+Xvt0kx+a
9kVOrOByyG6sK/9Vrilp/Hs+afAcLQ/nHtibvIjoMJt7ydvAvG373+tNos5diVbm5wN4Qr+L7lYE
O7JtEhcAZb4RRwm8K8hHIW3JJsYXZgnT6iyijJwoQ8H9ncQDIsdploAhSw4ewCmz8q61pNNsMK1H
CEnCPt8nvJrPQmBJiSCmuvs4Ei0/lidIPVIzhCA+JeL0wrx/YqAnmbdZP4JNxTHvbHMMSbGpDzoS
yIhVHqk/WLma/f233yCNSp9Ua4MTw7N8iZjm4ddbRljZf4ULDJ8Bhv8i2arAB/WNyT0ecANXBSnW
lWSEe9Y8v/g50xXqSKy5IGpzHB0CkKafaXHbeLOTNklgijP989wE4qpl8HwP7kqbxnR4+aLFxUSy
WREhCtmvY9LQ4OOX2R0h/VNWgSL8/quM6MC5V0ItbFBhIZ0WPb4XV4YGg+e8UdSSpwydBPEgqg9R
6JfWoWXc9xRdW3AggBD2RWoQwX6Pt2j/FHqSP8uB9DN/dz1CHTFndsYQmqjVfOYJ/27fKE5MOHAw
OtYYSQCKzHgBe+9jt68ki/T3Mr9Fpjv99pm0164oD5v0tAb8J44DUmRYhyyH9sSVQ2eM0nWswUFn
DrMOZC5hqXYBPVGtYJKjLu10WxzSmYMO+174WeOaaxp6CQLjKnswr5jdYMtYtF7jhpAJgRFbMsV+
z7iTOIdF5nOKMxcS4xFkMREwgk9XH4bWnFI2Nq/QqWdZnw9xxhc8IK0IgRYXpFAOwkMCNlnHCqko
dhth0MZeBIL/DU8UUDv99iH6UVKH5EtMdcGMa7NCdLk4jK0TCLQHBSeHnKQCytiIgvZfU5ik8hVV
sezHqPgD1GbEKya95xbu4aycg6+QuT7AvUZiimBzWSan12+Rwbn1MzZTHoymI8tVZbNQTIS5n8vE
oWlKyUwr5kzkw9pA+RrYqqky0rYv5Yls7lxVI0vD/prC6DhXZJxen/9iS7BVc895atbw9nHeQRyN
yCufxunBKq/v+Q0Sv0VcjW1Q3iaX6iKuIlw/0UK+XIjmCvIGK1DE03mRPnMkzUUqdRadAWS1DDv3
+B351NLi/1ecucAJPyWIokVtkF3EYjWEkR61PDxiHrNIVRR5mPY5Oa0ROtoMOsmENNOVs9pGw9/u
U4I5rJ5aNQriGTBe7dxc8rmH7QuRvPoL2YMD+SOEgKe9P+mk6W7xWAy/QnSkxYkHDGq97ivQJmMF
eqYSuZ9rTv1AwhWfzJqtGaAHrA2FO8F9GuGONov0C0tpTgKKTOb0Tx73Hw7F5VyaGQt70aLZs5Qd
u1JNvlyFb0eZPjrX1zpeeG37LcZEylDwuDTK3PkgqToSNwf6C+sCGa7xmMEJJrnhpA1iVEeQCGCv
FEGgXi3+IbdtvtWoMi4StAc2EcNCfkVExYixy7iSL8kxjgofahiGWAiLKXX7mUkTeU121HBTcbfD
tKP03ZTECGRuIcsmK8FMZRV0BD9Sdon+PV6FOJHlui2ID0uKskiLtalE/qHtx6+fSUyDg8Rn9O0J
I0Ox1cuB3GgIS5H5Jh/3HGVX5G1oKrIXdFcHYdiRWGeAn63KTI5KhagbzbW4x0i0NB0pko2K8yeX
Igl6PsCImWmL62aXhI0TcqNJAFVfborGoDRR5eAD/f0fnlplgTNCYdnU9m8aAlERSRpAcYct6TRv
EUwv5cuzu8at0GugS3LJ37Ip74V8UQqjlkCcSZ+JNdX5zOkm+D3eYixW5qDQSaG09WFHmnmb9rlJ
lKJIPZvGJ3JXpZoT0csWMsDapCyxNb4LakcriadxkbWSx0q7GAX5edeonSHKL4/vPQmefNsyrwD/
doanSaZ8RctsjVpCiUeOcMn7zxwlAZ1TXtgiGQy3KTF2Wnq7TdtUTptT8+4yeIAMdY8ao4w5KboG
55Z0PxVICnRJ0a6pGS+ajFSBFaD+oHDPH81ls3se91Vk02jiNA614wXZZN4Fs9svGtIFbY+7x6Z4
jET31w68zffXMqKZpNAa7v4BSpLWOwi/XkJ0zAFve6tuCPkLro2EWFO4b2vjB2B4jlY6PaDfyi+w
hL3kLJ/fmW76lpCmpD4L//T686NSg05b1+54DMXV55KMGhmz78p1xuA4vjggcrO1ww9FJNYb2pux
E6A1eyXj/KcPfqNYPPk62I0btOCji5IFvoxdkjWZPM9lLGN1Yh9iT1LsVRIDa9rtCP6Gd3TjK1hp
jQrEv364CltOqYdPDpGNdZgSr6TMXlXUp6MncBdrAW5T6PUmLlXX6NQa8AyX54o6VV8PIcS5rg03
jYgjRyiVSle1jxSyfjbdnL9Qx5roVsFplGKYI9X1r1lpLSdtg5o22A4JZ0nLLpmb7fDoMUS8YliF
Kg2kN9UessF/+mPhuxoTRYQW+ilxR30Cz8XYvOwHCFlvUEX2ywsUEN0Qng7ryZBOCLue/ukRD3wg
VkDhB8YqWSO6O7+elWFAf+GWW8IH6bOIYYnY0Zc68Mo8KOPgKZJPBppm0AQ4ukObuoBdKMo8E49X
eBsPfEuHhk4HCSF+zHendM3OM/XVr5n6pZ10IXfeGpgEaj/edP7DThU2j4MuLBUeBaGwFKFeoNsS
SSi2AzyHeEwtX0vIq3iXiz2KbKFdeQZU6AeZQ+NtcD5f+KXb7FSTgrgSOpeflLJTgt4waVzoMeZx
5IX0oaqXNkj4VT2kgFfvh4/1UUGc1N6z4lzNYOQ+n3aXlzZ89nELliJ1MG5omld8DvXjSs5DiqTf
WCLYJitFOntFTnPjNyUvGaJ5q+XRVpey7OJWwNIvFAocJlD3hUyR8pgSe9jp3decg4X0M7NXFnqc
/AD8iTZSziTzHhNBXoqiB+KguDIvPbbPARQmaCvHjxaOyf6lYrVt0IvDj3mzaHaVDazqfDbkx1fz
W8CrX405Hbh0v9dOBJUWCMzDL8AKMVgiBEZvdkl8CKKhIuwUh36K6nLXVp3QCC4N+JITsdBbFQOe
Me00+J5lIMTvi0cUb14Pwi9OiuWCZL8xSPw1nroeitaHuRT/edMneMagk/Us423xehUTRSRGccf+
GKMN9flQkxxMuAWQb2nh+vyFNKDEu/d05MUl0cN+NSBe88mFqspSqMpDM/vR9WdFkkt5oFgawRFF
RVJUmEkKgIe/vQ8GbOfQkY+D3plynLeapk3+D5SsOS4V0dsOzg9EyGaN4plZoJKnU7VkRqgyFDkz
eO40cpe57QR9Z0flBGi/FxbfvmEvqJxkxcokLnOt2Yd7BJ3AzGsteYzd08Yz4x/XfocC71CK8jMt
FSB/whcH/BNi6+JWJZSe5KJnf0OR6YWZaQEP6NiwvdIxLT9wTB07wlSw4J3DZSKvHXJI8CmzcJEC
povmNqNukduGv66CfuDvYqSnzGgKQ8D/Erh7W1e0ceSH9EMXLEEMKqggHPNpKNZgKbLUFYioFiLG
zEMHNMgWPMBJnQNIvonX7OaUKwip9qp/fZJE3x7s9VxUq1bGQle0ejb/Ye69k+QtkE3UoCtAP0pc
WviLbPksCTlMSoQ6zWKFl0lhsaqtvO+s6dHkSAFHpS+Q9aZ9RG8OJzF5OkXl0jf4W5bMY0iuvZzN
ldj1SWu3Dh9yQrCRzwW2CZM8AnLcZ8HBmzg4SL7Hq8osqDZGbQ6vrkmNpR317HkmaI99kvJ8bQv6
ySWbLKEs1ye1xwa6zPJJNjRnd6WpqwqGkGvJ1Xwqh8f1fqqY/DMGnZIUX5l7TI+CriXMraV7onBX
WTzGdO5cG5pGG6fONVVw7xMy89qkz5D3oROTK+C8zokL+ZuOnnTqZ/4U38AFXipQBk6GtDzZB9KC
BxZgKQfJfpHF9VqmNG4a57q3R2NJtyFvSfpLphiDKHXWnp+LU6t5VjmvVUR+jmtZwMMYfq6KGQ77
HfvH4TH2fa8ib32NyinqMDRBCUszWEscCvMOMaE/Dw7qEjSGbtuU7AIAJzgL2fQuy7r/hg6w4oHf
+0Oy9fsbbvvPioOr+3eZKD6hhmpegwV+1+l6+N9C1RXkTGwNtVFAUPGfxMe8cARjWyP2p3peby+F
JWvtM8ULk9+QKOA7Yu/eCRQxsWULa/Ll0csw3lwxx0n7A+SsHW4Hyo/gl0tlV/ycTL/m/xG0SnXM
+YefjeFgZazsFMH/3DaFm55AxmyFpTNjFPdDNvH3Ckp9zE36KtKnwkiKqiPhKFqn6y7QoimFaecG
kIxK2QejdwHfdr3mUKnoivbgqYzmRrfwWKjU192iOoApddttcangmz/c/UzuclmxEWviFvkanHw0
UZdMl6my6YyGzdbAeXWdIif97X3doD63EHL7C4d8jWXPMS1i9sqtx36Q3c3Lb+QQmHsDtnXhr0Tg
XgAEp+jSmgPu3vaRzXMZ/3cDWU/Lb4NiJVD6iWAeXHSuXAQs1O7w/8GwmeSSdMZbH3Gk+8bSSiTH
8v3Se8Zs/H8JIZIYJgoZSm5Q23YrBG9uwmLfdTtqOwmuT+Df+utzYKPcfLvBA4sicVIyzsgDUfL4
nYhwEAxieHjS0jA7W/5xMlcoLJMQ9MmY2tJX2E1FyvGbmLbRNivUnoTxF0GWvDcxJHEidJN10sTp
4IO5VYqGQdPDjTURuS6Um14PBZ5iPBWuHn+SUcG/2hjfzjnSzeT2xpyJ1X5SeAuNxdHuluqPa/of
EmWlDTxtf07EhAmz1mqrODpQ8FftPIS7a7LFUCP1Qe5lj1u/Oaem5berYdP8Xb2oGknb7P690Uei
dacFXYRJwZHDpCfoEBU1ELfNC39Wkv8fv14/RrPGA47fB2ci/F1jTTG71pNHTf5ArXbqCGAum/lZ
Fh0tYftFTmJ5O5vZj50eJF1biGhSHWzEQkkj2zXB5Qj5dENya41cZx4elA8wkph2njdhR09NSJsu
4C4GQHcZQrsguH0ZLpLiBWvWuonuEpMUqMxs0BnnaGynFsyq7HUkRDb9HOWNRE2XJYK9dXjihs10
hD7VF1T+5jaCjgB8pUWeVb7dCVxZR/m8g9hqe0/mfwOxpcT7D+5wHyXzPATGG/QmUlQUkRWmLCt1
uf19HKq1MHxd7NbxsWXohHV+QlNKHbtrBu4G4xEmdaz6sQUirnQxqMB9mvRddvdUVvjXvd2dyQDG
zowh4VUMBPUC7ArD3Dt0Lqm0eXyY0DlPYgUTbsXyFeH5lZCVEuZ1ZMZpKNrAtO97vifK0qIYN4WB
Wqn7VG2NG+kh6x73FEmGIt//j2+FNl6fHzjcubT3qLIT0VbWhXQKnCSjoJtyywl2H/7yO4uCEiLJ
yfMUTW9GAIwptyM716Q4TLUPGtQ6tCUiiqV39ziiFIcLTLIBK9p4sEi9DTAiirkK3AfW7xrIjsql
FFlbiIVncWob3ymDLh48/CMX7VtLxwNviiT+uHu+WIy+xg0rLIwJiO2jBbJ98Qw4uBhEHd0jicNf
2GvmLTH1CUd5l8UlxXCaEcdQaAsmTvPTYonC1kVCpusrfKrLWqLpQnDxQwtKOYELTGxPOzDb+ZX6
F52LiYrVi+Ny48Qo3T/MgDsaM33ozceLdYK/IrljIApE33S3DSFPkYyj3ZLVCYCYKJMDHWdFDy/e
qdIFHqD1crkdHcwNhQEePmlnZsgoE0xlNCwLCRbbgBQHnssgb5TMfMj9r96db0V4iDG8cZIsvpRb
apurORBwN6rWRpTT6P76sOYndsR+z7N5/mZ8AuhLcQORTXbg6TGGujjHzy2Dl5BgRDyaRgtr2Y9F
y9UiNhjg8M9K14tCzMEuXWwhkXS7dajZgYEQ6MCBLfD4AKJOFGs51r0Ae28+31Ev6ulDrA8Fairm
L3BJj7x8h+OzULGAvwMzMc+jJ1NrIxHvki/bB+ZObik+IIr2rPW1hnwyOjsjAUvNrVqIEICfQn5P
RZOw0VAuONYZZNdvGvLFaiRqVAvVEy/O88GXY6mKOa0nkkd1gb6bNsCkxCCLEAxcZYng+FM3yrFd
dT/BMBkokyuYh6WwC5FEF9uGLmS/ORhXfLFUSKBwlsFGtnnsdo4nMsQks5UW7GMz9WGzkHAnAum1
Xk43UxHMAgWxP5KSSeS329PjbzwVYHuXuoItTWCzsAdkbd7YcoOv4eAJDlv4cg7k06kTPwEw/Z2G
1WcnRUulKkPb3+dsXDEbX5Z5DsZwRYY8+ky9NxuVhSVeDUCeJskqMulqmeZf497ERJ0Xw74UOOG3
+ifD7l/hA9lkvEYX3wDWAnt9LYwWboYCt0W0opSGcrscctHSFapa4BzHqS2F7z5XPtUW0yPwlxUR
6bQO0eeYdYoYQRzu1t3JtRi18KCDEynHB00X6xgxMFiIlLOWnkHVlaxgCyVy8JoCp5ueDTt0Eoiz
sxlFB0cWGbvx9tGCqshL2mX9dNisGm36ICdrGtxNH484UVDk1yOSuw/WzlcpWD9HB+LjyqmuUFnF
vnz5NJBQ1z4h0weyh5wksz1lJisYXbomfpv5Nac7o30tByvUYbAw0tUl+fVjoeOffRNhSJ9UVvTy
x6MQIZ0NwYJxFLZko+OJ8c/v/s8hmhgo33/ffo8De0Dexx1OZebPbtuGwTiK91lgZaBPGR3WwX4w
tltVOyEmgK13z2iZU5ZskA0FVGyQ4kAYHISZYKPtKjx4krojTLYYD21cYPPbHq+y3vxgXEZIg3iw
WvSVeF/CyP4qr+krlscvA641+BPTHgFX79YURjR4z5SKKlDFaALDbAsuKnjfiUgaAq4F1w9EfHMC
ElcnIBv64d49SKRriOFJ3Ny7frx/A3Q5XuvCg2CRMcMIhv0oT79TM71CLvwcHFCQGKtkMu2IhkjZ
XnTl6wSE+20wmLtSHG2lVnHsVIMWcBNYNzrXNkkEEl4iTL54VhPSIOzn0ya586KICGKGIf7rJSIo
AURTvsmuVpvIWg3Rq9GZOg8vv9X4uUIciE8Rrt3+xjdFBeZVYhQrKpfPsii+H8Bb8fL3OBrHZdlg
RSXxO90w/ulxEGAWW0UyCG2P+TkVAByKno32dxwjr3+A35M/JHwx6E+NTVGze87/ackq1kRF7Mtz
5p9E3IXfOg1Kd8BHlGyAev+WJgup2tNEbF5HZEDF6bQ2fIt0VRaFfils69Zh7c32Hdxrlfna2OjX
n3UQnytnarOaR+ZiZMzIUkPIhaogS7QL49xoLCB4JPc3Lr8r3aEPkzGWO2Tkp4fCNG5KthtEcRBQ
Ji/KE8//fDf/W++n9M3zxShtykWUSOf3imKGcaunrAWIdOqObvL1l6oo2dUaiNwBurFOyLF8DYwT
Puy+khklSkA91DC0vZqgCZ8Fq1cZa1T7+Cc5YuK0fWCtF41rgUHk/F0LJdVcKi+o3mj+glm6OBbA
Q/djaWjvhA8M31x1j5CVCPAvOTpy6sMm55HD+pow82rLZEQx42L1238eXO/+vpKSAenq3A2l4Ccl
/r1kQEmPqBCk6j+GUsfL5eoQqvj+hEjq/7asYyFPcSenSiXXRc1Bw7MZt7eEAadF9LpOtafxtuPX
26s2LM8NedyEC3cqkT4KkPiD5O1nvlTWACWI7LVgJoQyCUAjSq1Kr4sv/ChgKOZhHrnV5dMi2Kiq
NKgOFSVsxO/2exVGhhhSQzO0omuBm7suDJhHqQRAfeODk0DIki3vuykgl3ENuGS1tlVWXl2Dq4g7
nlO2YZZ0FaLmmY22VWokQLgI64/aD4cKdHODawkBDPlGiFvZFOmTmidMx8WRebzJtZPIWMsaxNNx
LQuSuCb9fyYjxcSejPO0piqVBVNs1zVxsWwPcRSqch2ENiIAHo+rA8dBYDOKDEIzdb6y/TahSZjE
Ne0y+TMa88u4N138PrcETUZx0kfaiv/wDd3gJ3C9mCdaQr7n5Oqi/cvYw/hTQoQNwaNTP6d7hVXJ
M0/Lp1wUSJqs4CTpHpgOT2e+5kSPCtC8Co+TFrrvj51kzzs4Z/E3DBWY6WtDpWfhqGfBSg9W636W
a8GWYZxXL/Q6+pcPmEpvXhhs3fzAAmGCnYjrhKM1UErkDYtKM1kOxqkS0EdgUMIyPLE6VAme5A0Y
USyJ0JkTu/raBVoyq/OxUTQCC7qEoC2QeLlVOs+dnbXdpUxPb7AXYdNdUhCCBM1M5TsEAREwusDe
WyL2o4kZL7cm7t5pH6kKaHj3fnzjNuE7waMZDXFq8cu5biK5awFRl3YC2L1mWIQkoFVL/2VXAkz9
O6RYtl6fatekAoee7RlHP73vQxnc634KP+tH9XZ33rlJpSG1n2oVDZTap++NXPv7HlC5ZsdpHJuK
KJ2kYV5EYLlydSMvL7JWx/+j096BVCFf5Bo49Xh76TeQvTNm8BxFKXDfrK3+ryO3vo5OB/Cpp/Kp
RL2psQePWDVSlrZBxIs3UaR2kDEQfvLqH/nXYv2iq//k9svkeHoZdfQlRkbcnuefo5yGLrbBhoYo
Yd0wgTC3f9dexNzws+LP5hgLLrRtI/O2tgOLd3C4yCJmThJL52JoKM2j2dzZNvkhguzS3+iGNuM3
MbmfX9NQoHrXq0GytexFGn5dgG/j/qk66PxKHLUdpAtksa8/Y+octJF/YZpRUxpG1qOKKREg72ZF
go+QRbU40Q9mh7iX7715eJ89wzinONi4o6/7dU515m0iLQgv0zdXvE4+umwfSpat0oY0tIwSeEFM
uYFFm8JwlJPJJNwbzS2VNBB7RN62PwxNYzUEZz4ijPeAmwoVW3sR/tG+4n2xNC9AX/rIXYC2bRWQ
+9f395+psfcmOOiOps42jUbsiqgjTl8weY5ibNf9HtzbvAEx90lzNNLaU3YhqX0bJaXMtl8+2THC
sqZl0RKkGhyFo8nhr4n2Z6d3sDoT0JikImxZ56N4svHV1YSOkVTGXUTATvwVR7iTYZDgU8hWU+Pp
zGuI1/+EDZ1EzYbqoEh6dCKiYQzKv8R4symAsqlfAL4pq/xLpoXjxwCRCH7i+ZZjmqr/1OWl+2VP
pllki37dKQNIRYe6oNaibRXBg0wC54jVa3R8MGkqtU9uI4UW2JskORGNKDhIh+Sb77Xm3p93hprM
8/+crJK0gHxOVyGaL1Zf/PnmxrMPkDgCBQLxgyHNMz5pY5fPGqi2pCDgn2semXO+krEvyZMQG3e3
jAS++uKxr/CnpbvGR0gV6RpAr2jvamWI3DjLLR8jPj29zkIM1MPkjntsMAwW1NHxvrO+l4xywWvb
84ocgf9/UCNpLkEwCjNAwGtdB1lA+2+J4T65o4mHxOscpKwvko/yDe+RZosDBVsK0Wg4H0c4y02c
8yiXMrOlc9U/VS3Hwo8fuSUz95zt9ID34cfwCir+YF5L0rlnFPnlQl2UaPUFX7nwLn5iW4sD/fIr
LLsLutCztewqaiegcRagFkbio3fmUTNWHt/22NhNqFmJqlT41Lt7bkIP95Oi/bEc9U3e2OOhLBnm
bgXc4FGXsQFyrKubXrzBDv6vcri6wUdifsY67WlyE+pUyP4O0OGtF0rXn4c0MfGOO5YJK1MugMAP
DULYcrtFYmG2pp563AtmStMUUlVNI008yXkZq3+euTol+rxIAdZfPawFZicyqiRckO1gOnBA8UUS
G13/sZsBTv0gzejFJfU7LG9c7Y2ARWqGazvjd49s/eB7oTE0DpH2tbN1CKzoS03koHa9siOiBT/g
DmWKwuICnVMqZMEpda9FBAmmn2FamC+o5VAlpDcvtwRLDFYZY7x/n7UyzaHOVjuPXaUb9+Jqy1/d
bRBiAwN+HiNIhox447Z/5qs5cnDAbMm7tbtO2ZKqDLqkZK0iE1gG6SWc9/IqUebOtW1DUXNcH3nH
2UMV+UVc9XhgceQr9DiEFeISXxvgHDpx8wmEJ667hqFy8NqZdgg8veZlmJZbr6aWh9ulQ/ZrIdZr
Pdv6EByA1sNKW4vGedvBR+p51aYe3gjSxGWXhezZ8MeCJmlJqE0eWxHaVdxbIuoqEYST/G/TtM6i
OmtzLBIyNz2PgvcuB7cRB2Yljz6j4gMYDMB2kQcV8cOuUHX5jkZPkKxVntwmS1W/noiRzwQuxJn1
LcxGRNr0QlffPpFNCk2srhB5+03RLtvSQ2ctV9gOiRLD5OWm/fJw9rbg/D5+E8eV6B0TXUjq0RAd
pwxpFIeDLiLqTpxG9jqQdZ9YbI69dqJfsMb1soHaS9zyOG80yXbsEcpGzDXdDpzfutcuZsBcJGUs
7Lf5SzBGHNd5n9ISZqrtgIwBC8EFDOjm2Yb3l4zaaTo099xLT0uKrWydtsPtLbzgMvMJIR5YAwtU
VWLGj2It6Hk9ZLc82c2krpQ1hr5wW8xcpd9j/vWVu0zicoM61KyI4M03vTAyCIkJqTEmcZA62oA6
AmZsG6eQeWuTtkrCG43jOtEmAVfZARK7y1ZBTe5z+rBDY0Afd0ppu3pdWm7+HIkwXQnbhrbZvaDD
K7voWKVY8ramh3IUDvwPhLcTsdVaCwp/lKXF0aXnBIlm4cxkhQYa2lmNivAKEp67otnG5vILbqgm
e/UNhvHt/g6kisWROiqrrRBgUKts8okM8VM/4ggX+AvSQi3ivqeYinXjo9Br2/ZCqeQai1aBL54e
K5dY3RI1twoS+rDxkCreVPDL9N5RZxCdgIut7dv6lQi2Y1lUF0EGvKDhro+1uE1IXbZDNuo96Dvo
WLIVLk6e8NTrSfW1PnwIv4VAs1+LKXClzU39dt9B7gdKuUuYmyS3NS7M6NExynG+/jaPb649UZq9
vwbNj7fHT/lYFbXUbZHsRtXb0LYEefWHOH7bflk4MKoOfcVJy2nSO/FWElwFzGfgsCVwRQlJ9CXm
4Rcde8OVL4/xXw4KuujLkfRbPXkYl+fBRNSJCnp+YASS/81AQA61pCCO6S407cVZ7Z0RdmJLkLyS
NTM4E0gYgorhLEBzO8Jfntxp4+XouiY6FG++UvC9ArANxijlDvg7AP2VoLySvLGt5Lpfu5m4J1jv
TRjy7E4qwtU8V0KDtRn+9ioDXOBa27q3/F6KKbdxS9UDj44nxggoS98T5jFDTNRlZmPNaMca2VbI
8KGf0ky0DpSt8QZdFD9AelRLIfrbUu6H/r76aS/1e3W93DloYxsrMTjXCuLCrO/T/iq+oRMKNu1g
e83y/eDKhoi5mMoaJh4duj7yZa5zfBnxr++1JAwFtyAcORNvZj/COtAF9igSi68/NDXV+OI3MkXU
qpfYDWL/ufkA0qfEWadpjNuLoI1IB2QsgD1Q/K2/ofYVSlaUxMn2yJrBP59DU3fnV1XESflCKqym
BPZLvBw6sh/tv1z5n+PWLFiXCUtzialeMU9TmyxIBDblSbWiMpqWJwDmlgnd/CB57WMDsYzdvBlJ
Hdq8vmW7uIpunVJwfER3OGODTPtP8nV4TBIc8dEUf/F30JwYFDhoKlG+NKjCv2wpPUIflAuQVc1o
k3fxv1idRrTdCfiPXIVShfQ7L2RzEZWxU+t4mrCdqoYp4e94GP4KxKC36MzXL2SEfMRRNbLXoYLE
qLm+keuSfPWa/uxiCOVWzwUgzOcD/gX0rFOiErFhMLbwd5tAVUq5B1CKXXObCCV0utlFgp8ruQtg
9XL22iWU44Ja3Q8CO7uH2qSKAMERFbMB3hMdCKezx9h2IngTt7vW1IK6qyzq8NoMtC1R9GovTFfQ
rTHM99zi+RQTqyHIA2CHAqDo83Ph3+PMY5e9J1Y8tsqK8WApd9JMZTCdpv24EEUH67cxexdjo69c
PJfBw4cSn7pcKTfPwO1u1O4dS3oNNwC3fp3lzfWIds1I72E6Ohy6pTzBOnkybrMZH8AdLmjoUtcn
15i0nJPzRib/6+nCrXu1N9yJgqHEhOMWedwSI3afT7hr5d7/ZWA7Atu9B9XVw6vaXjOSuI4a9KZ2
UFJDR4pZW9NFd/ocrn40FDqyjZQ182EyzkKRWfaQz71vFZ3fnh83y9jzR5ozqnw9FSI8qUZ746WQ
uFdy/v560thvuGWBKD/Rfp2AZx/l1TxnNUvf2qjfeGyr3W579H8xf6X3sKtK7MRXFXnEkBunM50H
/Os2zbVBXhLKDUzwc3DRxaBnAjyzd3tM6Mkt8QzC7pGbT6R4IaW6VhaphVJ651fdrws0otWA5Y4W
DTYcw4qSJvykhQBkQrwnACUXr6tl2hTxyvLYM2K0B0OpwYd0XyHPHdvsMx3H3owtAQ8QJaVaLERh
xP4ZazO3ZP55T1kB1nD7ZiUNTVoooHYZaWM2nrz56wI2+qtypTXxdRAIC7Cjslrk5WQfOIgIeWgt
7o9VpQbe9odxQgXGmFul1WfFhTpr6oYxkvEB7gYP3AtamT7PtJvV/vDOhsWE1fvq8P0geJGkfI8U
aWBKjVoomxSM8BoTD4zGS03XnknaKC694cMTWsuRPd7VqD4jKvvMQc+/FgwPzMk36Z+NeYxtor6c
oUlfHJptO0fyN6HL7IhQcEugXT1a2Qu7ZJU0OiSAXl+3qb5NiRHi0cxf0GszB77pkm0ZUVY7wHI3
y6HLzXQiOSBcoSEvKYvDuzTeQqJRK26dVLwenayW7egS7mPW4yEob+87kh+eEnrHFf828lS6feIY
IPSmifPNhqSZMCKVqCh3AcHJ/AYcGWRjEz6vYC2+UM0rz5LSv0+NsdmryAcgQM+IFf0GG2Ip1UN9
9temHx+JBBYbzaorwBjp6PlBpEe27xG9RS5yqwAw6hEIUxK/lmKYnusF5ZYE0kWRhL2PO0lWMG6m
/EBbf2X+YfSYkF9TLZZdbyH15RNQE+JHf01wN5W8YXaV3WiVYcukpWSfzEodyNOp3qKmvUtKR8YX
IJd9sEQNrVRpBRt4p+9v3f3siTDWUZFR7gTR0avfJ/reC5QNNEmIegwtVDl3m7iS356CteTRC9RH
NiejUj/liMlu9VC+HdWSIyX5ffSVtRTVx6gHSj+DD8e13KKqyw8shoEaUAmQKR+hyzODzItJfIbl
9TB9rE0jNrvUlmo3Tpzyp2Y0izG+TYXLIuyhZDpXDJF8HwSqgCt85JdmiyJFmtWHxcTDpmlSwGvK
Lbo674TlybXEZe57rIiR4TMTjIixNPI4r8b2Y+wIYqUYEFVVnCunIfsoyYMZhTD64I9URYGAF7SM
3o4oby3d4IENNbdP0pnn+qruQ7JYuGxvCcjtdm2R7MZKHdTTUUPLYWQ7OBRwV+b3JzoyG7kwosfU
0ztqDI3jGW4VV4pZRtk3xIV3gvNmFIQaVi9zR325XKiTT9fiREGyFcDx4brnyq0sU40B6ZQ6LkIp
M8XheBmB9kfUoX3CC0P/f1ycfwfY6/iu5MK4j91JLGeM4RtDW6LRLqtmMbDcvT/XSrLJDfKkMTm9
mjsXdZdxU0I04VsXpjYme0rgAT1KfpNRdfw7ker/r1PQG8wQC3tQX6VN6YBk4vpcKg5Rt8Lm9NSb
7rzSpxDNurzL+13VWAPY4WX2leSQIsNtXJbsdC8stTWn7M4MK8ueeJtKrxOA3NaFZeXWgtY+Xdkw
rKqUzvnEFdhQ16NHIiSoLxGJ87ZACXK/wzhShQURun9AqzL1fuWhMpohwK5dA7IJYbAO66KNm6Bv
JREvhlWvBtMFtLf6kN2cG4jZh7503WR8rmrDnNqMJaJ0+VWmTXTtL22lKjr86ypHz8eKwxIqYojU
csKCewBWgOjt6BG5Ew/ppCn5Ct3Wb0vXCGKsn9CEgdyv90kaJMvIEZu+VeLO3u8vZN1ignXYkc0Q
M/TqeicqSRxE4pL4IODBUW5Ep71hhwotUaNqNxD07uZ+RRbcqfxku/g8UdvCgAoCK6wib/sX9B5Z
mQiZeRrTj5xDMC4H6QkQkqO7mc4of3bfYJfQHMywKEihFpKIhukAlPTiHV0bhFjlsxzmX3/pKSKC
SRQ+m0Fpv3IJCbba0PzExWmSdNVrSSTOcTwR3uHfNjGiK7ZYxOz41BK5jjX2dIlxG7vKLP2rWNr6
FH/EtN7LYbC8bgbPFLJvZU0hakVJmLUURJ+t3wkuTUCUJP5fHfgrjAexukZ+oxMUs8N1iGitprlE
pVkQvqnmy57KG/s9/1yTDhAMrsd5xehXaPgYeOcjxkNL8RYw9JfF6k0BEc0oYnb0FFkXOIImDhnN
v2i+s+ujVO5eJHQQ/tfCvd1QRelnacFoKCniROynmyWsuhEFmYNilKeq6j+Z81B3tLTHShAOanrJ
RUsbJOlMq5QZ5ElY/8aPrZ3K68maYoKVlByGPvh+uKvd/HwEoN80KvkYsZPlMmvCtfU8acWgQnNq
fr6AgJCoi1YVjnL659Z75KviinwaCl7Ps180Q+MJp82SkGGtWOfE61s5jgfOkHoiHajJ0XLOwPq/
djesYG+asRNkV29/EU/A3l8WmG17xFuzkcjd8Ic/u/Jh16E5dbUokihn0NomK7N5/jXmgKvJ0IJ1
GuQtrm+dR7Uz9gic6dA94ZlHEa2g2JiyXQBaeDidQ3xKwyCh+b3swGqNH08IUhKNgF4FuAm8+3lB
3P9kztiMkg9fLVlsq4P5QEhKxIBTNtGwOpcrMtYfz/2Ts02uTKOQfw36i9TsIvLQKVYMv1Js8EtC
UQilNTx+HRyW1b7WniYnEqnPO2kUxburJ4V1G9azBD8e3FgZyZehbohyKpQFFLvjdE1eCuRge5FX
pXBjEGGKOa3idaMQtaSPtTzAO0oRu+igy5ZE9w3CaJoCzcthjh4+sUmOJ1XgI6LnvvcfIdZgUOrP
17QgKNNEXa4astyOQ1VYxvCIbp5S0pPDQ8zFJL/ZFsRoTNHXtriWIchNuzRtHOR0LBETwg8teCqn
z7sGYMZxsmSG65ZPi/xF+ml9l58IBilTwlSaeUbdz+23Sqp83v0vS4T3I/xVVSseD6w08018WMRp
XeVwTrdpHkRasctJL2qBTHaAYTqA4icRzeTcexOt36B6JViymqaJVfX24rdgo/jshxEDVjCZNT3Z
+lClR32DYWqwFkUs3RXpjt14aPkybRqx/YXIDZk97vGp/gcKMvGuCDFi/Py7y4qY9Kgstqqd3eVu
I1u+b81JOqVpGeD+Sy/cqLJkl6ooGaMQAI11TFbzB/WREMxta2+pD1RO/B2hqNe0LwLYooH1JDVc
zcg7ci7abBMDBn1byBDt8xScwQcd8ETKz+MlukuBVdN3QIthPc2R4+gQ+72xhYyJGjpPz2EpUJ+Q
93DMdJPfHoz016h46OJAbX4IxqyIIGT3VV4czQNOrihaddjSb6mtPqgph2V6+PU/Wf6ucb+Flbqo
932yCnYlYwJk1RCXC62mjK7gaN/6rtZj+zCMnIcvAo7cAcFK4E7XTFA0YzKyUbOcqAaeTGs+FmgU
vjMbbCSmo5It9HN6h9wGONa8TZgcYKTuWVogMQQmNpMxZ23W7o7JU9ykfPZsPW3k6gB2DX9UihqG
FrTyXGGD+GYbLa/Wc5aTbCfSNIVSiNJzLzQPpPwGgJLAQ0Qn7RB6uJlplU/qbR3RcMFYTo1byYya
Mi9b+7BOqOPSsPRQM62LPFLdzov5TgMkrxe0DmZ3LplNLxXQaK/Fr/BU11NI9nmxHWIJY8pmSpXJ
VA6z5aGn3Up+2IdDt7nVjMerndP4tLDWdLpx0ci2T/0Z24KnIXpkicZRAOGYiZww3FmY163WOxMM
aqKCgbAcOgNfBnO391mRhRBfIVyy6CHKg9W2cpjw5mRtc6YQYvrmH64Iez+ygLkUJXUYAIm7Pbgv
kz6PaejhnEMrfOt26nGkcuMewXdvCqtbkepTU6oTEC/PwFe0l/hy9FQovrkCtNZSJ+4FHLmma37U
jj9A/0mCpsYzX7/1za9eD7E+0p1sm5s1tPZj0koC4dHQ1/y+51C1z5DUTfMxZ8vmK+LKI2Yts/tk
ZhX1in1B7j/SwU2aDz8HrBCSYd0JMuYiukQF7kEqJkUjecusGrJeEQkQi07OKY96Y88mf7fAmISJ
nokqrmxxP+Zc+3TkcgumHNii3cgMYpM2LnxgWinx0y8yFntxz7O/Kg8sEGSnsUkCkQZ+nTth8G3G
brMijn+owXaVvXt1atEh28Ll0weY5e/zEYwtRF/IwUB+d+w6IXEq1zlFOTiyzMQTIrI9bxDqG7W9
I8geohSIlWTdbDk23gwfwzszXrVCGxsSJwFKv/ezE+vgjs3SRz2gMqAK4ddbqA4uq8lOySjAH7D5
a+JADmTJ+njIyWKKRAR7sh5o2nf1LZaGMRk+J0u99VUkSnVcfzA/7QmvpjXxrUeau9K+LFtAqCPe
MzQ3CYldTwWPxV14jsIo1o23JxuUP1XGkeAgFQqOR9wDJwimhC5siSEXCLD/7SDaePaVYPj6Od6K
emDbKRyap4E8Q784VUpqZXszNE6AZCALAMxXcaDITlBAGg70AizLDGRAGnjy2wDg6wnTbnYmBGH5
i+t/vF20BL/OfTtd3Fe6cFGR/unavO92BGXRO7LPyGGle9GYyQTIvFzUKwx9zyB96JJPOYBT3udS
EhAlJUtxU6U1npeqVp9LKlfueUJ6a3mrlfKI4XulHxlkBQ0jw0jW05nFykTAiIClXpLnYOZTBPPs
cG2DROWZM1JCKk+iYG9911dQeumswCh6BLbcvHgt7UMt++napEI4RGuguMMsqyw09Ez8hnFEtW3V
piSKiiWjwWVwI0O8qS2lkCupdtCl3lgafrTQN+nSyTlGpjSyJSGD1hTKA3bOxXUsh+NnMreH2zzz
+ArDpgffN0Nq2ubVzuYCWxu8fH6EAAeuQNmpfSwWz2hHclyfBrE2f1FrRUjAxjH3tlRdnEnGS2Tn
n/PdYV2jZMxufICl4JnQk9sLTSZPV6pGbgtzzv7nMSbkc5kuWZ/78UZW3tC13IGkD5MoRe1nSxaJ
3lWbjMpVTob/5cxj1bQot8HVcNoZXnuuMCARUqEqkc8YgDx8RAq19FbiprmzNIHFmGQlfXTo4ejT
ZU55jhCUbpJKPogFBtk/KGU7UDvqCz3umPcz65vt0ryukKft1HAf4D3CV+7oysjj8G6o047etGsI
fhPeAWCMj6A0yt3BRhMv+Rzqc0tXFm813HQ8QasA3aNo8PofiF9MwgvywNPsuNOIkJfYWNyd3F4C
R1Dpw2lqq6oOIE/ZP6AFW7MUNXI3KG8mYVp96ZpFSExcJRwioWFSlkY3Gu8ngT9CL/C4KVUVlYyY
wztPikVCs2KQ60vvW5eivohMK9wiiMBTI/xOR9/ZguuLNd08enDpEV3bs9XEK5h2N0faJZsmtE1+
jwwOSCsFYhUlPYRDD17RJdT3qQQ0hvfR31IuLE2jH+pREdhycgXcx+gOXXt+61xTKj6oUTUVtjgy
10NqrFfdcVZypJzP4ljkQ7ye0hwqXa7WcKdwSZiRIw6oLkMrX5XXPGc05dTQ/8OGoWLfikLJFZl0
UfHVSX6J3VVLUznQWGGCqqlyaBaFtp9QVOAW73JOBqLQ62d2A+AloHZBbBjdXdRBNPgD31uwj9Wa
SBkJ93V7EdfGyCrGJVfleCzju0njgOQgpHs3CYx/UzXoRAre35OPBPfHGi4eFgVCtm2wklIC6WQb
lnHVOMgEb+2p4RZecl53HeVqMRIwfk0PVtHzw1xOXpM+vZdTU/QLL66KohhEH4pTrQ3Ch3kxexYB
lYI2K8H1bMNeI2fNYikLXiGOqqPKH9V4p8OPWHyG4fYJSMXLc78cT7gMLZ3dQgV8ZY5XcBvlUS8/
Ep0idJRIPxmIsxfFwTcy5fXb/UMV/sTKtKww8JxScchkOFGYmDwyNvb/K0476swOI+JbFMLsa8TR
1oAbragUic2mMxNbE/Mm8KoYioRwJDWayj44HScSj6lyg2U7ytbZHfl9wwoSGJwcurgub6JjkZYU
ZPtJdeB1xZ0IxJrUyWl40akoD5xiD539GrfvBHvgeHo+L9KG+imQMcH/xlVRVRWjhhZQZalRleHe
cLA2/uJr9904ue0PaRCA8bsV2TrMhTKX7hbm94u42XvVKMs5DnSwKT7yhNdooTcAwEQ0eA7EPFVh
HL5dCiGEnPDlOyT2BrogyXOpUETf2/e/2Cucyi+QuJGljj7xx37LPlyDr+isXLX+Lt63EkOp7Y7U
wtWNfyHvYO5L4yfPqSB1KQ2h/s+JpOkhUHKfz9n6ECOVwdAhpgZM5hSBdz0CBu3MABAo940cZ6C1
NUbVa1HEzXhjISPUd6xa6vIaZoqvPzCHALX2oQ/5dWqxkM9QuBzJLTL+h3FSCMQzAW1JoQG2/yE3
8dkPVey6PNePUjTvflWOgExzUeG/gvBN1uS4VRogqMT0skXIkKkkYqxQnLmMVpUnLhauGjovf+oc
bDOHEZlbDkeQwroKr0epNAoWhjmOxIxpknfuIyVBVIUDXmlBWcEYoX0g+oX/6CC0wr70E//DDH4X
7tM0cTD/n6d6tXpGGxmBqTsKW9AiYeoAsKI7RG7sUUO5MIj88C4tcrlTtx0xdOttTUCU57yqcv+m
l/8WVoM8jZeJTIZVm1Qy5suBagsrrJlsWAjCFhXt6Eo8jOs+jUGdCR6uukIKVcGzFtvnDHEKGOYp
LQYOuqUv2NW8vyoFFKGpv/CrCEuR6jJpgSmn4ZDbUvJXYAcpgW0y+trQlLob1wgU5h4NJFapv3AJ
a5DxOVJ746FZuCsIAnIjrdkINWeq1TSjiyf5CzuuSi6BSIKhsj/5fTgId3RTfFGqddQflLJ9k79H
jS5R6yqXLSxPbjd6HwnjEZmg5aubIYTQFNstNRFElmV5BzTveP9kzxumqcsyKlPDHST8pPGRIOIl
KZ+4So9YQ/0l/Ev/k/n19BE98xLmbcwEkiF7HGn9Uu7WfTG1wbpB/MhB/C3F8ttu4mxIv6xmvw4K
Q3V0LyOgW03R5kT2OErWEnXMGlElmH9bZ5REfKA4ndudLiW3prDmKRpRnHFz6eunXZZKeuStYlbs
YdxkMqeY0o5eXo8V9eU+qej/QOcbLyteB3OW3RaJQQXqqaAp8ntWTvcPS37yP8+f8nSCBqnrRezF
V34Si+v8rmzUtt53OwjFgpU0mixMffm4jU31VEfL12hmv7fdu27wojJiHURQ1F0NyihMWsIZbTUh
iZ/Eewe/tdYsbLFmVtcEHkBf8U6dIbG+WX2kdLj6XWft6icWyEoBcKdfPBmF8L1xsmy+UZTH/S97
GB5J1HAhZ0vLZWzTXDxmDLrfUOk2zKCjftM9eOCoFnDqY7dIKRK1f146lkCOa+WVOdUscNemIskL
/xo5bW1h4ZksE8sReCGePD/prendnGDRVcXXt7rmAyNZoQqGt5MvmUNeyH+4lFzKtSGVGH6gBmMp
IleAGh0id0xQxbAsweRD8iesf5z70WK9F1VGOjX0mPoWAxSAzTsNn4ghtdz25rnZGw90GqiJE18w
lsu2nprbNDwIpG6dgUXuphDSComQ5xea3jCTCT9/tIYe9fFfSBIgAL+dCr90RsdWQiF7ds2ERUEn
6d1ZNHIWyxD3yUXNCJA4kAHxFhAeI+DenVyfJbbhShkAsfXWANqj+G1sUBoDL4GnuClQ8PUC9U6d
0zsMHF5GuS4ED6b9d3GaL4qAD5/GRlp8HbMbDf44nqruL8/evMke80HbSO5s/uX00LlSbBo4x/H1
jILRXtXDv5S5FPwfs/4wjddsbeA2FQerKmesod74zclySuuUeCEGabCWR4UgpBhRkNy5NPKAVOtg
53WOOpkTJUhpZgsEOvCkVb42W/BpFqG/NbF2S1QZelQ/wv+rsiMDs1Ga/7NSRArLLHuaPSUshaGS
hDkL1Ib9X8yab0D/jF829ZhdioyT+eQQwrWiGeMWrmVe0vHDhQeyMTdkXQRXXwVOaJm+vpIEeCJ5
r8RWXv700LHI2X1PgyWR7YAR225hfyxkktQFN6EF5ZRba/9Msv/1v8ys1FXNKcmuH7jpS+jvp/6r
WF6anaJXwFAykoKPQ8ysxcGLCdB4pic8SimgnIr+3Yoqv0j/OA75J2Bbs/Azx/h4kuLBPRz6ARlM
ss1+o2+qMo+tghjocRgwseYVsPOM8QzW5JEDduby2nyn4fe2QQcme3NoKehGy6E0+i9PZFswt//E
XZUYs5z0xi50tTGmLcw5z+wE5+Kf5snIaLu06Pn3ljue2od1akDCbUtCQc4LN7kBjxmLt7eY2Qth
ylNm77WZzyssmujEQyrhIGfO8HQH6jq+Ogf7pjLUnChOWCsmYDErf1wnqM6btb41DGcavXOxAAJC
LHxLCaoOmIIi5ZSPcn+/++198m6kKnH8sibOnzMuCkNhktf1WUohIMaaWFv/BMPIcE3h9h8zjrpH
k+dSbNRMBVWReU2kFLEMQENywi94BcXgPU+ti9D5L9C3hv52C6VvhOCPNOyt+SQCrdLL0Rt63yV8
7bXXuakmFVn37N2XfU2yFyGcC2Mo9BkfUQOdVyU765voASroIZvAgrr3HNuue76aLhJAYjEsAkfC
nMkZIOK+3YIiSqrN7UCRfoChQ5T+6rYE3w5HPTAzLEv3J079KvO0yFz5UGjIF6yb+Ygr9A8JvKSP
P9Sof9/6CAwLnAqgUtU/ABgBy8TU6evplEDfTbJjaKkYQRHWLacJ0W2LGTKbS580m5nsonU4n3Xa
TnJaZs92SeKhLteCGC1JEhmvYx9KUJUotEABJkZXSqvqjEv7kdMyo73NVtyDo3iJrtigWB5jBdXE
6CHVdboIOCbFXsGd0iTmdcq45Rf3H+bL9cJcT0UteJBRHwVjURnaImri0uZfogScgshO9oLBs5YI
HO71A7jcI6W7Ch4QP2cu7JbRvN1iA4OwzQgy8X6ki/cqtlBRMhy4McSdXF4KSgBoQXcQ2T5bpSq3
EQVPLaMHH6+jca7GuvXgI1UzbZECbDyJ94bblpxT1dAYF1fBoaZYJ+vB6RaL2L6xyQ0jx0iNdxNq
X9OOKwvZaz5mORSdgjgbuGiptgINuc38QfeoYvFnROTm5mfLX2kegZLoQnlBHZA/pMauJFJIhkMP
IrShCkXrDGlsfAgogcQLe4BVb5XgeZYcN0wvUajKPV3F6xm62CUtrgnZA2pRuNbc0Bor7pGveLX4
8VoavW2OC+F19c4JyK4Nbi/lP+GYy2Jeu865iMnd0tAO8KozuFO1xN0VAZIgYriaPBQ/UsJBoL2B
gsv2IKA4KRWUYOfTngJaYyQCB8R9j1ubs6kVspdeKQFp4P4KPDcYdCvztf+k6zXZ+rqIEQxd7a/k
uR8mneuH6DBzflboL8o3qrFmw4W8LnrLTAqgJnKtLokjzRHCZKjw7kpYYaU4IIrlHUFX1JAQrc3Z
jhqRuwo4X37YXyyNJ5cKzr+8uyKheD0SE+/6reZV2iowuSTAhnOkozGArbGS9xSJE3Fjp476sFD3
Uxpv6AI13UZS8Iwtny/eQhncss7n0PWpfTx0Q6clQy9iB4NiMefswEgcYuaVyssXOfaAOx8/8PYr
cx+x7zs4ozTknnyzHJIAguCsMVbT1apsENFTAXngvdwRSRQwhvGAQw4YhsiKYqzRNPcIoH9GbLpq
2jw+7xffKOjy1XL9BaPyBvFqp42YtnBu1b+BGpqDa3188VRzPmQr5+4hMCU2YTGmM5nuf+jT/aMW
VMfmIhF1uNQ44KPh+EXbLwP1il8w+MYsFxGkUKT8EeUX9hGgFvPjBuI8Y0w7YitBzHfpLiMe00Gf
nvEi1tTdTJSAJJvzOzY52asDJn+JNeoYlZv60LvQ7WXbZlnQ2MX4DEOEXcRUOq7MzMRhsDIf1LRu
GpgvshRHFJYNEpylgULyXVdN6ErJdyDzG8y51HX3i+SzHbwYLR7bp6WK3xKlaKMiWkblfVJqethF
7Po58WChMfaPGarblbm8A+S5CcyttQA7zjTD6i8IPbInuN24xhRJLSAuWJbbrdcGZsScBLY1EIgs
mh+XsmqYqZQZ7S9q1ri2ZptSp67w7pHCwWjATSotROcCFH1fwL9N2Od0a6V0kT1HGi2J0qdpmuxB
l3wuzWBeWz/+93G46L3LTaUnor2bataJUKKA8F2wn2IpuAImWs8iHheJEbw5Gvgt8MsrK7KTeR9n
fizmhEPWOPJQqXgC27Yctpr8504sR0C8Z2uhXU5trNGBb1dIOrO7vNGvs3uinQffWLnkk9ODUAKG
/CYLHeWtcmXDDLhcfCPbgU+PMeettPU5+P87+lpiGcePip6rBYifEvh7lSe7TXLW+y0dypYZDH7m
cb8ywTwNVlP687ikWc8mPbgYfYxX/x1fI+o22UwQqqF5QF05bUMwEt3KoR+jyEEK8kMai22sYZmk
YEPNiwtTY6gW1ms2zpGkpYIAQp5sK3DCOojBZ9PlRSlXRsPqRu5XVtndfv6MpCz7+GGFmkc/Zu6K
ZkRVz1rsEeqzTiR5wEtzXZ74IUFu+oWfFmzwtBQZV+Hcdu6sG4nkXIQOlkr34mIt6pTHiqd1xULh
nKmW5OBUYhYLFBgxV2ilrHva/PD9q+c1J+HlHhcvcUcO15IY7HauEKo7K2bDqXV/Dxd8ZU/hjZ5S
hwczVKeL9P/NEmYLeLmJgS4Yiq0FQPrWEfihynEteAw2TAwuLDnhgzXpchz5brio58cE15drwbnd
2V+d+1AjWNO/j6XipeNRREWjOwNjdiBf2XWYPp6LywY3oVnM5M/IqtOpOJH+jGODBed6WoFG3GEE
zXdLj9sjbYAAEWNxCLeQExEvTKRIsXV7cvQc8Gg451HPAAScsElzEbEM/B6g4ZIQy9rQw2x8woRg
xbb7NzoqUQNprBSPMvdnhEUrQUdBdx9h9YQYAzBaUgE+DEz2xQ9fRx1BZxK9NwJaMG3jY8ooPxiM
o6CxfLoN2ri+u4XWPnrhZrjsCwAQiR6jW5tfenC2VKwK+604NBrutsnmkq4wPLq/9xlI40OwGo31
cM3AG6XtX1AGnmOK3chsIfoBMx33q6OZY5oVUtLdqYdxUBe0whZqRyBUUORZM4H3ua/t0IeXURri
kMQsnCr5BL+aZfcArcspjRPJ05mpUFivMfZw7WNS1UAZg5Yg+kEtPlUBpv6bNHP7R5KXwnnWvux5
bfPLG1qrN8ywfQfG41DS20F7j8cO8fnhxjBVY1dcjRFe60Je3rPnrA6er1QVY8x9mx7gBFuGZC/Z
NYfVDEx/xuRfc1wwDEzuETJIUGlHpFkt5GA+8VDl8E1etYb0Wft3fSFp7tapGJqwygIrH26ekV8R
Hx0inrj6gbZFkGJuDBSFIVgUXX2gXVd0fL2cjwM8abPj6q+NEXozT/AZXnchEa2jl2khzSYXVoz+
idHbPM5zKPpTqJMWfMnKpQxe4YSMgFci3bvealcmBJkwCqqONHFMt8IQ7U6Am+jWU3NhlJrundFc
lZMj+1MAT0q/ObWxEJBBi/V52Y0zFWONXJuxtpI8xZ0onJ+WGiZL5qfs/GwfK8RqNvPH29TzCEKr
HCHkrpzhzQyVva7PRqZYcZmWQKJ6+0PgaUADEj9U36E5NsPu9nP38fOCB7Kfj20rQ6ETudGIHvtL
viGOQ2b6fI7qabNe4Q4yRRNa683w1w0t3OJVNgnJ7GFDVZfTQGIKrHWVQLh8XVhAzLlk6RzYvt3z
9BahT86oBPXcHQvKK5L9TBZKEvoMYb4k1SOQ4Bk/q/tQvsdyrnfStb/4uM+a6jsdVizpF1/EDb2r
7CPnQosx5Val3GyiX3i285vVqrccy1/R3VUA8UmDWKkV/JJHxECDAD1wwRdpqm7kkCrl5vdXpqEo
Z9XychOK00YNpqHrG9UFH4jHSKZxZCVt8KRs+Qxl6OG3hnLpJK800pL9mnhTZ7phOPm9rz5O5jl6
BVyfuNXJIxT7fXycrpIsdmNsJpHen4u7d8Dk2dMqVVHtXtKTN8neuC9pOkoyUyMY1EmFmHGdzCAK
TQwAecF08ygsL/6m1zHGSozBrbJMbEgG0qRWuNJKI6Qx/DnhNhACkigjpuEmLkCGKn8mYIAOQ46Y
acaKbb50Z/L2mnSSV2MBispAZU+U0crp0JdHi5nZccMCLT7ruUTCMBaH+w0HbHzZnZqbylhvbHcN
aJdvJRMykGSWC8uG1mwdTzsMpLaV4zB0YoYlJMmPqaMGVNYpuNp9EQ9sDuw1ZZuezGCJcaTxLcUN
RSQHIkbd3YIH0WgK1wzcg8lXdZ7I/Wh0iWIXxeZYrq8DyGeuSdFPnEFe4ULmNej2czKUnHqaDx9K
VpYMCJSOXVHcPA1Vhvx22Ddyb2McYJ8JPkp5lciI/wt9R2xO4HRIs6KlJLhWMssOH7rymFndWQK3
aSmG0WoFgGKN7Wd8syxk3pWiiSH0msRFQGAaGzj6+LV0OTRJZCsscyu6x6kfMfTgaeKAfU6lA8rl
DN6t7dGuuS5nh6u2alCm35Nzg5JJACbF24Lw4pJEVDaphT3tIb6HmAhA9vtRPuggBjGXBTkQrMid
dVpC3nicAzEX4kQLVbKf0KNx59vPzrWfUogpOQrJvwSVE/7AUJRP1RPfJE8V+gkG5i62eS7KLZ6f
0ZnkLQyATXHGvnZ223zaerYbWoVPHsulbRXUEd8CUZ1ZDV/m6avlneQjhZDLmhOGkFTv643FKaR1
eOqSFDugJiyFyPeTAFJ9/4HYklaSGs0urwesoxGvFhyjno3I2Lzv7lzwfpXRkVHvwkMR1U57SYl4
sJjJlCRwSYFeTKbLPgtFbZZtx3B4wZX0yizO6Kx+oiaaUDhBQ1+SIJKp43pza+MgqNkZrBHrP23r
L1qxH3pD4dzp3NKkHDZpHbMDqnxi/PeSDhQBG5ODRvmPX6bzLiRFHaVUwhgQtmK69O+UIsGxtObG
diSFCSske/Ef/cFZE5cLhnnIHNdX/uQQoCohwsj+14OoH8qGHCyZw13YN0jAx2GecQGTU128KVP+
u4BKFwpji5ehdo7efZUjR5i7k8mNG6uvTuMUFrZr5+xk962+WyN+DtTT8sqkcxUi+ecg0g8jA455
kELrbr8uAs1fOYG91edQ9t2wTmkECvfMUEswtITAkT0EFrNTEmblVePm35Cc42rs6ryzd6bVcVqV
YOZjIgGz+OrY/ZyRdYYWMISAGuTWL8/H7JYbdLbvfiawHA9Uko/NGr+bdmvmMFG/6RA4ltYd+f2t
eIYmkAgvWIuuIgyWGlGTWndjt8MPcMbSmhkfBgyyhqm2QSnPxGtx35doUmnQ2fVonJLpgNcSBl1m
Ib4+X2Dg1zvEgAgBfRH+lJCKWvz8b1TCEOTn5G0vCJOl0ZV74wqzcex9RMiHzRdWGY4tbpUhWxio
q9XTs22fhNxe99aqWQOTtsRTbWFugl+zxuOfisyOdU72iAzAh5wXLl+51AarL3TFghKUBdaWZqU5
QJyjnPkiZ6QR8fcV/DPxifAsY5EcQS1apx/7nJUoDWVWtWV4atINf7fcfZvU3vco00BAGn0b+fq6
zd+3OEKB46/l1eOy6bkMn6FBjBFpn107rbLMw+P3DHeEIxM7W+hZtTlxWrmg7ZDsm7fPFP/mBXaj
sl9+wHk7Z9sd5U0zgQuvUCxDlb4wsERO/4y/HCOs61K7S+ss3rmm+TsaoBmNtPpEgA8LDTPwc7/3
DQA0O6EGdWy9oVbdTKP6V/VxTpUL0zy1WSvQB3Ko8O57x4XiS9rowUuawIQ1xvxo+8J2W8NpaAFy
n4K0nuDycFasPb7jXi8rFz7s7xu0ui17SrJdgwcTevwuYaMi4nXUvYY+eoruiraPNotoKbvErdeZ
adH1j+hTrdZFS6gqyn/CIVQEkqiLYXaSrYjcA7Ku9rGzEl7Xstb7MJa23r98EMOqTY57CeWpjOri
CawKsjTc/+/5970orcgELXyBKBC7g/SwiKgq2guUnvox22PWBb6D9wxVY0CGDFliErbTbIkXnDWO
zCUoGqaLWadBTLIUO2Bz0Ehes2rFE2fUt/lpuKZMd5VMECLaT5gaq/+a97OSwvycybqfcDX+B9RR
1SdZYduwXc8PQyqI87VRmRDFEbapFH4bKlNFJlEQ9WQh4YlDFlK2wGXCt9TVxJY8M/ucZGdBPFhl
A3GLHiILAMCqWvEFD7NdVZ5zWkrfMXvtyZb5um4VBoXS/NUjOTPbWaIIgWyhi9OH66GJRRsQMK91
GO+uXL4yCes0UGSUsCH9Jg5OOapTRVPqB8R5tjetAld9S9USWUJnE0VqwMqtwEYGLuQWCUYIVvAw
XlakUTLs2gAvns1oTzKaQ3HZqVBalVS4E2n5NWRbg1tx9HFkecT0gstjD9a0RQWrDYWvYsXD2cY/
Ptql1oNDRgbg6bKOsoKt5GLE15qOOsMGEw4bYbcFgwrtGRpeIBxaWH2zcK4yZljEGsPxHDqGv6om
0KCWMZp7Qc0CDAk1lYRkx4g/vG/SU4vKF91DOqkaQ2NYDBIVV2lCLe0zboSBHWV2oI1LLNDxJfXI
v6H1EpRAprjYRHSFwqZrCHleb9X6WJGD2xP8aEXKC8UNX/UpUBL3MmYTNQ4g54TnF0jHCorAOLWV
WG5uX/3Eyh//BiXHiFUlBAvOuznTEUrzOBrPxjg9WiY99HYpSx5kFBeC3mNfHcD78Vvri+fLPV70
gKOUU0cZXJq0c10A0SkH4Es0qiZYXkZ7wcj31sAmM+TViOgVo1TQ3jEmyvfHEmpV3iPQGw6PnHca
deqibW7GR+OdPXHS0RjjxOOxdmf2l2JUb8YRktM2cymvUoSYUorlZLK5r4uVMLVUij0xOXQRgXae
uszKUVQ9AD3ZRWYPVvFlvcib8+TOx+XQQ5bweijnlN+I3DxCGeid8Euv/NtGr32e/axNUaOuy3yO
H+Cl8T7cLQUmbTKX2J4GDoeFqFFajyUoINF8WaefGlkdG/6DxsNtVscBh829fW5SGj6+SUs5J3I+
TiZjsmKxQT3v9qKLpzzlTLXKeu5s8bBotXFwXyfa+YvRuqMIDRvY59QzIUGNG3u/2mAFMXJqtOpP
tHa6ge0yqbln0vNHEyXWdSXfCYbIleim+qddkiDgnuc71ZrXLy9ueNKT0tvBgezHQZtu073UU/dD
s7c4ooFlcoZiLo4c2W75W5AjxhANDvYmxtA3lcjgFhI+AdTmA+iJ/8R3xjbhRgOXRqbDh6Y6Ma/l
vgew68hktwONS0IbOfAd6hBLxKX/VLeIaimOU6IkWFX5roBveR5Tq6ZcU5slvjgRpL0ACVcdQx3H
Um5CzvYHz9UJCAMl2mnNfg45RJ/p4xLsfKNmdEXw6Fy7Z4j01JwYFYuDLn1uCZS1VVuU+7kGgFml
EkKjjse48YwPeEZOwxYvF6RgpFOziWmIS9iCpHdHhTfXB47PSSN8fHBwL0YiUaFhuJ3JZArGeb84
FdjN1H16JIMXC6Ca7ij7u7riKg7Fw6BG7nkariqzU778YTNjZHIFE2CRShLCrQBXUxSd3RNQdUsu
XY09qaTpTFYpkOt8lMjumuvIBUlwnpH10HGS0GVFWcb8QHSrSip4KXQaHK0po6lwcdMeJKvG0Cb7
5934M/cJDLt/tSsdoFe1mXtpIV0keBiXD8gxon84v9URgGhCQTYqlachTEWwBV8zrEQC+h4KakCl
8gT1n9fLMOzxaCkZSr7OChjp5CZkfgvORq/o7VEC+QIFxIHzbBPaUSbVUhpDALqF2OO8Rlg7U8w3
kgTKixT3Z2QQClwrWa+zbXRi5sFJBHw7rGuSTr5cdgpCRuQy1q3RxRZnSqSRP63lx2F1SePc3UGu
YfwTirsGcW8XaBTznNLQyriq4V4YeGBgJrthVNd1r0ce4WGOikgfUvZGmW9WarvzbGKpWI5vkY2b
xrc2DAHEk6ObRKOFX/mWXV5ghK5yBs/lXcfv3rvcOZt069lTVpGRRVZCP95siUeMaNhcxOviSls3
TbZeok6GiSY+TUBDq1yALGIACM6T6TUpcns7d/xx+IVYZZDwsDyuE9fc1R+9f9VtLh3Gkg6gnUyh
HKPMQzHWoucGfNHQau5b5g8xprRJTxPY1w8wW+cv3RDoF1KkOwSSkfZJgL0EY911cblFJCFFyttZ
QgVrSprXnb9IOcaNC028SVONlmUYHxDqoHXaGcrmhFJH8gIAKDDKJ9uYqL2mPWhYhTlHKd8bXxiQ
DkTKujM0O4gJwTwRpJIkC+Y5kDu+c58vcdiYVSzX/lOfu3vZW7EUw3sZOpUloeMQ0VbD09VWJjml
0dwndhm9eA8BHez3xscboxNY+cWAsMAkELWP1BYoWD6pPGAYs4HMlnniUWdIMo5/LNQL9ySQGmga
X+nmjRIWCsywPnbkXJy75+/54H+RFLN0TGoWkaCshwLRbIxU0MktbhkeHLO+DgIwra1bgBoD/hIX
aXSod1LFoBLBLLxx6xYOXmcmQsq6dhWgixG8dIaLQPTJ1S31zVAmeoc73pK7r1CVDllUgBKqtyC0
MlRH0jQiLyj8C2VPbdeoPxOjki+OGNlO0HX6orcLEwXs5H+X7wH2g6ek2J7EZsCGSoVAou0AIee7
0obx69B7AKpahyzvwq9mZsdXAhBwfjSi615iuPuls0F+kZ6Hxp5zfI802cGAMUEWiAlS6ehG+oNw
hnVpxa5E2nnsSHm0jEpL2JzmnSBQYfaO64A4jhQnqOsdTVfA89RRz+/XpkWBCWmMLjyPUnT9XXSq
F22GUTw46rHH1zsCpD3aCI4XBEILxTXBfFj4RSrA4zw9VjCRP98EtTAjUKPR1BdqXkwVvW7brP/G
wuAw1aWsHXwk+Ym0yFoo8oyZP6s3SOoLNtV46I/51/0G0v0oZOdkcGaks3Hzk2Ildq/j/UrrJYw3
nYsG9YFF1KKk+yrvlZGmV6pmdc0qDL6ZXkdzpfgyN0H7CWPJGPdLOm3wAliFzuLoag6CwnbnkcTg
8Ww0XdQ8Cprdma9wIHt5ceZbuZAYgUUkRRG2aLAD7ACHMM144RMHClYDZqhtgG7l1mjhftwi9z0z
5xs0XkmSEZr8dptcrGipOP8CighuFNLNUXpSuk5NPutKnFGb1bd/TD0Jzfn5R2Oq98FG9Ou5nJBv
bPGJaCbk4peMHcOlRIseU+8Iu8gdnZtVhCtaXYUwExTdyXlO9wInuWvFMY/BkZdTaHmuMNajzsDa
Wk9WdWMwKdVsKEXsf2WRB7nR2wJKG1NDdmS2WkZhRgjg+Epl7hTym+SJjDRYpqAQhjx3uVuDYg0v
JiFVAEPuwe3URLYJ2k4dGXY9SLMyss9ZrcaVnWbogTjLV23z9la5jrZ+7Z4sUOYu43F+saoqO93K
oCAiCOj6fm/iUmQh9lSw5e8lHq5ZoFBbuMC2YZ/TMjoXDmiw+24RqI2O3M5MZIz1RPGuqOPXG5GZ
PwXZwP0keWrlYLVy5orZPbDZSVPoCzNGcl/1lKTlpdPnwssHNP3PcIxMnFq/XkNBkT4aXk0jwlk1
X/5YDPMwMhZ0yUsggkzqCZ5AJ6usrKRWw7BBQwwQH4wHs23eltp4hCfuaHwIi4jFlpYPWQYho1/b
/7LhQQR7tHxWmusdqlcC0/Ty1QjJXSfcMfsvqT1m5pEjTQjE1t5t1htCbc/ZAwYUASly8c2RqZfG
2OSYFq1ZTlwyolbdczK90Xeu5BRRgB8Epmp4cUk1anp8OP7BmDF8qV81x0CnhIYBj6Or4r7ajLmr
/ihUHVixm69TqtAzK4OeDM2YovLf23sHE7XPY3q6JSECRKQ/2qSV5xzmtpUoFpkmqcAvljPmNegM
9HWWok4oUy03t7t1RcsrxFIdx208Czi9aslkstCecUWjQP2ZKlYIUUGWmsQG3330PHQ/8e1RhahH
RH1I4gWR8sZCZt6vzrWN41qeo+yhnsff4NB24CX7FcazKg1TlGXAAKpK3vsyCYfXfjd2PQeZQ094
zIT4N+Rci5hI90T4fhVJTUWKOHgDnAOSNDWYfT0ctW8CvsBuVxbkfz/g0i8mQ4LotDYJPafilK/g
wMKLHus1Hb84IRRRb5nxQchuBnHXfIsTV6rRGpXOHgRFg549dEM0PL6pO2efUmZCkPB4dDVhQSly
DY/gDyCxVI4kuW26O+5D8Fy1w8OdtixwNIvCLiI4JX4G2/M+CtymIq/VrKlQ7DgYqJa2L1KRIZXp
PQsq21gKk+u3bOwBXFARBR7VX/KIw7Fgl9/6hD35DqsH8arhOvUIaXhVGkJfVtyimMLl8LjdjW6u
IzuTbkHhSnVCTyEzNH/VlN7eZc0eDndJjbphphnfb+cwKMFGmXZSFl7BeLSvFn61DlKn+Vt9SF+u
FH9jpkeGntYppwCPadzlfmZxv1tnM43txmBrc8kKpM3HnWgKtG7tbT2X7grAVPNpJvrkKBZ9umXS
W1zUmpt4CY9Q70ikZu/AeiO2TxjEs7gVZLWt73RaILbDX0Rw4HlN849hl5rpRnMvofm08BYrvtZr
8A6HZ2ouTxPU0vAYLvkVWWe/gx3drH2JuIy2GgZQ+kjP+NTslwqwAF54bbBDm1K461VwWe2tY0dU
PwwW/zv0jxnOxGDFAGCRvPC0O5Fppseo+zeK46DZfK6iLnGY2ZxHFTjh4j+NTb8WAaFRiLvh1Hep
NrsaFTMGK+RltYPnh5XTxjwFdFpLQM9dgEmUurKSyPMVl6nFscnayGcmoh+U2BF+Ve3sOTmlpyzq
DAN/wDMpAUgIJEumT63WUyWBVfXKrywVmjpag+RPkYbwg+pBe8NMXpE31epkvlz4WRFHtEuohpUb
jFFGmPhe5vuXjzglz8bib0mT7G1cg2rtxo0MUx3ne16u5LfBs2Q5XIhygVMgv3ENVTIBmG2OdWQY
AKlowgqTAaIEpI99U9soAw4f4u0IaPnmWBpls4IR1iLnbjc2F4DrNd6lp/jNhbA4OUvA4rMKIHyR
ML555hPvC+r8jN9ovqH8QucVPab0TQEbH+fO73zBk7R+5H11z+JpW6WAljt0TRcxMLdYgLszjnCv
WaS5t728wZ2xHDgmrKyi2c7n+f/ZKIorhON8QH24LOkMgI7nkiFnC7AYcTkqS2Fgwt0HWnMRmdQ7
l+lR0aNgK7vholcDqf7hW5mePdYdEqs07Z6I5E43AV8QwErqhL4aoNH68ellO+p9evN5E1qp1hBZ
KK39wBRGyy+jo5KrM+naYavuSDBfztIyezU3gVv2fGLf3hmX+wo/l4WGw7dvfrh/92TafB7Zjka2
IP3xO8G+qzmM0g6YtZAHloHm2FZDz1xrYqgeDdbPwaHnAD1zBDyH8zptr9LZp/qc1kPx3x99hka4
fj19W5AZPdtwa/bcL4WCGSw+MLD6rEhxLvK0JMvniyoPxq0MQuyaOvmHXZAHnkQzoH0V0zC7TnMr
x1wl1pMpY81W66hwxQMcTwNElOf1tC7vPebZYA5W0EECej3QY3SqA6O3iq7upq2cAMljT0cHtgsk
ngP99878FwK+ov6VXOAfCj7pp/Cbzrt7mJ7cv2P0q7bfTgxbjWiivjCo4YLQDHL/68qGD1wxJ/jS
4NkdxvAV69KooQmt0aiTiCI8VkvKYzITjCV2DfO1hNaM5FyKcTwqE+spbAwVRuu5HioJ29YARmeH
2HKvN1MfOJT1pjNwIsQSfQgpNPrT7cjjisPlWKpO1lUk51yHzdCqIWVpFh3HtTk3c2FdS1/KOoPO
za3Vt6v+CKPnBn7ZEMXbZX2clQTDATJX2KZ3as33DAIqHME79f2rnly+4YKyioy4fh4b5y5QxoUE
f/hniww3AzHJMnu2YCbrPEg5mNVjl3k9wzHakS+sVU4cSj3QrD9SYUewJprYKA7VMHNN/fH0ULPQ
2cezFNq324iSaT/MgfYFaNoYvOQLXf6txGxOx3wCD4LaaXKvo55+WqRoC/7rScqdf/R5o9qmaf4R
rKOkorKL7foisLZ4vCqEu6/qTWcijhC6KlDRB48uz8BfAMDsDHfNfmIDONwpY6fHiQhxWhX/q1Jz
p60cfvM/B1A89e3fzGFFekH/2LNXGHF4lhv3JCJkkqCbj7GLq0FPJNaOGk9rqP+QovWALCKz3O6X
6K0mNJvqbs+ngrYULNDzmWkM7dNsiXeTLJehdyDM3sJeZA4zpink4mFv4kSPGaFjs+1XCJv5iLa8
1nbSuC3XNWFEqcivdtKqn4JokNIV1e4ZefyNi89kAZNdl9pZkmEEaG/8wbk1d8Ru8aI9gVTGw0s5
5i1AXW3pzDZI3PXpE9WMYUoLdcVmg/TP/N7tDZUrVRW1sJa74SINroZMsbYpmNy5pRFjyk9yb7ir
QlafzLsT13pUdk0EBHaLaq6UeCQV/jm5adgzEPTUp+nvem2+ZUI4LxtNP68aFAyxpcX46lcGkOV1
GUEuZcFxvYpB837+2isiCr3C0v76YdzKpqVVl1c670AqSAOrpeMidaGv4jMFeLiQd3QXLTF+yaLa
9cYuwx4veHEjjrZ/NRvL4fjwgOxgAcvcsuk1w7ea9GkU+PUXEw/kTtKfc550dz+Ktv7tr+FL2U0G
8eo41Aj+XggJ9DUNoKBw+mfHBB3x2xuFGsEB4CH+srzYVb/h6gpPlg67AbGjV8jxcaeDraqyZdrH
9rihnUIRVciwR1mDfop9c9rquXQafAr6/ssUTkIM1MCbBLRVw6O7WqL0G0vLDubCGy0xPiabQ0tV
O+SmSLw2z59ccmeS05ITeqc1EKwihHVtg9U0bYQbvzKEC/ohGM86oQNiFdyb1HNP6AX0skPWbjGP
C7jhk4cyo9hzux9Y9xSbpIM/+8RKMPOjZKti0I4rFTDJragRjy0uAKbMw4lioj69yhLr86U+uY2+
GviFXyH0xKerYYe1vaGZ0uhaBO74A6dh7OqM2nIZigjOA5rKsukPU3iJxVLqQ6+GLyB3uFowoYj6
+n6vKcJNdblO6nKSOaS0y1lkAEFhimvYW2IHnK5eVYlGaZ6UB906MoyIwntVIBAzz95ZS7UMo9MP
Lu7VaWKPOlmVMYGyl8QESSJxtcptgsD1hSVqQLSPemR3+rI+LDhC9jPhei7qsNvtePklPpfzIkAe
wgsD8jsPFdv+iA5xmilg3hcvUWP/bbk4FgyKqexL/L3blbrBU5oDe7qDOKQlwM4qfuacL8DthbYW
Faj1zkOrQYn/XEgs9RI3YNw1LiMj0qbxrOjKlyJAA1rOY2NdPg7jbftvC4JDwCp+nZHQNqg4/qeJ
EJC+YfMeEARAYSJ54EiCsfJZgPW8zc0mWqd3FVFNhut/vgcxcnjWbX7a9+VKgNQAAIkWeUmHB4pM
/5J/s9bcHKPq/uK/zU9mODjhG8cCCkuM4TC5WIVE5e6YzG9huyAqSrAn/SQLGlkOrOpIVwOR50FZ
DW9Tz+PGApe23XqIN+AYVhvftPkxvwnM+7LLsYOhKp5R3ZAM/TELHmmnj1hG6yCpBk9dVNHxg8Mc
3ALyayxhcVloojjDctZ/jThg8GVfN+uimntOn2uqwphBIiv6YZAPRFcwy8G7AezenHDe5A5m3S/f
nsJcDqCKncafOMSlk1NUVRF86J+H3xTTG3LvsGkZtnM2gGuqoLtDTv4PxXWxHKFwpxBTwFED/Wj0
oPjVJNYrLH6nPS0hHa2fJ1ojsAK/1fPVa9YugKwDNrrpJQzSfPWa3V42tT8JM007xh0tqu8KOup/
iEMhCOQRaCOJniRmDnMVupqR7cF6Wu9wZh8FHPZmSY8XqYkdX8DtDzJ0VpygT9AKyC58mnGRNpAZ
tk6JhRIakXlIBfZShREohTru/YbjybU5EoCgR7fCo2mUHSp+OCl8eIyA+JSPgc4foINBFf+ocov4
FNzpCqgzPkUgeohow3KDHLXGvLIWr4s8EJkNap1XDuAU3mrnGoTTOhFlHwXUJS40x9UizOmirx0i
pysKHfivj+/QsHzIIGPTzCtpji5aQ2nqULMbQGhWUm9eVFZXb2e3G/JZjlxgxcn5+OYLiifh5Cg3
SWNwl82LN9csuWfgxpjiX5ZLMhwdO6dr2EiEfPrpbyUoOdLqPoVfJkRyxw/F8SMH2JW5W9GgFzEa
eo5OJNWUl+hCB1nkSEHJlyCDeWinvijkjS8fqdWjJKsHQ5g7iT+BdyyaCsLr2EItpHA8umfEd1JR
k32qeUdZ696CUQcIpt/A2ewcsZS1G2AVuKnR7da5bASh6/te3vTFdU9e0hcQYBoLeXCaemNph+5Q
ekstGAmtErBVxHdCWENDxAo04qJTQQadiva4wYnEr+kHZ5hkTfZn6B08MYg7e0wxd3ck2f32tDy7
rJd3paHLp3nCaroY9xQ7J8wBqvQkDa8mu2RhI+htjBHX72RpmeX2fD5rgYaIovT4MzXrYWHmAfEi
SCV8zbAwKiAResA1wS/WLenGjtrf1gUEGKVQury+35wJreswk1e0lm7qJdT0dS4yKTV9XMUZKs6r
4063XF/ywhbOSPBvfa6bPWxcS2IlGeMn2MwBsrZ1NXFmvj3H2Fru42ZxwJw21/gxaoG+UvSSzIYF
eIJrWPn+/ML1Y7A8Zld/QvmL6bToNoBtp9vR6va5ud2QqHwXz3DrDb4MP5VcEf8Cj0MorYCaTsbI
nklyFjzdcB/wpBAiJsBWLyz0XjG4MT/czBDB1rdbXM4pSL1Knotpfz3FL9Eg2qFTdPUEJa8juzPv
FWEOlpcAs4KjqQRZJ0aJD3PvaS+uzFyWUyX0oXopshD1qnppvT/GIhdGd5QBfVw4b+oZZtI6p80B
PxwbxnMOBOTF4r89f08tQhStoT7P9jumSNm8gg9p8nzRdcs8bhSOtBHOQ75a/9C8Q3AeR/m8oc3S
e9LPPE2nRxkqmRCCDXY9ofD3s1LpmG+39qJUJFxPJYuhrtVdWA3zL+8jJ1epk+QCXtXVTE20S+w0
0t4A6S/VK1xxz4tbGsp4lro7x5XfPp28pRTN8RAgJkScFrnQg/MnxCVDs4TUf7TjY/q/n1oWYTnx
K5akXmzljbLUhG7Ufnoi7+b7Xv9MdIEfaHsnGsZpfv6QKq8TT1JRu2+eJBclQh1SYKxKun2nFbIC
dwSdLOc2FfPmHAJUeLGIH8NTpufT/hxXJloUbzAdjVaPijci+6aHWXZS3UPlNy8hZvDLzv6FuUVd
9+KI4SJBgvZRG3yV82GFrxSg+vHT9NJ2E3u8S2EejX/iLnKabLbPVSHHrf9+p6x5k3d+HGlyU/28
SfwV2Nm8boFdJNirhZptC1tG5xnP3wbk2MThCdHZnU2iS6EpRKogDoEjAYyQyRHenBkdwl82Rhtb
mKx8iIbCzo2Qj9cKDAnC8/iBTodkPabfiEYUsmhX15FMGUnKW6vlPQQKaPWg9j+25qd+9PNDIJgq
Sr7W1eJC1gYzAHZS3Q+ZrooAlPkQ3f08ouoat4Zg8btqLdAck8YGhpt6tzwQUXVOdQOfc/GekqVM
UwYyz40GjZzPdHejPMENV9PLU8a7vg4v+9OgXO8SXroG9+scL9D6OkzcZaeJpANimNsijGTitvO3
RXzrM6c8Kh3sq26DF7crJmiRb0TuWQ2x/HQJAMkKXlvgiPhS9HDTnJ0hb0FMcTkdnn03KWal7wU+
3y/ywfw8Bd/3CGKJqn1wOi/D41JoG17CIgc3voF0CNhAjLfW16uGjNEFeIEs4O7Zbf8ERYY8AE2J
QvsjqMSQ6Fxf6eJQJf64HrYTazNFNABjX4lg7d5WWSHNO/YNV88r6xdRlz78YGKK06L7C7zlhufF
3QE5PFoMrIraTdlip1KS22QodDQDEOOFUOFKahX+LuOfSA49v2eDZKA+M2bAhwJSSyxNsnIg4MbH
1St99m+f+3cwIcQPJGfvrbqREiO2gMVwz1DHusBCs67SSp6MdlrhQ//i8aOsmHUYsNlnuwQLNraE
3NDyAJSYCbQRGIjzbYPfeEEQaF2Rbi3zdbwEZXfG8hnQOVQFh/Bw8fzuxSB60szn+jIeoctcDRbY
2l8JFhJCZ+6WYze2fz+jBX4bgRfI4RPNqNWFgPH9fW0BDLfhBSTwJerOC3GM8XlLe5tyGdzwSS1C
6Ug5XL3721VMRoV1dZnloMyYO+J6qWXdvOk18w/ln5VwXdSN20y7zQbE9OBEjYSgO3HutI2CqIpb
sSW8lmEJ6cKbR7Nl3FhNrf2yGSMriM8eGg4h5F5oT0jYA8exitox0d3DysotscmI9Kk6N6jOt0DN
AUenA/vmGHBWHXcdknX8jMyFC+Qk2lHCccC/BwgDBET+Qk975CxtCXlvQv2375dtzR7baE2pTIw7
cypwz9mW2EgAJTDA5m0oidSObEZqNAcyT1hnK5SxN05rUbfqfROw/Hc8H1Z9U/3IhJxVe2PAL26i
3WTcVIUGQ+o3UwOxuQDF7q+NE2nAODRY7iegzv43ZzXHbfUQNt9J6iAjTOBfwJEt7URnpMet09xA
TW0YtzDxSLMnfQJhJPCuZZK13aog1LykNkTm1W4Rr9gE72Bqsc3Ww1fEUtXEZEXzYkweQ3oH93Ij
cHmGXPDM2wbqYFVJu3b6PWaeeJ1gj5W0ZiOcIkEhz9xPE0y48OW0CjxDeGiRPV5auF6u9bsNwuOV
lnRaZA0Nn8sWyOobPQAzj2fwsw85sp51Xz18SVLOzmh++AN/kAgaBpFs6VgYGnbhPBN0Lbjmdi7M
IAVLfCj6sg9CiISd/yVfZXQjdX0v2+tgvC1phPScYLbNnKQZd0I1CwOWUpOFXzD0CmYjll7Dh02i
p1pS8lLB2Opre1UTv14xELYmVTkMHaNVPk/9p+qYlcT3Oq8a2jE1D2tlA+fkg60KH9R6SXHbsWYN
iynMMk/5BQ9rlDUJvzV6RzNwaGt2ggiOLSZO3GJAY1R4fQM29o3XalMZiJa0BukkMN0qg9zbVGX1
QyDleTnt864eHhwqeWDglE+0JciY9Qx8QSJ0+oC72RgAADG+kXT0Oyq0s2yY6Dh1vK/9YA7Wgp9d
u+IruhYFSUBN7gwXkzq3i4y5CH+/AouWI3eOGj+BL7KLueT5rMqlNLXgDFpPtOmRpU7hk3DdYSCH
fqzH0XTX2DJpsHrXmurbsAyJfoSz+ZupLxOosnDKoa/QE6e0ZbevYSJ6rAnpoGq+FEVmTjfC9rj/
zUm8UsP20F0DvQ3evhQ0S5EZH1LDbsQ9Gw8tMncY+TcHf5angpBSdHVUSHfFqskkraeRHAZERtdA
ZA1pKZaG+67l0Wgz5hJybxVCtvE17uimFBMgwMbT56Wqx7cFI7szjDKLMYlcjo04a2EjDvBVs87Z
FcC/N9WNg2gjJ5DALOGnFIV5OlgUVkLPVMRIaQ+zBTXXnSh20c5MvCt9k5D3qZW59ZZGkD915T/s
xD176s2gB3CO9Mnn3G/GLKy9vcI4k6ofYwb4h35Kp0ti5uCYxcfzcBWXwHRUnAaKUemjeUKwmu/t
CjTXu3HWOTCczsOggkqmcZFhVKmmffOX0Uh4rbwAKH0smXLJs353NLRha15kHgSC4YCbp+xNVLHl
RHckNOvvBN8fNG2+Vrdx3BvmAKqm/Lj4X0zMygw4ACDMhWrZ/KvzF6vNL98Tyono8fcpY0Uu0RvP
+s9NLcmpAQ8FOtSBtvu3co2aIkIMLRXhmt6BeTcK0TbZQaDgTai8K1PdtpketCFudxv2LFS4dWNx
bWnn+99bxHcOKTVodzsbNYnckQ3Rz+ztE7sZzvcZWQ0W8ezW96zPs5fbfhuR6Jx+HQuk+DQhYUO7
aUAN87+dQXa/2ecI0Qx+pnu5xoHVLKN3bYAbKL8AYEqPlOPOFS2b/bbhwwDIamvlDfhFQvGM1d9l
MMP3AUZM5goOpCYvglJI3wLJtQWky+0hhnsPAZR/upL9VV5ZJJwkhU3y8MWZQoE2P+29Ook11riD
IDAe3FJTgPVBKVil74+d1r5h+lVOYWMOCApnCNGH4bzJowLE83UL3eXweshrLUDYxXALQqikUVdO
Ztb75wwNrjqiVYIN0mmMaoV115tEuEsm7RJndNEsuClEotTbRNIIYc1dN6/Z2NtmSg/0w8WZ/ipo
gAvIafqVg1C28LhPR+88ESL7gc8sy38H35eN9syS1NqGnFrpqmFSjeW99NntoOTOO/VeDo3SxQVc
17bQP5PVFJcpbRNag6HhwwEmkpxxPQhtPHEE0KW3DdXmbeMbk4aShICcIQzz7VkC4QlLaTEfB8OB
OEJYZG/jAuBlTfrucjjiNzBPY785BzsA28YbQ9yEx3hDEmzJ2cKEHtrnlKqicvXwTifKLHqumGzy
RHv4KKP5hyR4YutfpUwrg8XbGoSINkv8xVybnlhsvAMUXJ1EEKOO8U05L2ZNXkv9hfVGy3sgSiOT
727AP/p9kc1TG0wp43yTCKOvN8yUr6OR9Hg8VN7JVIeI2NzPuxEJb+YOqQkoxQFFsh5dT3r5dC0O
QVw2b4CYbuj+Lfw36CoaAVN178AQJtSOfs3HkI9AjBBnZhrZBmA3+pgKKZZO23zDV9bTspthpHZM
qa/hTg4Da8DLGgnWapSe5ekMokjG4rArLMKS41MkLVzpMyRVRDIvEn+iwgLlTRYwRmFbi/8Nm9LT
gVyMdn9/q3EAzeSSUJn2H4A1dCz+y1pPQI1gkTipmTQBaXOStiqqLRwu2KrQjYFzaH5G9T9JdlGD
QpG32YCpsCT4wUZcQQ++IJtwsm3Gx9lRF5GTadurUOlqSWWGYhj4p0JME9Qy3Viu1xEKqJBT6erF
r0MKp+k3GaqhJfFKlxiBmkU80zzHZR+hRKAPRszg/y18MbaPW0xahyYVUsjeQH7NTREDfcb3KA2u
kgVzpjxZuGcowoNrV+gBK+V5qAN0/tIFDs+Lxkg36OCXvGRWUC41a4zwR66WwrO0JNb9Rd6erW39
r7p9YfyJL+6eQ6Amg6pvMuLK8OA9jfnVHBEx0wmPnBEyLHrXRP2Aid+LiQmD560XPzwKJc7EnAvG
0BC7EA4U5rleLnX7fbIHYsnro/nt+2fvDXu+91HU3iNA1iUEErdOEWLqBIhOWTtUCjdOz+hQPfag
e/SUiQs+0gWPM0KLtIWAg5fyEGBzUp7+Pdv0KS+PgOQUh/QQ0P4EBoIHB3p8gDFB1A955ItJO5lm
senpSSxqL6lV/i5xndg4pxjbRYMo1FbO5gGxn9SE3WUJp7Bqunpjr3yOhdTQmYm0Lussgn1ZxQWg
jgPJN4tLB3QE+bQEV81xNB0vBeb1xwDGCNMwQSjAjfWShET0eUrQ7ZGSBxA0v0cZysU16+d/SKtE
e0TUhuxUPEdKQprTSuPxJaGU2cB3+GfDJoSXSky9iYCyGqbKYH+6A56DPhcB/o2R9DZ79qOiZvry
yC4xPdaDrR3ss9GsKc/h4HytRql4eLflzbjF/qmViOq5CgVngjO0GfT7AbK/8iTX/IwNgaB1rOfl
/xAdALg/EJeZ5R8YtNZs32qdtgfu6a0lMGpSeBKNckskP2+iHyfOLa+qtwcvUQkKft8TG+9YaHD8
JPd32qS4l/OORI7/cBNT06csU1dde/gjO8q64yIZBYDY3IoiVqxmhCrhRdvsbOWqst84YHYqUzvY
nm60N+zDXTogpjumR4osOjpKBily0FBKc44Jd/oKumiEem7mkl+jogiNELXr7NcRCZvWpB3KAoN9
+z+PoF+hjsHK444QL7p9BMk6C0mo7KJOxX8iNtcNnRmw4Ed60Ve3gBcPQdGf7+FGLDH/Ssc5nKVh
4xHgz2glT8tRoQL859r6r0AoCy//RvsM22V0JMvifzCY0qYOvUDKIvDsRKPC2Gks1uZEFy1qGP12
ix5cVR409TDdsvNHdb/8Io0xcCsjkxk5cIMymfguKcZS36w4pe8nRPdPxdyYk0JA3xwJrm35Khmx
Lagat3wXW7T8U9vDcmAqMxJCaIuobm2G/IyIlJkOYv4iBo2v7dtblwaSWE/TGRGxZV//gcqZWArB
N8hCl7WxaIhVl5jv1tPF363mpJmDO+CIKz6RRktxcL2bZdcSDy/yaz2AOf8gLpekgslz/NrLTBME
hs3uIjouA5VhU5KjSPYRGknugHWLKlEv3AViIaQlOOOI7Gvn+Vr2ppn0Nn+ivSZVWJ5GjFaHqVEy
EBq3P6rWJxH33JO4qQkMdZVwKEqD7GRV0pPAbXeL8wOgKq1RCa6kb4xnbfS+LjRqNsj869kv6caJ
F4G5fywZTqxcDgcMJ76rox3sSPXhgRQEfXgxdN2gUiKIMrSk5GYBUpiHGzZDRSV0e9IrE2lPdmly
I4iWF2X0OUKxyvc6NU3DXbnTNHAxBYOKKXanFc1gujzoB2unugacJ8S/HebzLn9gdck3SyyXUORf
YRerdRgPODDzuDpp27GAHNiyRL5EhnSAHKbGxfagQjNCD6Po9n8kHojp85Fs6NiOU+awfqOJs/Oo
s9atI7VTau7ypEzyw/HUu7XQqreYtWXyag5MZj2jv9ITyPkeFo+z39sE+bx3aj+rL50/Zst5QX0Q
+JRBS4m4In8d72IlGNJLtY5uW/RC1k80hX+kRZtQjiOKoCHFE9U8kgBrMDbZ3KNhbsw3J+zrXgd/
bKZCa5MxPd3AhuazUs7WdTcfD6KppBHs/+sfKcoaMoYhqusm3KCTp4f7HhC+1tdjgpxszhuqOgyi
ZhqfoiO7m+weeo2nt/r32c7hLoe9rJ5562mdeEyx9uY8PqMSu+AgTSXXOo5Jnh3E8zfm3KjABgQS
AkehM96QP721bDBumNcE+EbZoo9Rwgd40Uda9tHoUwIzCqpvtz/emNuQZRnngq7UoUz2k/lw+hq5
lj5IGvy329DHXk1++gBIOUQLA2eDqqlD0Ei1vvTERYMxygazwvIPZo2qM0/AZ78/tSj9MT/vr3nk
KgtipYaEn+1bhOqtUeVH6LXo3/r+aJbSmAkk/Zpmwf3+fD0rdytNlNhdVwgHKWL6XrPt4HxCaYb/
T0DpQGxiW7o0KcWZdk0p3l5SBLiFpiR5BK2+qcVVhzVUW8mD805qZFm/Fgs1vDTcqDsiGbWk5CWR
Vl3QAGHoXBd9JzPg/oxRVBa8+3+iGZLNVdp6oQPVuiltLeCQKMW93n9YFcuK2tCrIDeWdPgdFS4N
nAkbFxYXgHbxjLcjhYSDfWGWxVRTgCG9WE0JLataFjsurU4a8BvFKBBFh9W80b50Y6cj1N/SIsjm
i58fg6scXp3Qp85hunvhFqQiSTHcsXthAvXoIGT1OvbwiTA6xdiNpt+2bU2WM4pvXPuOhzxKSnVn
TiFnSov9HLJMFz3a3jydWkQaj75dW0N8LOHE5cyyaQbKSfCSAhOlFpg2kVf9HukSZw2sHDeBF1BC
79IVdzRPT6eb6jEsu97foAnF+0Wty0imz20jHWEO3pvRmDwPSliqJwux8LsTLAwpWWa5H9N5Odz7
iHAPMOADknYVPgL9DQ6HXXwWcfJ78s0PEcBWbhOhBVlkAPs++2zBUJSP2rGcX6GnWoJpzZQ034yo
YROFPk36lDC8wXeZVomaDql7APF6pxh1KRS9R/RI6UfzNFmvgMSRWqK9u+mfoQgV76BhtdKzpipv
ADE09oUBqhwjZv8NP6gHfHoWltyfhMdhvEiS34OLOFqgJ3T7q+fv+G30oCKO07rvdLyRtQXZ230v
PqlHxwLhbkmY5O2XanOuXUeOWgeHzAwo9O4eDIbUrjaJWzvkrCoHVorfPvIhMbp/7AONOaY3/zJj
XTSgENfThy0WqB1oR8NII8O4pI1XE5DWx+sFMbyVAsFCrkNreQ5lO1AL4x84dzBO4FGdppA9uapP
fQCko3fUJubUt/CYXXMrsGbgjrHvGJHgKEc1+1gXZ+ILAvQObV534FL4FOzVLsEEiXOTGvMZhKxc
CWDw8HDbDKfcDL601X5WEXsDxuGailqbfv7gQq9gStHZqQNil9KOKXjQvMvoQ+Czkja6Srrw1r06
5ugPPM0U3QrMJPuqCZ7jkbPA1gdKid5J09WCmZr+k5YoR6ycqF55tbKTOlUXsHGXgeI76lvLolJm
qYJV920rZxhHnV+3/uK3cS1r16lEVTi5cHuutWMm892Sr1bwOoTmRoZoMmJUt+jMvpV/lDu0+04a
Jm7us0+kMyux+Ek5siME7xPYezmjBRGM9vki+13QXQa4vDJAgDk4FugTRW7vMOY1+qozZyU4PB+D
fxjSDKvheR1GrrPJ9mliUDD7MScEgyn0KVgJ4bJ2RNgPJPZcv3xPa2HWqhyh72PYnCox3gn+U15k
Z3FJaiW5wDp2Mib1KxzUPPNKRF3puNnpJ3vNdiCtx5y+guW1qgcfWLOWtrgCyYRDkrqyc+XffU90
32ykXgKkeIi67TE1EJ9yfcw/BzRQmse7T//VA+1uDdEBcqOkFqkUoltP+hKgL/sNxTByc70eIrIZ
qXFQN1wOuZyGj6Pm/GIdJ0OGsb3L/sN8+hdaItdD5EqFvnH7g/e7oaqAt08trtxMcgDF5VBuao/k
aNjdBR5hATVKQWTs/Kb3/9NM9fUSRM9ZbzceJtiFVKiEMSVdM0yHimGsif2aRrD9a9FBXi6ccqtB
LCThUXaCen+T4LhS2P/GWhMGED62mCH+dkda0rafNhrIAF8OQtjWPOiJSWN8E3I8xi2eXQSaCv/9
J/q/RWHTXvMZ5FItllNUTuEt/l/gxgf6W/+A94NLhL87Df7Z/fUag20kBFf+t6OJm6uNHFKNF1gB
1tCCZY0OAPzh5MWMolrmZZbhF9wRz/aSB6KwGJzO1kAL/7acDnWf5yzl1RC9KyEjSvitGdWQEgSD
PwK3EXAdNR1vjkHjjRxca+iw1Yzjm3ylEuFA7h+WzutPd929/gHhJI4Zjg6fsOpm4d1rx8Rh75Tp
mbxddMIoRwLjGtNTHeqZ3PvxT6RMRtBJzgzBi2Rt5NkDRsqGNn6JI4CUXidZzqXzUVzwQ27j/Zcd
m+U2xNVXgUoPZXolyGSHFdxmn81VwgTeRsnszCjVr59+wzoUDbgQ+R20IB9sRuHS2DIEF8D5vx4r
gObI1bSbhAuexAfDCixvNBdY7LAcrsNTeKDCiw727/tccGzjWNT1BzOaJ+uNBDDgwUgJ2dxHCQgu
vKBZ6JNzRxU+Q/hUQvOonDi1LxlfzrfSJON6JDWRm9mXr8EJ2KMYdCoG2q+x/uCyiIcxIpeS/8GH
n3B5O35pXa4lDmmcASjcxF1Mp77gEWSfOmN2tRdMKKshPVRIEvgvbNqyPYUkmOw2qjbn1u1GMdbn
pJOfbQyrCBmXwKyJLo5SW4TnrJQ0+W2JVTZtLCXtn5GMEYnhboPaYhQwTmB/MOkTQ0WStyQETBv5
afZC66aUy5m2zDRDZscFNxk5lgQv9dKlhN6iEAcLNPXjQmTr7kj+0lawT9NSe4eyIn6J0RK54ZeQ
8TEG4ToLhAL7HF4510bKx61T9ZTNTe6CROq3+Jsc4ORQGSCiA2/wjhj+KOJKvhk8rd33n1lt8oMl
N48RhFezAr9csWcjAoQVfupXN3eP5QgFjkVFd1PYJZbehcov+WkJsgWBVvjrk3Z1UFc0JbETNsct
UpRVM/0m39xXHgatKbvugkx5Lu+cM7eJf7VwphS5Gk202Hh1T/qTQiz59EirP9AWqg5vLlR3Jnol
xENbk0nvWSTAmoYtiUGSsrILZdMgjDAfZegKnAKjIvgOEZHc7pRGRwIfyIYQf6cWa1hitsxh4g4i
93YS4hhC0GuOMNMSwJqQb7n9yBPaPHfXuV8URfV4O7ixUGLO+9vs2ZhOjPSMtb5/nDkwhpnHGEd7
jpD/7hhCwWJNC+2A8xwSDNrNJ+dJo/9oPqQqtPhFGTjTlz5syBnLKgf2rE5WwYKSWq5eVkrP/zzO
jNisWWqGkNDYCKJS1xtXb7GYDomiDOsM0OAyqeOjkuX7C1eruVULgBisEZIpBiZuk7cCgPMysJSb
wEAkbn3sJsGlMQHIGqJbn4J9LQ+gIzdR4E/51tG9wENiCtFWxzV4ApUY8T5CMmQeDq0MIXhwZGUM
caV2vn4C7y5EK5rar8KldleF1yhEgOOJb9QpMe/fYpZQBbCVVo8MRf+MSLKTE8Lthg7AQ9z3vJ6E
/lCyfWVUy+bgLhpMMaPRViBWj8IECi9FR68Dqcc4rfPRCifVCH66XUS3xikdE5uJ+EatWdTEcLo2
13Hb3ApllUwkzKahHqw2eC9UvAzFYqz1AGrnL8PU/SArMdjr3S9d5I1te5bWi2gtP3LOun4Qko9c
F43CKK6MBgzIhKMHtM5qPIzKR6lqEcJsBRb9cj5syt0HWC2etN31tPhW7quNu2ECtZv86AbGYZYw
ALtJ8Mw4owyiiU7FumyAm4/twpKxn73XubUzycme1HoA4eYAy8QCTH4QXfnxw7YKw5zSgYb7XwT+
kNldURg9NMif6oZd8Z0LlZsv2/lSDeFnowfzQJCt/2a4O16LeltgZYsu4mAWts7d1G3s0rgmu8V1
I1xx5H5PMtH9M/WgSK2jgiIX6RqDN2ZZHJpfdcpSCBDDVIGxzVhM0/ISlPPyE+HMxRHQoLPPaasI
cCyJ5vcbgKrFIW0KzoUHPBU9Zo47xFgOJHrNRsDaOghxfuqHshvBeRrY73exspKfecj60VFEeRuT
ob5ecbW58zw+qG25+xf3u1Z65yw7j6MeW8Q+Wtzg56CCGJS7W8d5Aw/bGFcf4WzDhiNG7b7eRww7
RQLbf1T1MZcpdoprGLtWJcOyJzN3mg7BoQ4Mz5GTkAgFHj+1m90sKClNvBMioMp8r+2KAzIx7DGk
+HoQYJjlqeUh79MY9tRT5j9Uk5YtG2JiDiJyxVitpo7RuCJsP4LYClqGEY+1CRw8ANi0Hcrm8ZWu
fYAmHWELtV2vtG6sGXWiOAJBCbFGD1ckjAvoh7RAximbc1Jq2IDGOWsFfuAr7wKIi3rBOHgo8kFB
MFyQLowBGSJMgpVFpTRTkg7Z82ucGV2JT6JpS5Xp64BKHgcAZR6Yr+ixBF8L3X0VWXcjzKyJuQrR
8Ma8iydnoL8C89NQVN2FnAeBXESR8Ex8TTZcgc5umI/JcmSBVwd+twhPrzhnr6A8yHnzgNCt0UpD
U1IbA86Q7xJ6di8CpjL7FXoYdg6EaG3xqP9wY3iwtUVb48xWaAWuyaZA8pgOU4w4VTH6v+coQDuT
Z6KWbl+LRRJ4s0GiwYVfdTnfYrThsCweQo8f4WlmoIjqHl2MQlHEpTYluW+mR8vb/WLmVZP+MTBy
BCmW+BSZQyvxE9psuoju7w3cW24+AdnioySdERMd+p2eu8LeRJZ0NkcrGmCijhZQfOWJmO26jpg7
T0i/APaKDjpcIj3Q5EH2dZmLk/KwSicHEDqhdmmnKTQ/eqgiYFn1khSuce8n+ZPm/mt7zr1iF+Kn
gzF8JC5t0xv1KnzTlaQb/Y8otvno133g3W01NwT1sPyvHkCXn096Fytr8l5iQP1qfrwexlxS7G1Q
P3AnQWVeSj2EOf/RXh/MGq/OVVC4tJpYIjf0dmdV7s3EU5a3pVoAILs+JLznREuxzJkR6WxnUHgt
EZpn2NH7hAXUN3Qr+DEyiKLufmYpq1GH7cWfEXT1ypZy7RTVyOjboMGPuP4Kzm+S3pl0mL1OEPrw
BioOXQ4NYcT2gd2R+0UFHwS9zkAH2j+VTtUwiPTMimgFoxWzFlE5OcdKTVb9svN5FakaOHJ2JMB6
aD7vb/WSoEn+uBvmrB+9ByHy/X4IUQoCZTvQCvBlO6q8S9C9/GEtdmz38PFj7BFsSRHsd3HCL249
bNKQPrZFPRSZprrUfEx47FTqO7FG6Vx0MT1kmNDwOw8ny38CA0IqQEdA+iTTk0TH4DP9herVx4VO
mrj2VmmiatjFzhhI4rNbpSROk77Jvrg9bMr43a0c/uEjuckQifxamFiVekxc/X7sXiemFwe41LXJ
S67jc8I+GLH8Q3tUxzOIVzphSL8CJotBVYDLCHzTkggZU21E+rKt/uGQo9dPR8+6Vd6DvLXM/5FT
lW1ty7tfmQKISKsK4X1hjO8+6Sd0oftnWK3Q9SPOBR153hZfqQ1zidbf1mphQa/Vj/t+wHXbh6Bc
pX2KkRaCrLAx7AnPfF1EDnRZyWy7s/PAAgDtJwzGVnfR2KJIuu9x5jMPKCmExjpRUS91NZVmpTkt
0lDai2vbMFsNl7BF1+aZfIrt2xcr9uSejIzF13rarL6ykL+bmsCsW5qHnYZZILdvmBzK8Wy8TlqN
spsQVnntFge6DDhnPkn7deNNzSaNT1lFM28UxEFIqIhl98b+ybhfPVynYaSsPb51PGf+uz7LkmqV
Fsk5Ef/DA3vmse6lRhdyOTEvJ0NMwSwfw7Vm/eGAEftH7LgdKBHldWNp4xo6Aw2ILsqXYjxAhwAp
xezR4TDPOmhpmNaHfDFHWER4keLesye2ou7xfQXBKfcB0zaXGgoLWydS7FaRO2KAEDVknLCVd6M7
l1pj1TMUJpto4xJg0AFp5+hMZIsR45fxH0pZXK4bRfv52P5FOf5d+04bCklZiSOaXEqrznmnLm/E
M4WTHhIpGmzekK79GSRNvKDRWIBm/Ep/jrvKHPu7i/bwnJG9qii4vr6n5k98nhOPkxTSGclsVgIQ
3QIMDNXOxOUr1YdUOb8Gk41SlNw6Y9UGvoBgAqwfn+O/tMQ0Ep6HME5Dr6XNAxRri3f9Ag5xW7ta
LCUIvXwJRSUKvU4EW9CmFb1FH7pWUReyBSPgV9MeqnlfBmM9ry9azT+IfnAmBpT/z38KUZgh+SH/
uz7x6KTWSn4IYEGcA9HJN+kVzFrvcHpClz3JMfYslEok0lF/fjIjd9fT5bulPmohbnexPiwVp9vq
+yoBCrd3djy6BX2IcB4OJK650vPSYBxVNlXhpcGZ4/IB2me+Y3f/dnJcUOFdFKXpeYM1oLX9IWaf
Zso1394NqW9d0fqx/atxPXu2bFj9mzNu+riao/jTIMYXB79lxbtq1V5V6NP77FCkWRvN/mZA5bGA
VZ7E397Fm+aknVAHEmN8OCiUcAo3DJacAYVi11czSiuuhBo+d/k+D2Fbe9ocXVRyitoOrsOcHOcd
dbdBv6q/9XQT2YBHsk7teDwX30hh/6sRhD+lYbNFAk2Yl+BnG82jjhp476n0VUjQ4aCiYi9gsNXE
LrdJvb9It0CdgPc4Jb64OAOtaTeUZXsVEerqTCKP/Jn0Qg22TUHGDgILh4GOMmCIq8swolTRjzQN
Rjca10wNHv1Ndf6hNv4Tu7zJOXxUwApYOkh+0ClyuD7umXOG/P5zx6lf5bKTCmYPpf4ijDpxUKjT
v/3X1IAJjMLRqABe/hgt8x7av84g1znVANIP5zF13CStmE9VMhfBoLahaISYQsaueC4oY+wy/xTW
owJ2Dfeb767H42yjPoNF3FGQoYvN2I5I35c7wU16tao56Ojm6gPxcdR5w2bibG11N4SiqQcZRTmM
26Cfapf5AVBXtOiUrdG3/xJ4yaeOpZPTHa16+IJj4TgqR0eb60ErBpnY2s5KUAGcWvCitakPP0ot
N4Yzjv4l71bEXnHAVc0LCKGM024Qq7vrZeu/C0VfK6IfFk3GOhUzLNgUMcOuYVnpwKbSsVf7vi/z
3eiQvwMrOMjwZ3jCLlJ8rW12BG2IYNh3JZb54NElrkoaajnumIwF4TZBnubw+fyKf8Rw+3v0ooS2
+UVKynaP3ABWn14azHF54Mt7MaIzSIuK/KS8kNSK7ep9CggnTqt+dcyRRGxvh5iiXr7jXoD9Su2k
aArjutQcmUdh9qap9dsP+PddfWvYj1Vk128tL2bK1+oJG9PcXhgIFZOmYJMABKzS7vyBzVI9vjVz
7a7JXCm0NfrbKbJxQzYqjX+unc3EaoAiTbu+Z4Kobxm2Z5EuT4veyouJhmUirHeaRki4rPiH6p2j
inrK+hvl8DiRXGIMgLMzs5x+iNDrynktocpQRwL/xjrNrkMUO/aby7UfIgKX+etXqauEhhUJOx2A
gQfuykKzamIRZX26wOPz2K3kJIYQUJZBwRR4tXprkecvJxqZV/8s6fii4RG6AbmoDrPrCPYcz520
Bw9cOJhzaONHbaGJL3J+Hw0u6Q+XRVkzkhDfNHKUqZSGwzEMS37Th0gZwPpKNtCYIMoV4Uya9HdM
vSdiyJQInV7TPH2GainnkgAD2l98X9QgFrobhNDMHH1Z367i4aw3kR2F2aSjoyH5GOacSEza9faF
8QfcG7gaX9kT0H45sj0Kbpsn7iSJDOKKKomkazZms4jbodu4TsA/6A19vzLujr6zxNPK2F/3iHCP
iiPQNUfFBzKJaVGCrQJ3IsrOkNG+xJb6EdpeU+5/1gmjoWMYdi7yUszFOWjLVucC6YTjlJFxixbj
NHcBdS5uKeVzSMe53ns4tJWmhlKxGnesc8Sjau/N7pM/LDLxLP/3dU5y0XcnBWp8O6azk+okW2np
9MFRW27tA5338ynm/CXQgcFmqOrWgrakJJl09ZzFJQx+R0DcUzONE7hO1tSZ2rsfvrPCAf0VzPYm
FA9Vw95CI5gAfHrq1njnUu8Kbft5Idt6+fH71izzjWtu/ZhtGim6WRbv2wFF/rTtLqBB70QOzHBx
IGOfRClgl/F/ZLDL+FeHpj9WQtmxbf5P25+ZgXRE6U0nMpXnt9GIy7KJJFbmA6ww4bV/Jnp+Vu02
XZRE4EfvVjM/Wneex/+1K0vEzPGIjR3QI7bB/mePHO2kMkDwrkagrLCZ2nHT3A2uFL3ep+ROpF9+
Xn3GrYCz3G1zSyOjgjiWmobfeXOaowzDTGolv6s0cpqqm+4CdZvUB4mXZiRnrXzmTbA9o0DJn1TE
hZnZ/pJq1a/yOXgTnE//d73EseKAnAHEsBDzMA4s+1/3if1MnMBfrMwd5fGVpfe3t0Oq+XbFWMOu
zfOG+TWN6bnNulCm7czka/RA335rFKyGzO1IpoiXLLdSGRnYF/pnFOj3j4LNPqToPaICmVuI/cXu
3PyPIK0Ri2qtyO4dy/JaX4X61ZUzIJBZMPJiLkyDxtNw5V/XndHQjdeYkrS813cAeLUGqOysygCe
PG4c0JajAT8qWF/NT5lcxrLBi4kt15SyVwQqX69J2m3wNSfn3QVIRy4dbroKPpfEOmD9iJAKgU20
YeU/7UxBaF6JhRrQqnePgG2IPmRGm47OuplbzN63F81/coLxETU8ND01j+ERxVj5s5LAJ1b2247E
dIbsbkR5+hnvRgIcZ9/RkMfGP4VVs4nffgGn5O+xtcedZP+Y+s27AKw8OqhzBgxd9WEmLLl0Kdky
wbg+oS9tgWRYtEJFRiB0dQmjP3RrTqEva5WT3QIfe5SpcWSo+o9f4FzTn8yBKjSS9P3Op1Vyelf6
5cqwn7XXV2x78BJddH4xp9/uchANPrtOxpPY28lBrFOOw0va5vzG7tuBGa2AEh4ICTeVjGmivRWv
fYn0cSQLm5y3mi0g4Maug1EhXmj2itrXNrJXcLZDXqsqHU3INzEOQMLf8b/ruSPtqQxmbZp+3Li9
rz6Q3v2IctGFLIH0cajFObupXioxGtT+EerH5qeeQVnj20IUtvBhwkPFeZSNYUJaTlApuF/Rk6EG
djVy59ek0Nk/7mfKAQUXVTnh8oeiFywRij5Duii/Nhuc5k2U2iBm8Hq2tV50ayc0OfR1wROtud+u
irB0wBsazwoa20B/SuxbbhQofFeOFWCRFAjGLuiBGH+sv04P2XlvTTdSM9VSyRJZMR5PP7j3dWun
qXaa7Z8uQM4FD7fbPlO8lqzjqPhv0UFbQOaE330FvXIkOzsWNnLcSfQgt7wkTxBiXnkS15bSnrZs
uA1vRkM1jp9Rll2LBEMhV5uikn06Fco++Hg6102Hw+nWgbWN1IzeKBHHFXFe2ViHJAOW3Ej8mFXH
u0WbrGs0K0k1KKggH60C54tbF2b53oKpp6Vohg+jtu4TlGzrJBWA7i0Fc5RdN/yU/nHEB/f5JP1Q
uZqHMuzTYVSHlWsbG+wSCtlB5iYNUYZKn6f9/sL7cJ1Qe82ZBVVrWUs+2nJbbvT6BzrywAq/MawF
jBMfC83lGC1BwRBMdW45x5FQvZKMMwl/qi6KN+X3N4qoJPpqk7mbi27ZFBEdm75M2t1ihrSe2jqZ
XrcR5lkHF8IlyGE7xzLIkLgCVLxP7sLwkrJkleI76fsWBqDHZvpskItGjCiAYWHIBgKNKuJFpbjw
NSeA8oxWrM8rkxKDsQzS+a/DxGxGfCmlgFYkrMqFbdgzpoNMgmkDbTUhLpp+o7fR2PQY82IrGri/
yjZrxNxkGOijxC/XsGmq6gQlCwP+tQeOzIA3bqTKlcqzV6vyr4n1M5PoJMxzF9xbnn/4gacy5vBn
kX5iZCX/QOlHCmdvnrRHZ/wG8DiR6HHSe9xNluRV+NfFEm88ZvjkyUX8Z+/tBIl1W6wsz34/R0oJ
qY6Ps1H2FUhOCxVP5jJxtdHMBLuw+zzDjzXBT53RiGnRhEqkDxr+pYODaxogDX9thPjrjy4d4l/s
YAYjIlXKtff70cs15kUH77e4bPtvihR4GKrMM0bEE8NfTqfmSoQdfHgx8vlWn4YT6n4/41/QuOsV
UhloslpQF2U7uqNAzs85RdK3aHovN9Ci/nZ3NJOLN4x0RKPiFWqOjt2gSibkrW4W6B3NtRo9hikQ
Ym6qaqpycSJ238GFvMtQ3k0UGu9iWAtsk6v3+UMVKdSRbrZLz+Yctsg2ZsYPeDkY7ujRpRhuzl0T
rIclWpjKW96idLY3srUA2XK6/mQPI1eL88+UClJifKFXI0qTK4QN2PXj2ZZ6vU+UphRVCEgmv3bF
douVwhU2h52vc54AgsjOJ8llJOk7cSQ8jsh1q8zL3U70JhF+STXRHgcj4cMoVUSwC/7/4E12eHZd
vTIoMRo993WG0eDe2H1kjooMLf4nMA70iGC2RDBVMEJgJPeZo7OxA7+VgJpf3ERahHM12BhUcC6t
zHZTsY1GIKGP+NRTyg54qO5OKQu9eS9GnrJ209w0+CcnLI8lsEGtCfpNeGDw804xfk6sRwd8PEmi
P9wjKOWSzLclCj+TWTtjB3POsMac8Mxg1basF+arIWsjJOR1WC8Igm09X11dt8NgmgiOxdYAbKMu
OQNDZXAKNUWL8K2NbuQBhw5At2mbXNkbBWcYLVWEv/AP28Tw2CS0E44r9BlfqQaOk5BRXTm8Rbs7
1qI6Gi5nmuZa+JtPHCFcVs0iQjtctoD0dbSaTYAP94ZVu5pMZIrhqM3P6io+BX6owPkPoOG7Q1ly
HNnN8wK5N0dg8x8q8DSht4PKtdCuobO0/LDl1aIZCVFu2DS1c9vErDhc5X6IVD5NSIkd+AjOzOn8
Ik5Urn4EXZ8MhxEfLhWDims+O4htBw3vQoXJDOTB4aX8vZgKgDcLD/uT7WWCU2hfmPgnbGUB+ZlH
zK+NqM16SXoEob4VcQ0Ej9qVAF9TBZF44SNIE6Ov1XWQDWF9sPrxctLawf7QSXzgtxO4aYRittSq
kaYyo8M8MAlHUeOX8ityLro7o41vQZlUHOOiQHF5Sq2hFjVM0iu+wrRNiH3UBN62qybieD0zfb8Q
XuaDqjqzu9o1ncmA0QrCsM7M3CPAIqF2eIRmqO0ba5Ldnj8j4sRS/Fwgo6nDl0b/ZeXhB2snarGw
r07091FxUGfvx3pE/W44mWyLXPuslbGr823owCN0hswDgqpApEDwYkDPE3dPM+oHI78FsEBXKbME
SvSd2gUL6WSxvp0R9xAM06e2TiszV3GaEZifeSlNecpwpxAhSDBG83Tx50tlkf5u424K9tmXa9P5
OYa5qjPZnyzwAmk8px9tHomj/1cUiCYwnXfkdcpCNEcQguiuSBnG8A3IikwhfGL3NePQ7ly3OVt1
ri/HpGHyOxaGWXq0GHBxL/6VJh1nZ8/LOADZaRlBL9CzgHXgQUcw8qlayfQygTAwat+hZza66Gbo
wskmwvFo+Fg83p87tquK8QXiDLKXikGwTQPAyA2ko4qfkalpycAm01t1hWjW+bOnp30Ni1XH+0YU
BrjwhG+JoJfkefwt+yJ5jrkrXic0wvbP+xGEeW4M3jF0kLqowZ0Zzg5vaEcpi7XsG/xOYiXCMTTw
waZ/flGxHGJoBDm6kpRRK/F11e7RQxzpPRwyaObTVgftklI6ZgD0HRJSKn66g49KkSGnFM7JOtb7
b4c7INUKpPMr9EmtLjz1OpFQGM7kwGfyCpbRftz3wpPM0fqybk9gE7QSt6EJEQMrmeE8bcblMtDR
atUb4TpdXlUtUqL/lxj4zgW+FbdgEvEzRlZY7J1tCEPT8AfFezDuZaU08hPrpZZWvekB7wbXCzEJ
jUHfjsa9iTE5d4iRdAhZgR5bH4noW0DKtjIeB8WgtEMaFejZW5f/CngYPn8qLe9u00bZ1zCaqbO/
RYkvf18cKpl6MKB9KFTQPcZb96AnApyrl18UxY2afAc4N8FGJ2OVyNUhgGrMylSIzbIjIUIyXwc7
c53wC+ftXTynQE8PLcTvFBLtbTLsoFPlVI91Wb/EXs97pYLCN844Nh4ynkScHA2zPjDDTAHvo3UG
xfdgc9v3/hhfdEAg9VKn3RcemObqesVbqnZ5fETPxB9tWOkRh0ihs6EA7I/JIgLMd7lOlb5bBsF7
lMDJHa6LY288qLApR9tRXLfOoaQefjxBaJGz64fdcgEqKiyLgj4z0tlgCRjCmo0Dl3nSiR383NUl
XmlwGDiiYH3Ty7bUj1rpki1QKLu6IE+um3Ibq6mwDjSU2i6dtamF4iFeaeA9MtC9VMFCmUgGPTt+
wSdwiAlBd/VbwxZyX9WjYZWHwxLGIdi2+0pZUCWmGTdL+mDjz0T/k3q26kM5nbbzRFgaWFynzdkE
jy+PSNZD2WLRun7IFrE+nd2mzfv2rL+y6eLAZffrlk1/RMCkkDKG76wwmTW9qinCXHVuEs8OIp2h
QkJoNvF3pUCJ/IZC6QiKSBlfJfauHC4QaKzrt9FZrKcnNMJLxwzwRBCJMlvfnPj7RTjY+RGzJ+2+
ZeVBURX6y2/Yemze1btOUICg0toUNz7w/WUVGXNI1wM1eDSNpPZYE893HXwX1e+vuIinn+eWU+Da
LBemZWA8vAtu8lzMAeHLYiAJ+X+O33nfjzS6MExtJVvfzdWMrPDqfCUqMMyz6WgqARsoIOsixYbB
he0WVeRcMlDYQomJNWGHDUGgORgUCXqJauBkuYD4eI+1gkSoskujDHOcNAdsQh5ZYjyIqc1l+Qng
KmhDAz6064dEo4uudnqF7MDXPyJtwzmdB1QXlbYYW+GzAHMcTF6Hn2zEuyBnzaTENdk350o8Yfwo
ArA3PYUs9qjDj/RS4gLlRkonjQCs+J7jvhW4xrcuHQoPh3wKfJaI8fAaqotr1b4SsXNTqiSCnKYc
14Yj9mnbCx4GeFzJp5r7CWK52g5N4/aSwKxANFv+8QhzkAoPGXKyhoU7wOnNi0cZZhge1D8EoBSt
Kz4ig3JI5h+EoZt3fQiIBiDnAEm8m+d04hYX3nj+Oy7vPzF6NQNHZPSthWjEjHdkJWbklMAJbB3O
rWyZdN2TRrBkcVGhwmMnIoxnz+OKQ6q0fbE+ceIZmQbkO0eqDBWiC70cgwfy8s4hecoWBeQCFEQo
5Plm1MjF07pJXaq+EJmOQU4U5dHpR1E/AUlxsBbiMWEfGAaG52FtHjHo5lNbFLC3S8otcsCx9uq6
4327RJuBHiNmRzL3AkXeeUAk249gwvvu/B7BFShXlWcJ2V6mv0IO8vJ/ZvfGAeRD854EkDm5Y3s5
P6BJ+IeXgzwLaFYtr9rKWKeKB7uKwC49xdTX+FC7eK8WAPJR4EwaeYbdyOZra5+ft6WFjpp+6CcG
1t/zfybJ6LJDGcv1gxvgKkAiTZnWfOe3iTSoVi3tF96w0mXYdc5Nple0GBQ+XUZVxmpZaRn6be5P
0r6Qes6grS2zaLFbyyOukyFiQV8JVPQiULWzZvxR/LTO5P87NPn9+Azjs+LLOQxtWLQ2VmsmWNYW
ZcQ4yulvd5ptcTDc3e34ZiGBq3KP38Df0uVqVCj9Y3sL4WqRsZbe5XFyJH5woMS6EYu6l7pQYIhx
z/b8kdEH3Zs+mw/C2J3XQImJix9a40zHGNLpvBCUTRQ8X3UvsroSzV16Xsx4ItCMfEaZV7APz6Jv
/1Pm3qA0CIJ2LTmYtn7BVh0cLqA/DY2qreBGaTbxybxa6c0PpZXpl/H9dFo2ZnIwB7U8X5Myh/7l
5dgrax4p8xn3FhJtNkg6J9jUU7CwyGaO9AOK8nYzV8N/ufAdzL3+Il+wDwfuJ1quUBhA8dgh3udm
OVWiAw/DyVxwRgnVQ8y71hcebJ5K5WO2di3HkXAPZ+CWRpmC//jMheIuUkwRDST2ofOOrppBJ0Zv
Cs3AfHgevm/Nxo8yROBxBA1dDTfWqaqDPR1/8TorOcD5RI2hVDu7oAXyCJO3icIIVsKgndTJ1cVA
bs8hdG48WM+tZzSPYx7h3bWB6nCjMaQX2/aYTt19P4jEiFTwT87fBsE4faVeQKhniYqFCL6IjxPu
Abrta9g3TQE1mXqjxNv6bIdXts99eLEOkoOxiCH6wRczehAfrtcPHqzT8loUBvQEV3whP1TJAYkw
fqTkYhWeASooItMUCEvKJr3Ktd8sXY8NFiIUhZI3hGWaNeL5jPr4D2MU5Hrtx5QtkrxYHoQB0rIh
nvTsyrnFXHefEooDte48q6J8/2JItWCxohKld9Q/YLuOcn5EMkbnH+U4MVkRqobHz4KGugbqS5As
p+u+bWcMTTdAy7NKOxEOZRzpmud4/UMWq8g44APNwMC5GxvUFK4TTri00Tvi18+HnIYJnX4dpdOJ
uKOrUzTyIyVfcKq5mgOk/uj6QtDBqx6uas2jhgaG97+bqzL25BbGQjVnea0Hr/OJhNPZ3Tpm7NVL
5qMF21FKBC5vc3VofaJANDGbrpixr34wtjCX1+77ceH5+zX1yafZW2d3xiZtGpVFxtG151OLxsfU
Bl4bhraKjaDcxCjASzICD4LUzLdt6HUZZCrZ/ChTpGdngdi8HAjVZMW/aiWVcs1H/e70gKiUMHfT
qvxQUI57tv93vw+esJSOagYHRZxK+Ila0wKYYCQMdn3mrdQe0qpWAqgqsLcSiKhpIUBW8er+UNZu
aI1DGGWmuAKNNDtnmoBvUqhM9bdhckugzYn1a1BKvZNG3FNmam6mjanuCDcq0JDLgdKLiJhHqjqU
+RChED93VFEnTC19db41RoCMjf4UbqC4HqwFQgSYleBvzYAAPfzZb0u6iu5q7a9CStOwSDXwrS8B
841bsuULbQJdQ6vp4UgtOvepd4uxaIhmlGz0KlDWDw+R/rM4o4uBu4O/Oc8zqpf0WKla+cuFWeRS
5ia4wLHdpVpD1pR22oosBN5DMShQMGafdf7TuI5bSM82tHaci055FPpC1YfgP9ivopuBSNM+t8Na
iqPveUcSr07vIXChyFxtNEw+bEV2nfzj12f2sukeSHuROoAlwDv8ByK9CrSzno+Rn8DIbLfOPcVR
TWxsWgjIDzbfxeZg5QfYTDIoJK4o7X6WEGC1Rh7GWml6XKT8koDCOSPb7TQA2vklEOnSkZgGwp1v
G1skmfUp++jeXPrFNSBbKgvWVXddtP6OhrLTA+PL9Tmxh+XTop8MpIn7hh/HmWQslUC2m7GsbbfB
oHrAEdGvWRLiVP3VBgg0UbwMrjaz6xyWmm94WWnHQFTLBXNAjRou5r+lcX1MtpSeq10ZDhuOHqz5
/6VSKxc8o7r+OABWBmpums+93l+rJlSPUTZxdp5WZMyznY95MgbETFpOSJEB78bQXQFN2T37umf9
43F3AhoxcL5OhsMg57vhPFSzd5nNNWILzFWEooM0ejg26BgHTuGybp2k9SwPOnC75KyShxAxwjQd
DR168usiIXKEIymVkn+2AWUTJSqeWxqe2CyE3aqrk39m9+ac+JRVpgyPc9IwNloUzzC2QwAUW0Jt
9AgoIyygcYK9CrXXSw1ipD/gN/NhHnGWBEPc2nW9Z7XkiFzO6G01xIfBueB3OQJjqG5TPqJX7D2n
hyhggZrlH83pEiD4t8sbGaXExm6zHhtl+j+0TLnfJswWtd0eqpfrrYJFKoITFlcc4apegTRqzcdX
Lt2YT44AUhz/X+yTVcFdB3wRBdr01bnv4x05wWAkAz9djYncKgzcmteZRxS/Xim9e7pmpVUn7NAL
ZSXWFEpq27/kutSFoGw5GFga9/6j2ift7kh3cQv2GeVUaZyCgd6va0rMBli/1NCkWkiXJB8ckKru
9UFWxOYgs+UtdsXoDUoFw0vvGpAL2nGKNH5jjkx/blgYrdsQJ68CtiT1aIc9R94NRJ2JjUhG3/aX
5Auc2G+n8P1GyIpZKaM9herTt4RbX8HfAPmaFpik2RlAy8Ez1YQFyMCukNGeDybZ64T/YdJv3tZH
cLeDrdByje9Rz6ul2NfQHYBnUFSkkLq8svYwsBgkbdwYwOUQSdUtbiiwTdBEjp+vtW6e0cM9LULY
jUd4sKF7KdauEbeGfpm6jnvVeY6dwxaPOVysdTS/o/FifawhKmBeAX/NqJoKXWwy9JHO1JQoPBaJ
ipi2QD4oLCRQ+OkQP41fZLry5uD5Pmhrsrf6r2gbpnH4B00ECf/Io3BcA/stwzmAOmo2YW0B1Nag
ApDMSbJxB4dKfACurqAmmrseK/LPp2xN8+QW/GhdpowAusHGdIZV2kWRjL4xrqnqoJ32O++r3zJs
Obai08u0UOpst7EFmTPfUACn+E2RHxRT1+G8dgU8SICHPlLblnj5L5muuK0G3LDsfESmEguB40uF
XkUmCSv4ybPJQMTPN27ePnJmGW9S0gEPHF8iEtxzx/kwfWSPO3Gb5ifrhh9BcR4OrEFIK8VfzUOZ
YMjTY/nx8gpEgbyuabtWHifEP/h4HPzZlyfiYcDSntaSbLQ6HbHE5mv6XTgxcI+wRAiBHY4mYjfx
pWdbdozV+s0ji61yrZWQCO1vWz6YJKE/rAj6IH0kAMR9LtdMhIdLRkqlGUU+lV4+O9YXI31aSxDS
+oNmPdG7hR20K2J04SB1rp4ZIZ3hSovHUh6jtUJEfzzvWw37FyHHdQDy4sIZsT8iQmKjWudARx7s
0zeQzo1cSdMeLD8zzaCNCTUkv7VFOv1JPfYZy8554uxSLzP+mWRSrLQPBJddMAMyPtfcYKbM7iSY
uInevAtzCySRrxJJsgij+4h/0rjlIrvLlypQc17bBMNHYqpNUjb0k4Ek8V2A9puvr9MHp+DruV45
e1qMhn4Cn9RrI6o0k3QBEwtjbg3LNoxmyzI9lH91gyuyhVIkAIZaGe1uZj6c0KugTayXy6RdOqQX
V5V5eOhZy1w5g27e75uvXb0PGqNV7pkfZEcFuWlq93I5Qlgn1FX6Ouc2zQubDOlIZp7TW5z8Zrh3
VZW7TLgp2X1HNVTmo5PhQkWAFWry7eajhiNCBuMgQnQslSNWQ/IcgQipLE9sT4gxbMOi99AzgkrZ
35zrP4hv6gkW+Okdb/o5BBKNzv54ofhpRf3mzWM7lokkSClr7Du92YiowwmaGe6mu+fGPzbc/auV
7Ucg4AYO5okZMjPD2GXHTU1ZZ0Y8Un2cwNzXCoVUfLFTzNIvTeP8vyORB7PGF5sMUwOZMbzDmZqJ
A35YdqQ74YR9oFFVgRwkbLO0QvfSuZDtNRqJPC6B61eOrhmM4wM8DSXjZUj9+5kOz5Xx3BlaFlN/
mKRWcNewHpuWxUI7yJTbCH4LvRMRt9KXTVAHkfES12ILFohEVoWHekfR/aszrtj4DIIxCwMtjtl5
/nkLAhbT7FX6bQrroKtjAI4F0A9f9N3cczfCBh2Ab73sAybd3tSjNx5d27ZWe2CuJB53aQtyxt2W
Ofyeh947Jt8ZXx8qrUSg6bnP+zcIxdCPSYI+l4Y89Abdzs7p0mOylMdsyuhn1CCdaao3/pPGnmeY
+ICOi0VYB54gssY0oXqUPpwyhrp21HE5A/NyOHfYUfu5QyCJ0+bTsiDA/8Su+VHqJXB7NPNSorgo
/taf9hjFn/mp2O5/PGTMIgxmIDEHDCHIUXFIMB6CM4ka97Vj+wOaW5rAUJU+nsWOFB73SZbs5tvd
QLYGKFD0KQXT9g/qjkBMRlJ5guA7NooCNYxv1QsTjv10y4LxFz/ueER+Q0Uj7Xf/DEz6+sy6elQY
VTNEqtalzKzrisX7x6lLqMwzcAiJ/vESznXREp95BJMm+6qTjv1eNkpPStF+6yyaW/nGZj/sbiQW
NBTursy9ScjsABLnaHP4ng9opCdHMrUx4lxUOIIzCfP3u/vcHrOgCOSckQgox5ZkH7LtllDboFtW
UZfzwjiPcBMTxpHtmVFmm1BYygrtXdq5/xG4jcKm0hyvCp/IjX4kbubx1vPnc/kT4405BFAjqGfa
5+W/+VamJm+8xcECbd/Wy4F4yd9+kUF8lUCVTg+y2IwdlIMT9/V33hLmmZVotXn58D3DzeKFsweu
9NfcE5xWUTNCa2Mn2C+H+dRSHhBBHp0QUebTwNs1ZYOQZJj/dIyLAtsFMkUO05gu2qKSG1O+46YG
s5E22C98aWZ73WZm73oUDO85ZXZBjm8E0oShoH5ds6SM5YTQOF6AXtO7g+3LivdIhrxqogDam50n
cNO+pgo51OTwyFYNcS19n2RQmorbTvRiWZKNK8jv8cFdJC7424AlZi/WqYQmKE9tyUWQTpSPNuGz
QxvYC8xwkrRU4j5l147uLcsVJLX5DVxo189f4fK6M3v1cJW4xHpxMutdP2umH5o1S1e2AJozvuum
9QtILfrXNO27CKgswuvfeIHtH/iAIybBlD7o7/GnVsrYBceBwYFYeEtcjCJKtamu/tqjwvSWZ53P
8cRpBZYlf5kcwkYv0RyBaHM10Vl4sKa3FwfbvCX49Qj5a/KQLRPZ3vGcfu0wagl9HDYycOlMef65
o5XTSXOV5m2t2IunJ9KLcRJuYpFNdtl1SZr0SzBxioQl4HhQ5YDq4EBasRLALygOH8mpzko2T4nY
J/9m4FpQ6jqApQDRCwluycFwt0sTAd/MQipVWYIdWucZ3KKsN/cT8JVvOussnkCumiffq//Qy1oH
lJrEV7GN7HAZdFsDUOeUv2LmA5sKjhKtGY50qIT2nWypqZakRDHQounJiZtJSotU13LCmSBSgYY1
WQfGemfWWzw56M4HAt/mt38AhwY16pfSAxa92vO7s7xxphvK8rdqobrxCq5KAoEK8nLLIRnrKNIH
UquJydiyjFO+2CT/9ugfu+MZEoCpgsaFSMvZZf7mBE9j5ycPDsUoxmvA0JKB4ips8T+GhTrwTgTi
Jvp2rHV17ubUUtA0mAETyVFsruMDCjXHPfn6dJoFnpz5nESPU7STgk/GU9abqsldbV2juAabKAzv
VkUl5sakcPXsygYclIH0+Uqb3BMTVyTO8ie4tC+QfMjbsxTVQctvufzku/Z2IQyeqmlmbvfiMxSn
bqtuVP5a9YBgfPOsNhGwI20Q5DOMtITZxfKekPSQvXQT6EMVE7b6p8eSvc5mwFTtMnoOdViaU4gu
7XF8R0S12p2fOcQd+qNYfgDQB5mHj1fvmDgWllbL1NrdbnQwsPmM5nVTThwJ6Mmtw2XkkRlBiOvj
slJ0ya9N2nLiQ2LSDnOOdxVwBos7jKhMtaj/RqsYuNx+zmcq1N9oM3qgpKUNqDoYkzz7gLgfaL/Q
+mCJjiM5B8fv/Y04E+dk0GMHMIQn3aIpeFivnsbG786Ax1CR9KS6DhVt4p2VgfKYeFit7gqkmHG/
45ToxDwliY9Mo+nK/YjItpbjS3QSqYxKXFYtN2oumUGAh0RPeXS2IDk/Iw8+tA/0eVG5jdHFwF1E
2uj3yAJBjcEhDBzo+bdCZqp+usxXoQ0tTzHxp/9tlCW5/JPs6EMBuCWjTvX4w1uvJZS0PmSQYAmb
yxJte5xvZLarzvmIaiZAxpwjx98eCVEwBgii/n16nDS9vmPPaJq/wpvC7rDBrjancjY2YLeEk3f2
uFHO2zOjfnQWkyAinjiIfZAnVLVybWYdcmV4i+3MZYQ1K9ytH3354/d+gOXELbLiLIu99c0GfKrm
7WWpiqDWzZlORha+uOTevKZJV509l0UrZFPCZutDBdX2YX1ysxG6aOo/e2IKKb/MtVXB1IDhmI0+
JwTNA9G/jzVl+z0kbUXh/Lo0vNwsdB7n/NARjWNxv7Tj22Gt9w2LOs4wp549+o0T2cTXFAlL844l
7eNBuMXT1AUTISIM6kXeGTIxwttPe3ywA9Q+uuRvhiFNCwzmLaP0HasOn2TRT2KRw9dLtdtVzh5P
DUIiHBullT3a4LIvFf9NsrGujG4uRAJg0oYI1akwYCCepTqvn83yXKdYv7l5tn6eGpm+rxiK/I5z
GWTZDR5e8DxFjSYiWsDsmU8OYIJ94+0z7ZA8+3ZbuGLK78gXcFoB2rYevT/eOdqqTpir4iONRtIA
1dVnO6cIsZFXOwX0ILyMqST3Akj6mij6HRykfLXXMSX5zwKzA7vHS+OL/TSdm7vUFrcE++lWCP4p
7QMLWixzdaz3HzlTthgNaUo82t11Ml50nyoLzF+UDE074RAfKRq7XV1fLlDPQ/k+OdqaBx3402RR
oYq+Z41NI3xxCROmxGqImGzg54TFQ5Kcp66R3gIJsPUC/I9JvvrgitmJlRzdJNZAkdXrvcgOAalg
T9ml58OBdlcgXJ4SloKp8WEH8wSblyDTslq0l5fbzYQrJAdgqGwX8fLORx//pUI9iBZgt10wJpRp
1Pqs8MftUhZb7N52blbM/LHZV7ATMGQpbxM101M7Xwx9ixT5dHJ2OrRDuPixQDhi5CWVduGfn16p
aJ/iICWPJVvHTDjajRiBMGB2nYtg6EbHa9wlLVJpPreI9BTPgrH+j1E7c+JNTWkx+Iu7L7Lo42kv
1ZC75viP5E3FU42kNWE8RaVa8bFqXUjwAU+OzcwDGPFXTbMcZ01UwHniqKc2PM/V4G8e4ICJKASP
SxW3Q/IEHDS7obyrOJOIkw6qSNp+TV+XJtLJT5k2Hnnjx3POWC81rDmysKtZ5O5y2E3Ze/IF3dE+
BIkqmE9By+uGUtDjd/ZcTsF3or3VLzjxpqUk4U5x8D90gCN1CIhosZxkSCW30nalDosYJnDuImCV
0vlQZC3rPc+IASqP0vdh7UW0A4G8brwNpgzklaWqQLDkcbRg0lznKeGWZHG30SvIEcOZDCTwDmqS
w3QkAL3WAf16KruKC+ECIgGobVro5cGbCcSH/XFaRHmBLYTnvvJEyya30PgFpJvcyUJdDryfNTPt
AE53f6LhnKNRU3zRSVYZqK8JATTYBagfFjo2B/xsCrfnFb9YZFNVXgLVEUDpx+/FQU0t2JiBI6TI
7V7NquytPAoGsLutxw+dW+sJtl3uUnnsFghW0KaxWX85FrXFX8IDnYI+nP6OO9kuQm2RJAPuHjEq
bmndIuP0VHYgrlgeXokm8+bCwCD+VDVth4pZFetbz4aRFBFQpI4C7cXq47P3IPVjKjeT8XjwbvuK
NotR3mnkiXLz4jv6ANAd0ovyOMM0Nz1PV+3z+jJN3giaiq4q1uSe0MO8VOXnLQ6SRNin+iK3RZPE
0IDuOuWSE+OQGVBLzeqgiaHXkZ8VRTPsn8Gx0zyE4wl4n/uSFa5y5nlE4nJUAMEKGXzFHqgWyJIy
0H167GBiLORli7A/zXn4kvC5b39l9OZ5XA61A+SbLQnElBuUpjV+VfyPza5vkynj7mCuFJqOTImZ
NPQN1q4NF8AGAZ5T1ZcdCw9ebVAWL4MPhKGHVHmBpA/pgSvaUh7HPeQgFPVBO5SALXuCz+a8Vv0r
JXFBTIGgYNZ0fFK40n/5FJTR7oViqU+cJUYyXscjoOTdDzakKoiSGY/tNff3xkKpZ2sDLwxYsY85
aaIW2ObQw5SPZruHL+ZeBSNmr4rbhFrKv5V9EJq8VNbjXhl4A9yq7uGrl/vXXrCO5vjA0L08NwUp
P0ywRNPZnxechHkmToCNWzdE4FvrU/y8a4UZ/uRPKiftIIhe1LqvkF6bzlZYmRu9Brr0tjMqNby/
4yVdUoh3StyUKmIQ5wuuI4H+HmiK5zbEbnPJSF16Q6RMoKGWseuLHzPFZor0JtlLrTGTMFlW56jx
zNtOvDSQ5omQm5l/032Z7jIdumDlnvwsQCC5zjBVAaNDmcH1ETASuHjz6b0Qy3v5c4+1l/24kMq5
/Hvv17UemZpp9OfznJR52G59rKgxFZWNcBayWUd+95Q3Uo8GRSeY4y3ptQ0bqUCkibLI6ZYFopxx
0QMvK7ko+DmlHYV42fzwMmYN9qjdgnIV5XLG45+URHWfEtXc8vOyEuhGmlcaTgMO/+vBQwPqw2OW
uy0MQCeMU54pT0jbq0wgXsSz7DWsIE7oJjltlWQnwNZ0AhLn2U+IfgsMg4OitJLl5FMkgQvvLR2P
1dFO4K5QzuQAxh5F78pD0YwjE6yajwmRp2amHCt8NJVFL+qHfGM6WrANjBVvNNXeBi0Tx9cpNSHe
6sglmlfNFDMST8jfewza00/CFBqvVQ0+YOLg75+M0N2Ff0LVgHgxUCJ0xcJyAmQofMI8XenB7yjb
ZUmHfWkehS94D+xS9Ifh7aNrFdo2IqgNnNciiNCY1AoTL454iJSucIXl3GaUKNWPF/ysA9yDlIt+
Ww/Z8z3LKoe2WEUDUNjwcNnYephTsrt46j/S3Ou+sfINhE4QQBjQ2pUv9sj+Yr6dhru8gVEqTwuA
lvRP1PlIm2RqDwRwhBDNJIKo+9NyIBuvIAJsKwMXyHwq2Rz5PjOXoIImnVlVgSGr6j7vIeoRL9Nd
oekBeAPxU9Ea/pAYwSWen7v6sy6Qsq39KZ1HuznhziArNeU8pe9NSc+a8acC4ZTTL0tYPIkavsG2
08KhucvPSMrWM1nBKZ1jOdmEIuiNFrL0bt5SWyo2v+q+CQAJqJmXhcJC0tqgYvjfISMlfzOYdkJu
f4xrtDcKo49daP2jRXX8fqmmrQxX08YtOT44eUQ/DcH73q5Wtn6ty3640xGHWifyLvrT9xWh37lJ
2j1dqVpqqIaTmUOwBvuHG9kWA69XarMxXuep97JJdzIOdW7s5whsv+mMG0BC3mz7ykT6yPfl186E
z0fEF26jyR6xYcdI2oagu0O504tRT8Hz+87wySVUHAwJ714tcwf+TGU2mER0AoNBum2BDxNMuIcZ
qPJsVYfQOhaAxoH9JapvRisG/QX97uEbrmPNkKzoveMgdeZtBssiLY00qsoBvb3+gBQSGiZag6N5
ixqOpiXP76qoeZBNx0DSWAih3U5K0A1QkOotPQPycONhJcieWKHywUjTeKa/iRCgMMBWH1GWGznr
yMXRD3KsGm4TSstg6xBBMgZYTM6w+QtLeh0VGiUVRjMr2AH8zGxalyKvd/5DevpeNT7dXKyieUG4
04anfxxGQC20WEjLWuvAz4eub9W9DUiyj8TWO8y3sXp/ZUWPr8OvTH2rh5c5RgxYv6CAgq4+NgIc
PUL8QaCwF51doR/3NjEQKyHjnqHkJx5n9U+MyZrcyMRDtQ1xZmSkwPqrgCkyUSbOpReW7doOXIeP
1ViwIBmCq30/5kvr3wRiOLTT8ZAtTxcqF9b+HOG9ay0DMq0Edqox/+GZ61aK5hM+kpjmifr/kz6L
snE2gSCtPqG1qHUsC2gjsc154C7oAzO7Fr6Jrm8vJrLSE9ngfj6PgFfApXe2907sn7ROC7rFsEP8
s/R873+B0bsKjKMkucKDvJNDsNHihQw2nDxySjaSmLX+wYqxoQ3CgaDY9dpsUJvXS52WSDqqN1Nm
57NxRGoMu0n7ILkGCFWy4W+O1IQ7SyM5v7cSitpi5G42ndYAbkS21F/41ISxxveY6w60V31jeRQX
kavBR2Rpm1GktWuGBGOt7WmKqLthREOZVMBE8vmr0Y5UDNPJKLS7xCsCeDbrKMy3uTcRGbeJuV1X
vBGiRhKYWnrXw+i+ZpHStZp3ipXFStR1oOqqNTrM6QY5PHSpkuS1+vlxrEmeEC525QCTjq50az2t
kDf/Gsd4MPaD39mR/NslQZJGIoI4a9XHbw7JqZysEcGtRGaXhEP4WqbnLKbTA97ohfwfF3lWo1oy
EXg4ZSYQJ3UunPy3yOaHTC+WjqRAX/vrdZAbqeB3UhJbv7F90gVtx3Fij271Ot9A4/JpngLpNtty
J64X2S4dEOuIq7sixc6uBwLD7oOkUeiL3OKJsmYQPmfH7ODEXfjTYhA/adhcVsJj6ihrYgL0glTW
mBI/RG9u9uyuin4OBojkIuatuGlY0VvWkKNDelu6luTtBxVJZpWUHp2eYDXvXJLWmXt1JtD50yUX
butFVxgS14yFm0qAr4JXGNQmXJF/cNwVQPKuiMyb+jG4eGL4Fu/7o5nTxu7/XLpUMM8V/UwMeBVr
++vwgiQAkky8/CMqYNzJZ9YF8TqNFf+kTtjPB5FHOOTddQwHbxubW/BXfhiBYcYrs0foql4pitN5
t3tynurvyOkJ/JeXfGFPW2wBb4obEuLFbmufi5VTxKKvGwWAG9V2eFgSOXf/b5v0vYb3SFHv5Z5Q
f+XjR7kzfUGZHLsx+ulrxtxmmoZrl0cV3xZygEw7Ko0fpuWxbCzBsUAa9nvHAjwgyKJ85QoiClkq
TuiVM3UuUEPpayebWlAv6jyxmEl2/kW21EOS99mQJQtlzZAnuKlV0OLgvPNITtHeFOEuQAF1XX/o
4OM8eISftl0t3iEQ9Q8YqmrTfPhJulu76ESGUc4zfrsfBBYAIXIXF5bBI8ph4RqhwdU50cYTyXL6
oHAOd5NJdWIhFfCPtHE6leSmcAyaexqk4zeDvg7damf4FMH/6z6NhFvNh6mAk7f4GY7oD3hwkTrY
CgsjTfRIbzkh5HnxezXNzJxZc3iJXaa+wjFnm2ysh3Yb8L/afsGAz7P+mW4us7yS+yNoRG3JECqj
y2Dt+xw7ljubjdd7N5514hn7+GLy1KZ2y3nWsKGCnhxhtxV+8s4XT0xNSUekufMaC6EK/wrLi5hO
9GUqe5P9aP1+4TQ5GX7roVmcRNP22lcuwzn16z9OWXGbCbeZbZKhZypbfwdygS1cLlM0Fem7H8em
ucTOH9/LbcOpxKDkJDssXmulBEVg2QULmoQEmicO4cnOWlkADcDtZ0ci5MeYvUbx7aqNZb9n4cvS
oYeM+J3Hz9Gpt1AiLNjC3ITszED4E298itJFVqHz4U+m3mDz0BXaPNHA4m4KmaG3A9QOYcevHtSW
5COHO8nTJsH0TpsG6lzHyFkkFVIOLGtyfRGJJVX8vZYAFaFsOiSXyHvE0jY2YMnjlKw3LWpumexA
rd8ounGcqd6CzHEp+zqktYBK6CX9f+iiNkA3tgGlNnEN8hdGn4+dOnK1A3EQ3lK3cf+WmpOU02jm
naBNlTneO5ZJVM5+8CLYP1ha4z8vCKciNbPmmwip9RwxT+RklfksJ4+cQ2ytjHwliEzrO6qGPcur
g8z2FeBOU92IgYxVFKZq1/tZcTNBNF8rV7x90h2U8vrLNwizX5aLzJy7UrVeaqdcgRmPgFcY3+eB
UA7u5fmQqUxBQrZwWCKyWuOT1YwGl9zHL4akVDgsjvSplXvfUxoWCLqTARHTD1dU+X75bIIVGeOd
JjA8I4s6voMHCZE/0BXGLPLz4SLp/gngEL5zfYVE0z0epal3oEk8U043WltjvRPxknWzOL5D+jpr
WAzGGS+p5/oeSVa9vXNkr0G8feuC9v5johjDdNzYSeIGGSia2V4HGjWtulHz87WDNfZMdgb0dc0G
3g9gTk2t7PDnU21V5ohNLhtHNREp+yBl7EeFPg48Gaswi1n8HqZbtA9qyPYN96rBdVCHkc+n50Vy
98LfREQlK4G3yR20JxP9UYGY/nrX0z8TJM0bYgAmkzb1GuIDRP6LZonSEkPNV1BhxBFbpnGcJF6v
LHa7ISa2QN3rmCw6MpjwKcyYTiK7yqz7BHqlzM8Mj0f+F/i8Ku6jYjjOVPs+v5Y1+WoyeqrDl2LA
v1aBRd5h5n2HDsGj7TT40i2fFDoQCxhLiQVNy1Fi8g0qVdEG3MSsyq6MbYuYjxpb8aa7LKR3FvtZ
JVEvWV1CEs7peIb1FF9qNCpxAZJdTINRxeyFpL/zFe19QoR+nqkY71AWINs3uBGCSeF0kbLBDA9q
gLoof8Bo/zAYRlDNvNTr479/Ti21tgQatlI/ejhlrWk7w21fJG7HZ5IkIu8aorLAi1Z9fb/5hryw
cn9bd5np4m2Xbks+Sc4HmBxtLN0sSIB8IO9VWJFZGS2+Vok1cFVYGypqcL9PfaPgzN3WJovs6tUL
/Mq/vEvoH/yUuSdDmOuaIaP8l/ZnfE9+z05SntDsqnebDHWg4+BULDcofw5Z2cVtdfzomuD98cPV
xRq5qwGpmewHjJgmCjahniMTKB8mIdqMN6UKD/KJf2JKX0OEkn95iM/mjLvTrUpTrJkynznxVrPF
/BEzUwhIHspNnDgheUSySUZYh0s1Ze2tVfAkvkKRMnxv5Ow3g1e5Vhp1pTqmOMFHfbmX4KR6USBm
BCyLNJjNlZ999iK92Gpymk5Zznf8NjJ+GgzccYf6bAQA9znaTjD6xiwS90o88/sdirGgJL2johP1
lsQ67AIt4tuY8bmnmhvtz1Ix2BF4vTJR5oLgzOhP5mQZx1hq4yQryrdDnvyRM4q5yj309JRXD4ck
d7JGoNbuNE++RVLTmdDhaSp5NOaqGF5Dacn3SD56zpLy94BTttjl0vvC8tJSKrUIFfLyS0x3apuA
Mmb23l98e8LrMnmQ7fXA/rdF5DYATT8LMu8qQBFEa4XadXXIvJR62mOte0E8izkdSyHDJbraROSt
LGKNn/n3J/GArBeyW/QGI5KI5oS5ROA0tE1hCemn/kGj+xVg0a8q5uVtekYS8AzEP91A3mzSHMgL
Z1t8L0d0ORaZ+9ldTdzK75RbQlSgB3i/PIl3tNqMK79On+UayYsPdaiztjgj6w9wqLmwka4dt7+1
HoANfoFvvlZMaEymG2VEgqS47/iCX8Jgd+Y9SI1HRmJ4IKn/P40J/LykNJX+mYV1EO7nZMqEwd3X
IqMn0OiFIb90FOQnQFgy4BBB7ssLiAXDl9hXWizdwHmbvJMHBkg+Io27B6OpbUMXLb7mCN9ivCcZ
C2bQkvlLSmVBW5yocEKH2qRaN5ClvF1bPTo8My8o+tLSoiL8c2QUEbtx2W1xQlnEoL0awglWXuEi
TIdih7XhTZ5fSXwZtQVNydTadB/pLvDlVAfP5Pfaryt3uTdh0VDjTEjtpLPkXY7YBW6eBjHUoraD
8P+B56VPuixQUzyhYHwYtpNJ8XIXJPqvt8tulbt5PxuFSPmbJEQ1tw++KykCp5L14FvGIZhtc/GN
REukkXQEQSwRWqd0hkbyqGYUID9eKV7+a5hEEs065KBC0sE5OueyKtH4ev0vSuTq/qOPD5/fplvv
c0IQaoj8+lgy6ai+4jQXY3xoUTWPpHIMmluAPpZ4zJ+jKNfvaNAF3hQBCcp6pwhf95ho8w3yJmP3
eYqNSvTCMyrwERCSbfZZrO8HMH2Z45KVXov2did771x66jNT2YvHqKX0uDXNM4et9YgzYC7RWqMX
CgnDIxFbnYis2ofLa2RwwMP1HlZGfKVBkN00ZUHZT+ZxwCv0eZ+asHFHiQdL8eSzpXnooK/uvT5n
X25wPaVCrtPfgka8iEvkNhSszhHtqWt7Hb4iR+ZXP1Ry2T0sV6tHehO1ya4jc651cUR6U9vGmuSd
Nhp/rG3kgIjIef7HM1J471EYYoUDVrSHCz+skrRTW4vznfgcUF1aw2kRjFc90NFD9XhporpePEZ6
n0aoP6rtzO3Ry0pwoi2KfcqU4D/pgXaiWuABIHncVAEA4F/MY246SBB6E40xsgLNXCyEce3MTrcx
XdXfnAiERBtCYxmKpfAl2Z8uM3NEEb0gBhG0cLouyL4WCcHtB9JauRHyGQUIXepDAY4fHe68ur2j
5itbSZh8On9oPsuoPTxlo+iPOguEIUnpkzeNOu/Ktm0zJEFU9Xh4pladB9q7NkUZZNPjVsq5Ew6U
iweIMOht3LeDN9O+pW/+pTlKmGgs8QdDO0Kx7nToH1Tz7H+aeIDISlxC+PTjAqFYmLIfV7Sa4bQt
4jH39uWqK2SNgP2cf0AAu0wm/3/9HLx2C3GtXUUNjZGjIXI051qU9uyxqj+46dr/cIf+2RACO34f
nP6fJ0RniNClGHUNStlax0eCZ5M2LCNorATqlioJqIpB/BLjpNP0Khvi8V+v66djvffEKjyjAQ6/
CYIImr3Pmcb78TFmitklwBzca1+MTb9lkYnla1Z/Q9/uthINKeEjEXgJHXRLMJWRh9eToC2MSkUt
lmhbST3BKOc1n3VjKc9i/hmkANnvEfQXtEDGExrZnmJ9KAmqXDGpo7Wu2Tgn2YkMlFNFYpaQirLB
HRouG0RAUxg3M1ma9eX+ef72UQqSHysh84KmC6u+/5jE94352mI9Lxl19BKqtUraWpd+ddnXc5a8
a826KKXiINDBAJZdVxpMvFMpJ5XdNK6336+oBc5UimDAvjGxkWG7OIZy05lvonAKc0t655TMFeh2
T+UZk01EIhHh0BsmyYFiw0LVRjSK5HNKkKWv5PhlTXwWSI3vV+InqxrT2hUK/IVrp880vVQ/QbL8
qELuLov8wJjOnNlpNKJ25G7EE9tibzq9nnDTlGjmrODgJAhgV2IA0f2jlYxKvZsnu4RDsBnBVTjb
m3qBN7r3tx602pODajHuyCz5JsOYWyY5xr0NP8CVnX4UBdd2DN+k7VAIOBmrWDNshPkN1CGoXskv
c7xGQobcvgnqidhEipPsar4alVHmqzqpckPubJzMsFmSPobb+6TJ+jBqQtc3kk6em8kSCu7e0Qd+
9rJPxksmC4mtID6LAtcU8GioxpT0LtrfsTkvWKuCMIvj4xL8ozp1o0xfRckmHGwVxWSZJT67+OWL
4biOarN84tlDD4p6vwtur6UUI82RRMZubA8nzpzTzm7ebxey9a3PApVItcd8ztr1BwWcky4Vk3/+
8i9Dlxyp/j0t7DcFvESShwbU3gZQh707yFnFAMKafGT29MqpO5NIIVrRbUtQ3M2wRTfx9iW9RK2c
rT09IJ4JhU8DuvvYSkLan+WpsWfkv5n6CdWMfUI/hoBMsTCj2W+DiQuzr6XRbL5HjMW8A9byljS+
oK4ADoqlHKgdYhu59UjRMcR9BGwouQNHdRcbyZZZvHhN+DJxxz2/HTnm9AhZL2lIfXmPzRbndiaX
qW53hCc3iG8PrrB5ZwV7hD3orWg76rW+qX9FhuWjsashMxCFdU+rFnevsDamO7HY+x0R1SLPXMR9
NRo0bVA3NXWONdE/QaJVdkbJgR1wKKB/daSBJD1aqE5lj6xqz+zu3rm9Lb8flK6C2UQW13HPDVt3
h5RF99siqy7g5KDFVLNPFQ91mM9ETGGRf5lgApzf7LLFbofSQyRa7DlVXVjYcE3/Y0GADp07uYmG
7K983qewv5CyTX5mMtu+UQPQ3Y3CI5akLi7tOGWidlkbucLiv75gm/XcANPAOk+nlDNKHpNKRSKB
UoVbsmm5jz2nIai5qqu7AOeKJlJ/uZI9DBnuWXoFvWSE+7CLPEMzSyI4QUVBywrbbhWgpXwX9UnK
6ExL8I3c0cK+Q0qdpKThS+lGJPqP9hXQv0ufP+RPOBR68tFlLVZvlqXe/Q0alQcs6Nim2+H60Zra
ggq+EZoGmr7RqvB5BB488FaadTgXT2lT4AatGnVKWhhi33YosSPHfuCCUH7jsPTnGosH1zHK5bBU
6D4VA+7a+j1C38ki95c42Bzq3ry+6A5Gve3U5Lj52XZsFu/usU539txfXxHT+EfC/xi8O5Plqs3f
T1ZpTaoTpACRT+cBEy6Ve9ZkRgdFRQLV+v+bMWA2mvaQWP8/ZWGrkFNNEy9V7u+f4FWVyAbg5mf5
SHrmqcFwM5eU6sAsvvTUc4uLKX2ykCQAtqE9kVOd3tjW1sjZR5z5MJ1WgEp03L2AjQwXmxNpTs0M
XpJhnLPNqGaMX8n7l0xm4hgw5JvVxbeORu+fpFHFa8NHCA4xG1P+NvM0gGex1TEYn3QCe1Psht+Y
ScG577PpTkw0RSOLA/Dclt92YGJA6NU3m3EzLZrc4vbt7c7k3sXOq/4E+Sj4eiJhN6vEIYzBnduy
xPYCEe053bbcqrPOYR60nBVNPHcAVNb3DlYong6CD3tEIih6Ve9/8si/ti7TL3wW8JasG9hW6ICD
x8h1+K4wDB2GlrcF28XikhboTEztonISLaJR2rRxyfhZf1OUzRE8oybg5WNL0chlZkCALUR2u085
s5auwSRFZyQpQhjVRHDfBJgFxQh6mxyLyZbo2EJztFEnGsBbqdH8lAz1FYgqSo37gmlxf+hqT3XV
JnQ5ICe209wWca+DcGP1TGiZFgvkKSijmKJtgBB794OYkGxs2OPIR8r1JzC78+88tAa/uhKpuPwe
7aN1fvj0rw1nJglgnAVS12Sg0iafpsXeULHZCFvbrtJi/XgL66RmXEyqQ27yaAOf+RkevMJ4szeU
fFzAFh6s3lVdW2DkwkYiE1rgUUL8PcnfokbK6nzMYwcbe2DGAYCR1poQ5H7Bi/HinIndV89yaxVy
fzQEH1D4hSl0Mh2G3HWg+p0MnG8CA95qCObDb7eekUW2G4J7VgkPKAThFjkR38lXRrDpXMYuqpAD
LlhsZ6oN8U8/m1X8nItLYs/MKC1kOJ7sQBuxpAceLMJBOuBP9XhlhcEzOa+za/2AyjD3PCuxn/4z
CO92apeimcOGpuNZgbaEtMM56RmZ7q1EfJgMqAsVgk3Qg2lDPH7/txI+x1C5HIZ0lbZa982lqaCr
hPw6DLQJooZVqC1yfwgqNeBhwX0WF3L0rebN8FfdenLwXMlg5n4Pb6MB0FlOjE45hMPaJq16ke1s
9vzeRwvQmBYdAgNuisQyodsVTcz9TPWLJxWv7Do36SjuF/uHkIIRoLdXG6l7Nn4K1GXSZlLk7X39
ru51buNmFMDIuriaV2VtiiifCXMgley03gVudUyCd5WznGusFKfdxwoJWJW3lwpNLML7a1IzM55T
MVd2vNyHz7Ys4USyxF9zPkMybytG8j1coeQJh2FefIkkFWx90779YFDYv7YsSJSer1r4gV1QOKbZ
ns2U9wmjtFTlz3wRrAIZBLdl7HxENcAxWjBrrxkwE/UXgSjZRj3RA4xiF8opT0bdHcLPxktvghNE
AuPC2KsXwAkt1rgdX4Gjoobd7HCMVsm6y65rdfo63di2U1nmOuhEGsdHsefFm4irOHxsAx/31hwS
j5PJ80e/3bUHQaLhepNDEQVqRUzZbLXTYdQFq5EM63CTzaIJ9zIMobrIUM4If29/m3mnDuTexFLS
8VnBxJmDqQCozCTMg8N078D6j/kAWPs/lP//0rL22SQUh0tlOJe9HMjN+MThlLDyVPPQQPf46yxR
lnwn9dFxGdNRxPwdYdwAxe4klLdq8tnINfQAfzKSJgguHEQb3jAi6x9p2FGUs6yg3k8AFQdc7jEw
r+RPjtQefHR9CCNPdPdmC8FZ94SmZR59/IrKkBrPPjC3PGiKkoDfbosA1JZJfKcv7vLFG6eOXfA8
excqwWsR8KdgEHJIJY8J7txlI32VW5yWhVE9FB60aLWINFlCqsuSS0HazDJyZPfQS35zheADd7pv
R0AUVMTIJW+4dnS4JEZWThH8OTOOH8hE4m+9Sj83lV+Gh63yLb+ESv4y2WWivCJyL5nYP/DUWs6s
u85Ugbj9ykMqFEV9IBShgRMdXJBtx2P0wQphFZNFWzWdFruxIC4lWmbZl50SUbvpeEPDpyagPS72
X3RdYukF3WinXJ1Ve9Fd1haTcHlG0hw4NFkQ5dFfg3m/A27zjv6RBZckzhSX2xIIvZsnuOKwrZBl
HdWMP7yfy5Qqx7MdvZqN0MHlekI6lQMGw4PZxWhBR7ropyaCHzHGjqAj+VnwPynsEFk2jalQdMKD
zF3ZMwokliDR8bVP5ahCd0mJQq+2T8DZbRn76RYE1zP2msg/J8/QD98qYGV5wMRgJ90iDfV+uhT2
g0+oFNv5FEfTAMd9uyLmaMpUxy2B3v90lJBrunRd6O7TC6ccjFnQ5WBxXv8wYD5ymyrgPeZxATtF
T6uLtVajCwHnkOarKQ4jWVhyxhJGIpv8ZRb4up/NApHMFpY1+x4evOBOg4eOKpmLldC88mGKqHTu
nSkbznAKeWzZTq009kktqIoXlm0e+W3bELXj/3FL85qgOtripYwY7vbgohSM37I5OBSsKkA3t47b
vskv2e3sYUKKmAM/cwcvsVaKyXtbzMCBc05RL3jNlXthJugkYJxi+3ggsuV0ZyqNTs1iJvLBgV3t
4nTt1HMnWwvJq8U/O59uveTPYE/7Habkc/fZ5lyCIloF1qJcYCCbjeiSFkOspmO7tAElXIFjYeFL
SYPZy6L/82vhww4c1FH++ZDxFLi7nEaNG2poMMNsIC5Gj77buMYMAMA4piAThR8WGPyA+0jBNqqo
AHnVu8xSzYvE9Gn1OpqR+mKIDkHP9+lLL1F9iPIWV/IJohc3DGVNzwQlF+WgvcklHN9P08ctVbcB
ZUP2rIHTS3jTqsvLUIcJ6owPsyq7iEvwrw/XAFFc3Lx3a9RvX9hp2yUiKlCar6+FWDy8YFmMaFMV
Q17cAGNtAUBiAUUaK+bnJPBxHi7DAxaP4RLlDF/KYTlPkHOmJLgQz2Wj0oqciMDpVkDZIhBGI4tU
zagCvRAO6RD3tsDll5ch1/z1n6xpfyaLImXBNc3QwdmCoUIQtitDBzQDGBmdVNgj3nC3PLEfrDGl
8ShZVpk0YzQbPfxkidtXUpaoLPptqJD004yjpHqEKRce5l84idJ7q/Au27CZP5zk+GWozkxdq0XW
A2fhH7BhhBLyfXkS3zN5HzTVW1LXat1xo30SltDY64U3j8SRnoPkcNSM1XpxGoApZ51w9M25RGJU
K+Balg3IncARtoV4emhv9GIVb1jsBcToZDe5/1gHluNncfaFRitfEugAuD+jg4UpAg6cYtCpdYra
IYOXyEktKgvNhlSSwwDnqCdqu9fM1djiUIto6tXPSaOJO6V+SaOJjrEw8H/GrFOoxQGtI7NuUrQh
4IKItgi4fqSNAFw7zWMt5UsntqnTEecMmCQxjEuzF3+bjvy0iJdoNHbBoKO2vBuFVq+pS0QMuhhj
5d3NWfJvd3AnOr3AFfXnGZ06ljG8T5fvG1GQzwV8nVcoSnnDxor3I+XtEr876HsGSozw8PeLa6jJ
WjadNeFFaLbhHszu3mg9kQMTAjPKblLrmq+o3CvvzHqFm59TnXdtcWrefec7DRJQOTyTu1jHKfA1
EodkSW2YH3qKJxtPPbRmo7j7jePPOv8FTQfwMqGXVKc/RrEJjivW8DuOYhnEs/lFxNs5FGZsDE39
U2tv19LZpS8A38g2u0EjzqmcSJKOFsrxChFJJvrkbUnxXiI9oRRJ6OGOT3FMVmuNYX0ojE+i5sB7
42VrlsEYenreMTYZlD/2TycAYANJZJztrNHBcNhcZ0G275RN6exSTQNbuwMG1GeY3+WKgjr8UiaA
h2nIo4bAWs86/DttoPUraKY1OYAuNqJvb7sjG8EnkufmvvSXbS1mr1HhTK1HJHA6LwwjU+zKezKx
zAsikqhg3eOXA+3nnoPFyKyoEJ0H1wt2JzEky/8P4x/U1V1RptORuwfEC55q6oWShWv2W1NKN7tG
pwMQZ/9f2+mTMrNZWDCWEhT5L4Y0zci4Tj3AluAy/tQxngeSENVSGFAdXOpiVUWSKGFYaY4hNoJu
T/T2CNgo8QVSNeN+E9D7mRsFE/SgoHyYqon/y7JldczchlL2ADncC5lfpfelyIfQBoXkwdIvkLGz
Rj2bFMIgV9My/6HeErjhu7H/q0ppxVJnlvjCSXEPNEXTcjPOwmHCsXiNGy5BF3P5FIAuRPKc0aqU
Fg/IL+gupYfvQk6ezR7/ye3l4GOXD+XopiuH40LJPaukZtnJW+qQKi70aqXLd/9z7fJRK4ogXW/i
wen6HkVyImvOZcFJedI9jqt/1raqr97LaPwo1LofvkqJsktBT1AAq3ojLRie1rDsE+JzZ6u+1AzE
zbYP0zaalNkYkcjYCNZ1NBSs2KSIu2KyNQ4lfC0RGJhaAeR4iQtmVEk443SaGbbMvAkAtH9HDqrZ
TJpmxwisQOlF+7QMst4AB9RFMjYFhmDAdRpooL/lQdo1NBIqhXBHGCLlAl0/AAbff9JVa5R3/Nh8
2K31fGioIrANc7t6rin+V0EW9lsvbdG56As/0XPC7XFs1nprbOt+x2sE52K7tQ3GmeT6vdSkc4WP
sZAwkG2ClIA8/+j+GVcq2gxlZK6kQ06bqxv7Ms4BO82zt+8eSI6OAysnUVJbJXdo1kFDzNuKG8FW
vkWUuN78J4CqbjPCsVhXiFqfCSvS3wb+1uPUhVtpRHDcmDcAEXdSXfcDwp9Sv6nkZ+IYKx7ii67M
9VC3EeG9dzpDBEosPONa7ukmkbtpYNR2gnKhNOTMHEJmSz39YFz6fkpdOqHgSEQaASQCTrwYdhJv
wxNB0OtTCsoX06QSKHU0KPCi7TT6WczFvO1GvR7BYBTHC1qj6zc8w1Wamk2aSOHrD+m3CSQA6xZ3
J0Z+vpNWGvijBAmZMkbx+s/46dSbk8ljWOB8XHn7YtMFXq1CcTzHfE+fvzIY0Rs+1Ewa21YHlJGw
y8dPkZxJnwOUQ0r4/4zBDyk7iMd6Y6SDLSbZug7YlWaosnqw2eGXwDz4WNiEWnqjvtsO+LMC16Bo
QLTxt2ZM4T328SLaLbcH/8m8d/CmGS1xVxWCeHL5pXUcii0eXZICg/309LxgflI/pCwrd/DVbxga
oGk6t6Rsi14xlIdfEy463rUzMgHMum8gpcU6suB2KF7iBKib/+gO+qsV2621tTxNyL+PATycJQgm
xTkiWbk4E6zarFxAEetrKqm1uObsGwECK6VcJGJU2c620jps33R9sXuTtaiBj9kvCIHXeyson+DX
bbq1dqMBNvZBbIHjRw8Yn7Ntva/haPDMrGnMGYBbMQnnU/GSgJVTQqG2jr+ToUNdqMGpGyltFicF
LULIQ8nt89FvuJGiX3nR5x+N8yjZgA3WoP3PEiVAMvKGrWxGtMuuXDRFjlIqD7v2aiLFQTFbQgbs
nIdqQxR3uwA1qNDlHD94tUbkZHYWvuztCxrte7G3k7I5T9B1b78HqWIipUxxqBiqvCDJ4EGZSvus
53TlQTgoilvdfHLkfgm0JddI4+l9cygQQt3QNPPwLf2JOFZBqrxvYslx4ChbpLL7WM9ooeaOUDRc
qOyRNJkq3RarqDndST74FElzroA8Sy44Z1v54Vkyzov68DjCWMdzoGm/pL6pJwCfUgH2Z9IVUbMq
RZcnZe2uSi51QRp+F7NxwaNuWGqhMlN3L04jXS5mCyuFNdY8Dw45utVOS+2bLPIzBkJd1Ayue8pS
oKngC4fQ79GQ8pqFsXxXSm3Pg6eYrVnX2WumLiypPWsN/jk1DqSDjRChvXn1D5NLf4yCPg86LGAW
12/MQuiwRxUtbG/QhG1xnDZXnOvUMl2bNssvVNh17/Lw8swRc8jj2TlrAXiU+8tR0kIYjdT+DROr
daprgdgTribk5xPoCC3e7xp/aA3U2AazGBkqWhfPm5KPSA5zywBitbYnoKy6fQvxShJMgfoP2AD1
21HYXZm0T2DuNZUKsSZOgJKwGrlPlsAoM40dLrNa30VF/y0wDiNKsK+cryHaNCeBZGEtZOBDwEuB
CIoDR3nAmU81ap5gosg7booklma1QsbIH00abzFZcZ0io3Cg4fa4tpxFAb5WOV9Avl60O22HTQIn
LeTeZQ4D3Z54K0AQNsTrZhq37hxADFj1cnAApBuUA0kQmgt8YQxSqzymlU49cmZMfJ/ceeEONq4I
VXl6GjvyDg4z5evWCbcCdBirV7MJ1UPLVRvBOk6bJw7ylpMSWWcGHnsxhsqTI4J7cFhcZQ3ARakD
0z4W8j54PugL6c29m7z/zXDM6e5jyRS+4Sux2N2U4dRB9vlWicodC3aWAtvYA6GWOGRJH59QtbLW
jLVCujikp5oWKcfLUhIAUxFO89F58UnFMZMSFB+rGmu4jzy3ogd8/+PTjk+QGYAsX5FnwqC2OdFd
Bc6Cg8t/cjLtisleYVnzzrjSA6JARuFp76YZZR6YmzPOY2jxn7bgwMrkZmClxZnMflOLWUTjYZIY
MPrlH0m+EEIQy4AbvDkRDcJDfeilkyqvwl3IwqsyVwlD95ACDrhq3TBbXuRG8LgNOu9qzxvXNKfh
FIzLXM3Eq/CMM+gAY+lZKHIZR7y0oLBryvY9MF+zBeWM5W/D9qBGTMmXvV2ldWWNhjrx/1Fbdmul
YMyc90wtx3Io2ObPTuddEhavFl13wmnzMbbV+ZzRkmGBx9eqMTTNG6j22uEC+hwj4ozfHQ/E17tg
Jl0u+LmlJ25+oooL0nBjYod0L3Xk4Y7OJAlNr0RDk253tVwbRrH3hhJabeFiERiYs/NJn7gt9KNm
YcGlayaQY6SPhvvpGk5lkavFmLZFfr34MFSxDEAqu5Og+kwPWRAbnqEnPBSBcy+wbEwOqFtO2dfD
8J168a7+oztalBL4jhteV/C0ykFFrqQabeyIoXZc5vDsuXWV0lJ/ovWo3+AOEMWFkbLqQW7iLW/d
D4Hykdg3xSX+9sLocaafKCSq3Zwq0bQyqpn+syaGzpFQ8mvu81hUk/ViIsV55jOp7uipqk4zeRT0
zAgww9yeBMbXa5CiyZCA+yx1vC4mDUg5CXHY2JyJlB/azOHNVHGKoBZpU49V0PtK3fhKCVp0tSET
lS6rVEkSGW3sVawgc2mjFrBpr5eLsqibtCXJMBQEfeQvunI+vdV9rgZNmFSfGmAzwCB8izI94Hah
+HtxXCNfvY9DCcTf7JuNYlV2lAJE6xLgaxUzwcITLfTgDab1uWdkYt4BRN9dPeBDD6rYemauTYR2
Vu9bHa1HGHSyxHB1XNr1CYq6B7Dj71+ehSJMMY+925SnkzHwjEj/uolYcJdALdwowlyehS+wQkGD
r6EAEBJX8qj6GiGAuopWoKXq3ZE0bQA1KwanTcKPEwWr2AiqcygffNEFOO+rk7ezyR6GOaeBh8TY
bFlX7onDqL5mU1WR+dHDD+FJetFeJtypNdHACX7vPjnQ9HjncNRKVZ0ZllxPdTC/ZUngd3mcqE3s
Gk2BL8JbNPSU4mzxLP5wIEvuC36xBkKBGgLcxk2z7+haDHuvy/50xtUET3sMGKucFJ6xMxMFXvlT
Oq+KnfTwOMiRtGUWv/hOJzCaCnNCvnxUnQiXJhwQhttuW2yIEXEpkbK4WiysFxWdnYsyuP19VomA
jo8bQSdPeskwjmwmzt/CppUXe9IUZS7ZeStbqyb3q7+JtAy+uSJTRRq10VecRtGzACpRD0wVdXu2
FvAK2TWVDHRUmdJMWLD0r5KJFdzPmcAm9QszkF4gFgfne5rvNV3T2KJaGXaShxC9wdd1dY87bWDC
ue/JYDoZJk7U1tLBnLySyvjPvbp54gEGvTgi+nMJWC5TsnSJoY5ebfUxqADBt8BHIu24iSyKEdZn
Y3jDncT4SLcyoOP2h/xNDwzpsR4Pyl0M2GmWLQ5bj+dyZNh+5LeQQ/YDeP4MMRHSr8Hq2pvYGSq9
sn74ubOmZsEXLbpGCyZkRgskiBTuwoVgFlJ4TTNjxlZ9qMyD9b5bcvo9r50uxJsQv2G1OMdySMrl
2VxcvfvQaek7hHcfMhnKYyPIZm0RtoO61e2xuqvQu2/jlUVCE6kyIkOG2rQ8lkQvLDI/m+aDi6Ux
iQnO2bxMXNtnJQqCxDoyAgsuUu/1XjqNqiibwocW1ghXTc3+Ic3U04KhAasZCHKp4/52O4P/MBoi
GdjcBr39p+m4eceoyDMXn1vz557PuXYn/ujle0/NQpIu4Xryh/mHFRKloPdlZXY4iWIg2csZU7Zv
CnWvbqPe/Sy87zTm5WsqaO2XYu0kA3Hasmbb1wIt4HLIVIOfUABz6pjD8hmspuod8QuXIlSCVj4/
mOxcAt9DB/4nTfp82rKt4J7phxdxvXcMh8iiEd+Z6Mq7aUN34IVBA6NzK3h/vrFwvNhUIEjjaU3Q
AOnaqYrfmeVjti8E41vFD5eSE797VDRt0Em3gRPakGLzuoEUtMzUYp+SumFwfrMtSDjNoR96BmkR
h8XRd5dmgvPZEjic9JMkTbLEj5KytgPulgzWAaqSnHIkifUkyygpgQjVcva/DtrCaAstxMdrsn2w
wDAttL/+MfomvWZMgABY2owkr7YOHHgxEtt54G3ERSIEDwJfqrQHNJkQZIeNQujej0iO2WXElY4Z
OYAdwj32n7MubWdI7dsuP0b4BI+rBH0NobI1H9xDYp++pfu72C96E1rGp18KAPbLcMQTRoymi+ij
nmseD/xsoVpIjAuGCSkfFRB8YmaC9NaLaqCA/71Ou6BLLPaC0vStxQmIjNK3S+KNaIsXR39Sxh+E
jrqDQmEh8Qc8ag/arQkdRtRU9b2yTwX46im10PqphPHDzsFUye07D7GX4ucRAJa6R3fw4B5K9NjS
ANNfucf26Bh7bZOsycieHHPOp80F2mq90G9/XrkewLgluHfW9/JR41uVeCwD/spjn7x9Xb00Tv3m
m4o0SbKKQLylRMq9dcOo5BGDeQdcvglTFbSOtFpwL7CTPHwYC8rmvMv2JWlCQNJW5nI/sX2H6oqF
4p+FCuaqpCPysahzrqDUzWywBihiBgWKE44I0xYKOVZmY605B43/TDZk7WEvoPTevc9f8cjTSwM+
V4Fb3TT4bdqptMqLDHRf97zG7Uo++poqI7whsl0JU7aWTpITnJdTjQj1DCktLgW9Zsv+EClUbwN3
/tlWpQLUX4yXpPjOVFH5PhTzjZQW4wrwod/xaM85e7gBAi5npu57ShE+fARZNAmB328Tbset7Pb8
1dA7Sby0UixNh7sPTRp1u0NWbjJs0OS7tpG9f1mWoiulesNFFGUCrv+NVfOGyJhFY3TGzmJL3sDG
RLEhZPTiV+Y3pNB4aBfkrnZL/YwBYRvNOlWFShDthNoYMqvlsn7Lr2igjnwNVrKt98Vu2h18cf3A
M/rLC9UuBBrgKJT3KMklLB77VLap+CjPFUytC2a4Lm95K+M3mQXzbznwfk+LiKiI9uWUlIcdIU+c
v4WmJYUm2RJpOc8KyhYlluKSOFg4boXYnxVxv2TeGYNVyTnZdWNYLdrA92b+yCV9+G+qdfNqbF7E
U8MPKlGHw6MH2M26736T2WGs3hJEp3FYdJyxGGKpfmUlj/hFKhgI7oQb5/8CcBy0sKgI6vq/5nAA
MoIsDlx7hcjyddaZLbuxTPErqA3LvJje0m93E80bYpcUI28wy1zJsmGaGfPtEVxKIkQnQX6fYgRa
vstUP2caPrnZHoexXlElJZ82gwkvT46/vJGR3TkRZbbqgCsdhD3iKqxT1Nk2+23pmDXyz2A4Qdq+
zGz1ICx+K8/vh4YkiwDB8+ZxIVRH6nsfOWWmnwr4Srm8nYOk1s0ojWXq2L0x2scnK2zOImLtuHKn
j/Iq4U8/oQ+sp0LfFOZQgFmAeQ1ubdtyJ9gVgFlDhGDVB76ON0OozEPk42atBjKRYQyo0Ml2lLpD
RLdi7snDaeZh5nt25YF2WKtbK/MH6Z0qvgrs7Nv7A+mR7vvDeHXdNz74nBWQaHOTi/PG9OQPxC3Y
LKiVFf/gDP45UsqgDkg0CylQN8gKzmThaYCcHVkpEytnHpKMldfLgOKuyocF7NAqnrsGG7dfVWJP
u3ucV1oxYIIBHezJU5kvBmWvUkU65yHWAWOTIvH9nu1Y8vi8mBCrbiL+QA5JisLiWdI/yDrjJGT9
F2zNOc+jAdcFnnN/t2xlP6wNkeHvAXkkdQfKN1m1rW2T3Kv3eyJdudcgrqLTVzkDett7VQTRnIEz
heAy1M+FalKFiCkmO4cU51hF+h4CKy1g0Qymh1yfsWiiykcwIxknx3nI87WmG6UugIcBq03gCic3
OHaGtHqW3XMTHuY/YvaGXkCOL1BqSRrZZmuH+00SIBWSGPNVrZSdlS5egRTcc2v+W1GgLLDFxwRi
7ggMGq6ViBE/ooA75uJZtHla2qQUjFEvS0SYY6rWCTn++mgjMGzoT7i7BnqkRsszrf7pck1mY8EL
ArnUALaF9eGwsi2fV8aEt7t2Mi/mo+jp5g5gX+zMQy1Tkr7/4Cy1pFhLXRpA/8xtIA2rLbA+AYBQ
RMUFSnealEft96ckBhKKY32bwYB8mpKaLQe1rgcUvlxVIdfAOV9pDpwiiV1M/o4JHA0JRot5NnpZ
rSCM2lEHvYGZ9NrWOP6k+WnZ6bG5HaN3rOAQ9JEYF00QkssB40YlErDmEq2ewZs1zLO80IBiesd7
sbRYL4lONBSQr+VuzrsZudyNt9VxfgQapjwJOwhJKU34ZPwUE1w+kx+iV98VGM/H+Fj337YuDleu
IR0abMHFotCuZs7PTmjYPbuIJk144T8mvaXFuUrhjQj10Kp8ubrfXUKaVWuB4O6x1HhuF0Th+T9G
F9U4C62tkD5oVvb7SPdWlctNSKPHntW4OHXlXsAuZY41CJFyuiVnWNeoeVub5O/eE0fjRzW/33xd
QQCv9qLd9wc5wbgoCcKmv1ZMoI0D2BAQDdTKHVobkLGDaPai+zzWHyuAU4/dbkY6+gfDcDQ6T7Aw
dUCypVPqkwmk+nzYxwpbtBbJY4p7u9m1mCWQZ2ci8+cQJLwxSVAzVIG+ZvzPhCN2OyGa2lOdEbbu
1O6GeynFkMtIjPrsTCHyoybKyt3qeGxSJ9VFHLvFqU1UlIJmsXHItn8g8paSRvayadPwAha47cEK
W1YB0c255hLdb43noRRFTQVRU7eXkyXgDgyarCnChElFUUT3nkfmoWNrfy8HeEcSRNxYBmwJKcY9
1UZ9hACk8q7BkvIPDizDLNfujBP5cnrLvE2n9qWGCFWO8+ISy4F0y/ZtL4QRfU1Xz6nVx3M1StLN
shQ3IiK8MOXNAopTbMa6kN4lh4B8muab83EhTlUDzjCapkN95zFKiaQJFDnDY9JVAIuDmrUUf/HD
euk0VEFuoMo2ZQvIVOy+wdQD39kFGqv+4rGZJ5+I6wcw/LjUO6zF0dmKC48PzL7b1VBVxhqCqcWN
1toU1V+w4E1uvAzASGDb59H2XEKeJ6TcvJzWqLqB1BGcm1oOtvBJ8NKVxyDkJl5wDo/Idp6zyq9j
Vg7YnNWZsgkHfSCF7DGCzknSfl1kwts9FmFAqTfrlsonix4nLUoSgMW5xxA91zvcHYmKZPmOdofQ
94O7k0LoYGNtOq6uayjzI5s8Asyb+/fmW6sHDsSkeqikvLqRNjvvUKq6NEPfKuEOJ5Z9Lc8ToKE7
lKFZE/AtFL19x7EoeRr6vswHz4agDkTBSRvRUEebojQnMMm32NRqf8iE9CbeC/a0JIRutSkoq2up
5ENE7DoAv7qoMXKkwd9xS3ZtnRv6TURfgbfxsixex0cudJXa+yty9KdUoq2laN3X4th8TkqXrU+h
ERUm+2UaAs6soLm4ZnrL933ggj/cKOt67KWa5wmQrIo6epaQrX4cNQguRQgcSPTstt+qV9/nlxZd
aYeL8suLEoMkE4TxuscQK/bSMmaza2I9lxNdQkkXPDZHV7hpqQKPfhAhc2+/9HEQaRK7r/XFKfd+
XMYkvO2Nn24JnFVv/ThErxZGjeyxqplJ5H5bJpbsh20swJH8sDXNk+zlkDMtusMBJTM/zlHoKncB
CIevNa6Axl5Qo0ePBqJ4/lPIijAm3KwJoBUMewWWIrzXzQHaWCB+LMsK6uhDDjJLATnbu2dd+08B
eNK3PjMMr4BWISCo/S3WOldqTemN5ZrUShUTu4t8nji8fZlCoq4qM0tBlUppZJIGwetLC/tJ2Oko
akT1Ssn3BPQUtEkiwvWTwVnLx0v1HlBH3rnsB3RpvXxHVKue5mMcoP24A2ok8PlXEmPyXqHQlTqd
9TMaXl8/Yz6JFJlIeDfZDh8N7891XiigeFpvlry66htCtiRyVAq2E69oHrDPOSJst9vIy8WAx1u7
zrVviQas+159lrX0048YJhO+g+sAmc2BoZQ0KYoiKl2kpkGy1MNK7Yz8UziyxJNuMRwRr5T54VAs
Y/cRM6bChUMqKCQYWyELAuRhfTdsL1qpjz/yNqWNzywnM631lFQ5lH4tUXGiRl5pawtr8As0M4/U
fwBOuMOd1M2E3XYo7Rb74NGQfq4r5LooKTh/arypILGIw+Hjl09HDqEE4CQdkzs4CJXyM08yUUl8
a0/QY7Rb+DtIojlVYFZnf2jZAHzZB0HaErgjruxEIC3OYxJOBYb8PXA5UEhPRYwbKehTGhxhkEMt
FmWAFGt/AnKpiE6OJL6Ta3pUW8kd2y2AUsZmWdeYW7BhewsftYkbUnNfvocTnvvx/a/Zhgj7toh3
+3MnTDgxz5Nm1qXYZm76/xsp2iG580K3CHWsQf3tAqjRfmdJN9emWXZ4WQbDyeC4csNCx+snhR3D
qF7Z889rWH4roE2o7uLrmWmGCMjS1+DyWlZ0ua5Iq5xcNe6oZSFMl7SIoR/vPz9NMeMwAdS9mHq1
uI7i0Nwab6v9PgGji24PybiMHwFv9QZ845eT3MCSodiMUZPqHURRSBwEp+1TZgOR2kOx7fa6GEcV
pICX81niwCczje7CJ9YhFpRxM74GRbtES+HpYlRrLRy8zAKm+McfeDzzUCRPnjLooOjZvu5ruDPf
aVokmxjOdpD2jMBuBQOF49rDsj9qRB3MfUe0yTQiUJHLzRXKutTVpjaG2KfLrl4URuj40HC7hiVw
KQGzJYdgwa6ZQNG2/HwELqRf2vQoV+ZWfpcRtMGOr3VbyOLq4Bloqf5BIqsu5A4JrHDzTYt1rIE/
oBcWy0ohWSmcWqnMHspRq9/+x9R9XeS7lxSk63eySEOU0aUv0zWjovbG7+wOS5BoA+rGvk2AisSZ
1QkJaU2ibazsupZtuvP++sRlLhML5z4MxTXhwNTPq2ZqC3sk+8qxDAnqdbqdQAyO6kz4Fw9HRK3P
pt6QEw3VApFsaBj8KJWFSvexoO5Q1denlBIeELuKujHzPb9zEVrFeZoKBfOdl8I3Y1yMS3iLlzVw
IzDu15LXx1oBaYfRAVQVlFDxz74/IyVwpAWInEyAih7r7DaidQAEEUtyAQ0SpQdDzJrWHEJkwQM6
FbC4H/szRwURO+pj47LiNN43NjrpGfmi5rH/SY+P+HOq3S741BGPn5gOASeXkorazKVtw+7WZ+r4
Wx1niR0pQDFePM3eyrX16h9w0k7Xwaj2Wxoia4SmKZA9SQBIZc0rWWocG94vM2G12lHDeZp4d1i6
5uPq4gWNh2gqHjcB1Wkshcc8/Ukhdu9QeANgtWfhios3Xyuz3aKjuwS3nKWnI1JzLCraAt9R+TJf
dVbO3GMEdNRHp/xpcaIbrKpaVy/zlfmD7k10mNfgjJyIZ7c3rr5jWFrA1ZTI3o7KwyCcwysxkjpZ
7H2rxKj4dznT4BH7slzspZ3t3vXhGEqXvSyxi2tE1fiHOJB56QfEjWE2rxcDn2e9ehxbZO/x0qEJ
gfNGV+hbPFbXeF65HfyThW/4fb6wUq/f2Jiu/fZkK08SYF7UrN37H1ZqDXb8ehqN9u34xRk5CCH3
XMHPmQ5+rxTm/7BxVgfxNVZ841WzpKmEibWmveNilrbDPKDWhQNkS4ZR10dOoN/YhlDx68dlusGK
UC0RtcpINzX1G4Ke2WSEqXOcuDLiQ6G5qn3Om0Lgh8xzo/0ObwuLYqZced7ybT31r7yyc2dAlMEt
4glGmQX0OUN6VeV2oFHODo6KlGwIAeWAv1gk3uOJPcDyvqfiBut1cQVD1nwptbEZ/HthCqAkDngQ
Ha93qo4gPpoxWACUBA5wH4RjSM6RM98+vC63AiYEy6tn9JC7QFsXNxYfHflEnC7Nbo+DSVQVNDEC
afoheVPSq8iYdGf2Bojoyaa4xT87RyeNByO83Keh4oTqtHU7QjTGSaceCR4jHC8M+LbcHnaO48X+
Qesz3DRrUxtOSQ7hq/kPE+aVQhfFr+UKNaHYM7sRhTiLFB7ECClFO3m6dbZeSb1toE5HoWwsF24J
FVwSqmuEZIOHUHRPMRm5pRGnawIN9YRxelAJWSv6O7g66nrvXuMtcTB1Y8TPJLq6PEBpQjrZzZTf
zLi5edOGV6tbAMnVg+vFLPx0ahD8Z5o/SlrKal0RLtEoylcTQswfBOBF5slpGJk2sQ3eNRFr/6Ng
GKG7QBnabIe+MhNh2Izx5BD90+855e5sLlMzVKYYgULxtyx4nQTAzDGlluoag4gT7sJBsU/PqF3A
l5ppztCK65uOU12EPBImrVFFEOZW3oLd4RnX/cNSvToPIaUW/Y+72Zqy2UCNfS/p/OSR+XTtAdRS
6Pf55d+E4HtGwuhLUib+ViOTMbqDLOgDXCECOO/I073y9CWpR7aJSm+JgFFkV17lbl35bmbNjlhH
D0dkQpnZLk2eaEmyKrT4p7YniQoxFwX1GbgxcKJAiPLB2KErZjmOwlhtu2bV2nAY2RmlBxmuQp1U
4mRiIYqGf5oTgIxba3TPmbJVBIhaxg1cWLuP/ITa+jEqKWAYvnPS7fPsRWcdfAqRSIx6K80jB24K
0WhIDDat53pB5D4ivTmlLGwqUv1yzS8pw+8ra/aD4N8GM+Ijwj08mVOYKydXzqG+l+FJXYdlB6Xp
1EKtTB9WH7y7dnXlqELzbZT5dKm5SsMlyLzw1mzH866e7xTIwCB5KhTAqYeL06aVmJUJodeiNWrg
sCghrveSFS5TmZ+pl1rrJONC1YKeCgC1JAUyHycmD3V8YcILj4dHKt5CzPd8gHTGUFvnRnWS8SYi
fE/47EEJf9nBoJ97FjqTXVVODWD5CzyLjEZRULyMnmKC5H1hOCYFdlKWW5yjVtYYyLR7b5bkCuhl
ju+ehGHHxgYPMGtXj4r+1kYT2Hj1U9NkIiSZBLzA2aw1iTzeelvvk4A1SzG5g4dEKlKFWcCGCuj5
1IkBRaVfiAZmu8ohL1oIBraODl1gOMSYGBwXXRV4I+9L6QKhw6CrdeUwX1n0HbR1XQNfIme3SmEn
v3OvMTOlidgqWY6TRlJb2W7JV79bkAOtxG/IofGPz2HshqzHzdG45d3+VgZ4V9qof7jCzxShXkhc
SOjQrrRuVwGQbe5RJD5SGoh1mDbh+i2s8fg7CF4NxDZ7NRAtup57bdeLjS85KbZEhoBEBHkF6Tt0
SSFKrlcq3OSDYA3H+f+0TCFz7yb1ZO9EGUndQWIp74C+QcSaCEF3hALfrOUgleN99Mz486/qQIFX
u9SgUFAVwHhlRiv/yJpl+XZ8Js15hRSRpPalgLGV3r9nUfvUAVppLnZdgqv4Z2KG8ELAGEYA0pfb
iE9RKes6abt8P8Dd812eOx2L+ducyBlZOZrvUkozqnGy7N0uq1g9DckLQVlHVRHGZPwTcSNAN/Qt
HQQPm8sSIQDfG+rAdPeZY+m5ziaXWWHO0aiUakAWKSmjHFFiHlpThEdLDZiYUcJ/3IcguSj1R19f
jC0DomnxxmqO5spJx8adg4MerLR6DornnaPIi85hga11exatkKYiLtBbhwjgOYLU0RC3gg0eInzM
jLOSLRpRqKVAIhGoYUBCX3yxz87CKHxKtJNovzD2gz3Zi4a3yDMUS5HOM3rEorzo8t96qewJTaX3
FWst4opsy4JobhHJD8GJ+/jGKzX6SD+1ZRDejamlShXs5M+5kJ1Yejx7E1kJKLrXC+s9zjDtZ6I4
zH701O9Es1ZVxcNHVbCAGryqGD5ulRvLgrmfIx7b4Zwbid4HqBJNMN7EBnjo6XLuKvcVlmQOdiF5
Quql6kO1muDqUOukBrwEFllD4eNphlScB3XgmFYhNIrnWl3dlsNkzSPmjgKpC+XoCovZ8jSDxGWQ
ucuv9psOyM9ZhkeBXVTco3p6VR1LjChyzvX3LR4aY7PYMVfZHHYd0AuylvYuhaGFqmkco+qq+ymg
jvjbLKZ7fINdzVUNX0DyGlxuO2ceIHnBbl+eiV3b2RRR2Tr8H0fQWHNcryJFBTpgBhseWosSqFxq
H8ASpR2NjvazCWdjamFxJsckSiqLY2C88KqY64DKLMFttf2NCh2hfOTgAF+hM3NGPG9iZ/kkAogL
CEJB/YuamfX9Tc2kkMeqp/s18dnr/6GF887nT/vUmUSDfqIwZIdO7LeSQ5nt/vhTYsS7Jel5PgfY
M/DSMi8TjRI19sWpgiqYR9UOZq+OPMMOUT6d8dYEVSPLkpaaLEN1qN6ON1hiLfFCOGj4QWrYbc4t
4d+F1/WHPOd5b1+ux7dqaGqJxZOOQ/xA0GWmo7fJ6niVqD2cAxPhiVrIjdgJ44LINa3Rx36eHM2W
W9QIx9CDIF8f1C+82lIJWa4uGRlY+bOj+u+naACWE/Fd5TGkDnAzKGkLjZtm5sdMjcxUp1nWqsaE
YdFBGNpGI2hrhG372abXsnnAfT6nFedGcRc74d82wJzXoFYYI9SbBS/hcI8Pn2qrZFUJRQFtfuMd
2GscuZa/a8tAT6S38a3FZ14XoUx0jwabirn1FnU4Bjho2mTY/lS8ReNVF59GqcgGsreGAu7s53JG
GoV2O34f1qlIc26xkxGsmpzXnT03yENfXeByFhIUkmn5lVpWZyM1vH1Lf5uYC9cr7Ji+idDN/z4V
mqo0YIMHLPUmQXc6RRqzWh1+Y57jcEUxu+yPHpdQOvGt5uGvFxV5pzAdeuX8hAzbkjItNfHSdwCH
X0LHxK3jwHHZdux7iY0W3ecHIb5wLPetk/yF025HjCWKnKeaSGSM0SgOwY+GSHealIrKyFMtfljZ
/IcMZbyxB0Fru8fR1ykIw3aBLwAYhQaAOHcLzUYnO6ttzmdZUoonLiCTS+Dl1J8fv5XoCLq6mg7Z
0qxV5PAPPNnmGdHc1J0AbZelNLTtmsozif3MWkGrDhiRJDCeyg3Lr8oxIAUb/C3nP16PBK3DvnWr
dO1xR29K2bv0ydO+oRfUuf7PYrt9KMgJ/1CK/2l11/Eu/PQoqJEPXi8C9OGf0F1IT98kMQ6tlI6W
gnDnZSrdan5pfts2yvezJs5DEiqMDKN5j5it/+emwH4fGjzO3E+PBWwTP1GQdaDYsP0LaoTM8nby
WyY8TvrivaMM2e2QSEEHK7qfQKmKX6T54RNA3zVZk46DiAYV4/5/xpG6LXQ2+MLu3fgpSsXCbqti
Ymxt+aS0XC4dkL1FpbkF0Ay/hp0vsW9s8aCvSytwb0FdNgtoTadLUbiWro4o2jP/3X4GK2aFjY0L
cYOM2SP/pWJNkAOC7M1cO1G/OVhBX5PTpuus63EbeXoQL8cOirsKF2+yq8HRP4zjuKk7ZbhOAXXP
XI3L2o+6R/6LDNzaf3OcjWK8SzaBTuYq/wuaBQRDjTCYcqdY6kGsbX5OWT2D+GmWfEszBL3NF3SU
A1nGrB/YeJVWs8p884fiVRKfIVK9YHZvG19PNDvd6gpoqQSFbkZAVTacFdUUfE6d7GrRzVpeoE4B
6426gghIPXRCiECNH0K50B12x0p0IxnfciJsjoOBhIrkumXJeEYVT5GKV75I0pLYHFE8kzMOYY3i
jjAx3/TT+zXSoiOkDzwnsJ1xYlk7/JEbsqI0vy/uj/+Qp6VzGFMT1LD6Sn6/yLSM8w8rkdzAjyrP
Q1ZG/D5fJ4RNLxZR2Sz9j4uXVJCEgVDxSt9sEh8Km+p51MUo2N6L0KcneG74asyPQwHCYZvG6+Re
L9vMgI02deORN5s6w4Qk0XaloC7XldsqKHdr6bZ3plKkVDotbrO2t3O/M7PjM2f9g15Bss7GdEqN
0zdO8oftRZBLUFwp5YxeXzaANU/9w7KTuJHl07vlGCe/+s/1F/5v8OB8B2tMRNzoaKaw7n/a+Nea
Mn62dsuz6kaTBmpnWF07NFlVowkpdwideBgundDTjL/qAt8bOHHiAtT7Ja+74YVNWGRXKYfxzApY
SWTe/S0ax7j7frXPwMrn0bk+s9oSq9EaliYGeJtcVSpXllozwW/IOVXpmb+QbSCkBlpPw6JAhnh4
OdkHKi+0pUnLcM40XdM9tcUy0Dq1aKo8hwVKLSDfQ+jXhEkjPEhnqg7yTuCgnSChZi+ejoyQeHMc
MDg19F1t4YUWkop5xgMj02z5yDGgkLs8XDc0xPp2nBE2+C2ogzwgee8LuG3wHPs8ZlicO8bnA7UZ
whZbwB3LY1oFR8AOzW9ketltfLlK8zANlgMYQm0RFpEFtui7LVoRko2ZpU2/IMRH4Aj5ygkw8nYD
DhTjGJVaGO264Ukg53QkOMb5Imi5b6sGWVQJ03JLmO3h4p0nF/Q94ciOkMchmUZt8C9LPwdFz/Go
TI+5MkAEiRNpXs7skW9M6pDtmkTbLyvgiqL+kKVUfuflDaVZ4TRVL2XYAv0nDYvW9FzOp0/o3+jJ
ZS3Cbuj1Ktdpv2FKIrpE4iB2Yd7h5+6Itp22Y+0ZtuvvZzlXxiRrzGrqIKLt+JKGbvl2/3X/oiU3
SszlZf7LHNHt0FJ4BhJE1QW7DQ27kU2vp8ZqiyhYhupSDIYRVAFCOyZHVckkwVSgXUnjRXKiQNra
dsJviqS1TPPqBR75nVZQBx92Iw91GbOsRFrlsUD+SHxT+1etLxogY68mLyKmxrQaJsqyj4/1R5Eo
vgCZ9QZwSvl0rifSEYSIw5XqyFCQI0W/2A+T0aQlKjOy1IwRBtXo2lTNruLZ6HOBsYj0A3oaUl1O
5z7QLK9cWr4392BCA6sZo9w6MYfR4WvTNN17wcMbTqEwOTPexATWQvsfxrD0wRJvT0TeY46lplVf
Bdf0oNAeAfty22o278tsyoR/tzTDkgDh3CHnCWOmJlNHQoSE5kqVqjCgwF0AIF7u3bEQN/5KNPLP
1qrZlYzhklMKyeI1RmVGr0b9Mcy079sTX6MbJXvQfukoVmv+hjG5ORcGo8qutiIr6+c3mCFcrnNJ
eKNWHzIE+/jzHtIvFmmlOi1ATxwO8G+dJ0kll64H39wch3Iz8AvgzCFTTRq2P/OTI9wmXWiRTEvW
CktRq6AoV5mQz7mU4+8IEPcUZQFWNSaVkr5oJSWLnNBAQPhNL4uA+RHc7Qk4LtbFtcjZd3bJ535n
YRP6EWv+rPKjEXmDFGqRfH5KjwyISU/3XWXE0mmCfkhEWSEck2ELB9ikKRVqiXSLshAAFkWw29N0
dMmc+bsaIgnxthxCYlQJJOjYrpr8MzvnWgmYde5zt+NMTg1W3cfanQCl7mfgmb8o8C7mODbaOkJk
mcO1h/F1OKzDADtg2cU6LUBQ1HX0YPHwKqwMMy/Pf8mhxR8zp4Y6Ld06xUjI2ATbyoWRs49ihhj5
hYOb326M/x/YL+QL/ud518nhabMPAQKBXRKoOyYh3s2buT65jQdFtFzbxGposK1TWLGnu2EjfvLi
UDcu4UyCE+vBZSvkDi1K0pR5q/P0lW8h+/uf5zi+NTitAVfAln1TqlVJHTAT5pjmRGgV50HHYGCE
6kMptaZam9RKdtTaIP3apJN6oCYA/tsbZf2TM6CQhBUB8TEodNFFGdQNmoRBakJtlnVaqVVrno2p
IJmWQMRMhI9n2Zc7BqPdwBunDu47OMEIcU4fT1oAK2payiQj8OENcsJ2CZDUSLFda9ePqRAZuTda
49vw+DIXUT6NSIhhoWXStSaWH1rDVBMzxWdjdFLdi8xkEZ1VzhF3zoij4cd23zvrQQxa+ia68I77
GUG6DG9Gx5DmonNsdgRPyDxeViit3BhOMg2PHoJzwjWyzlr6mKSVSH2/C1OEX6QBXyouy3WfhhTT
goRw3SCB9LUdOfmPv1IsLEIEor6OVDUDWEyqkthC/hWlhEScPVooCRMp+PycmZx1IzlCM+lfxujg
rXC9ZQgcpgz/AcEVcNRsr5zZu6rmKNT4FkcNMr2i+SnQCDcKIZLzwTho7eP49g41UzF8rEIVBZ3R
wJfh5Amn3JxpsIff3/VYLo+1cRcW6au242JepCAMhtfxW2SYWCUVi6nA5NX9oZgRFqMI1TomTthX
rgaFfLeRRBcUH87W74ZnP+dWvo0rOJqGXX8j2d92KMTZSQiaQNPOTheASK+5GlzOKxFuk7QZgZ6M
y6vPkzekuAsNOja8fFp5YWV0Eo+R1MDotJB6538Qd7EdXZuXwO7r7N+DvWhPVy39/VLoTTn8OGG5
d//3ph3qecOsuB9fGn3FFNSXjxX1JYW/ia5U5hQw4gcxNMuwdQvcZg3oXYKko9nLg1yPWyDpKDeU
lMYFzimEvLCyz/KW1l7lonNAsoff+/GZN0/lGQFuN/l+0RE4roBp5W7h6UZqBP2lcTJm2pasosvT
9oCRAWwdCrt1QDnxHN4pIxAJCJcg0f/EE35br9g8y28l0xrVWmH6oghv+D8s/lilcy1X7Hp2ita2
nBQK8K+ALSSGiksH1hhHlseu0gAHbGXZv5LsxM2mh9m4Wbr+DPXqHoBTDpwZnhkZHXWL2dQDvDUE
uC9q/MrlAsI2ecr9n1MOlJxI5Vk5fBtgdejPpkMQmqIvJzZzujxKRrL9WKP6eWEumfOBlWTzyhXq
ON4nClQOMo/TAcIrscDVOlqCPcUtZeq9PliIUlrFWutGlhO70j5Nsm1a7FmYZz/iKPZT/05TkNGP
YXZiEVqOCOtSmVTPihMTmzvlDGxTf0vimSyLjxDSVpMhPHgxm06yQWn6RTmArUq0cYyE6fn6yUn8
C3CPt03+JSbhzNWwBx+W6zaJNTmOU66WkLxTzQ796rBy5KyTUc9VQkFZoG/8q9kEOmn5gOuMjmvX
uS3W0JuptHz63mGHI0b32YrDs+9tJhQHPtLNK/k3Y4FrV4ErJuFZFcV2tYrRmEutiLDYJcAz5rAZ
LYaX7e1EJ05dU0wMZenRs6TRDTCQLB32j0zpKqRkv3yClUN/7mzFnJvS1mBG29lW23bUbRA6hEj0
2evURA6QgssL077P2eBae1FHKunaxgiv6J3XqpjlKEd1Kg0zL6WH2klUn/h+S1t3VdG7Vh/dfDqN
nSE442GKc6/siuhtbkdgTJCOSftxd+fpjxGypupqlPEumJh//ZBhIJAxDgQ3IBuduke57oAWRGbQ
gI/nrgn7VFaHRXVwCsIEd+to0G1zbZEcpkFNAC2jrnI1OVwRAbxRVVhM7RT7FWGKrHQ0DDA3MJDR
8TMTyzjf9Z2M0H3C/3an2NRfnceumqMyC37a+YYWZta/jS1DrvOKvjq2u8Ax4d10T7AwMRHSFJmm
rzjQTzaSuvW8jvtxtJy5YWLfmYW+iYB0T/gMqDI/m6b7PZH4t2ZWv17fMnGTEkumBpeGZAl59x18
Qah7gNgpeijPXVW8SDhvGiuvMv1sz4l1OJER2DaqrIYSZfRoI4AiPHb+6F8gb+dANzdtTUePtltS
gzpTd4p+svNt+SQVSzW2PPYP07xjCt52piXd4/2yCIAKe6oNcfk+wl3BWCZ2kzIEgAx6FJlgymPF
EXqBrKsWv63KO3CYmD/1Jwk0ymFseygMTH+l0Vcb3e4YD/4KMuCfkP0Cke0CgQAub6q6C1gJcFZx
BiSr+lPQGPH5GqbaQeaWPADyyIxxI2dZhv1HkGzvjKxtuQyh/E0/5ayKO0pxX2rfjhE8EyyMYCOb
q+CL/eFcBI1M+uOUzenD/nMZmKKIhfe9YqqDCnqj89a9H/3YGQQobGfIxMcs2YVTB767gcWaRTZ6
JTMLnwcj6NulQ+sIcZLJP+8CB8q+nwBU1ozZf750g14y8AwxkcvrrGi+H68llVperZo/1jdxGB2u
4OaW5l/I6qUAgj/XH0zy2rtokr1ScZ3duJ94zEKTrh1S8czHoiVMUgXXhiv531GeOzpH9ccCe9ul
MzRHwelHJDLkAcdXBPosgiHNs+hvRgbrVwc5cwQXVLgk5QHBN+80ppvhtwmkN2xEX6PpDWewzHla
h67XleoQ04KWCsdLz+9zt+kKuKVre58GdFuTmgFRm5QnylZPwEzGYJnd4NbmY9cb58M6wjPcEzfw
/IDl0rwKitQBJ45dQyWwcYOE3bpCgPxbMyPU4tsa1k6KUs8lUdhFRvf3X86p7Pe6BBYqgqsmPl2A
cGhcusJ38rZbccY5nK2HfWtCwJVRwMsH2mwI7MWExLEE5IwtlOfDw1ezzB9zVYwQgJ7rSRdL5txK
G9bNGQGVbCP3Jl/0Ovmv7IsQAg+vhALnettKXQN0bs++PFcWXtfwpt0BdShjY5XM01oz9dVct0Qo
lYqDBLkokTKyG+E68rAr6KeTVshW5BkBLHWAEJWxW+bzMx3f29qkw+7K3dpbEGqcXH5xyfM8nDff
K1bw2Mv95wTrKUj9m+9MmPkqqRWk9Gy0kfLsb7pK5b+68M2IuohHDGanM2DAxxRntN70iIEze662
9zXi3Sg/6cx4z+H4PiXlPlQ9lyxh/WWaWV5DGxgVAVQXXWCe302RlL6Awyc25eE2bqJsrYGeQ+dx
SVFHGUyq9dEZtHrKbPVK0JFvcKy81SnM7FEfqzLaAvaICZ25NERfMB6A+tyPOB/l5K1VAdZ7vEw0
9Lh/1faOaAsTXkyxKAD3V74oAvtwaNf04DZEcORnJf4iQfI9DbndHBfY/8xgL5zHQNIMdHSjRijM
LIXWJG9y5ZeJ97UEat612VCy/z5oV8IEx+yC0YXkEOYbrhkyw4HfUPpCbZSF4Je/ACHU9UofsaZK
OUSnMXODJEIni5o8xjWAKzVJW4JdOOI/f594TtUB77zRwO+1vjVD9XhVIsJBUpA3HtwZ1f2HhArF
hhwuVEA/CNvpaiSYYko3CLHI5iWXPJEbIqjmBSAoobVjyi7iaNA0TJgABwgaMW10kqVqccyQub4O
cQxckRBgQGzckC+4qXv3LiKMZxTpkc19w/gPa4DGO/mkkN63emDnJ9apF9sAp9f077AyiSlgTOoV
TrdijymmdOLkr45rbIlT9xIpOCkzOJb1O/ELic5+x8J1aUCZdVbEpf13Y5/rabLfFOO0b+gQRC+L
bXHQbrj4SUljlQBsKdtP3FxZ77uL3FTek4oKopOVgyftyIulfyBVgSFRWQTPTNaFY1pl9QKrXgTL
jEIiEZDYX5yGx1Xg+cxQnBb1oRNhk7ueMO+E2Q3H2cmAQWnGCYPywsXfMy8tOvNCxHaKUEIKyklV
+O1N7uRmR77uSPHthumeU1+tpcFvN/zNAI44Yt+r+j0tDPsqpWchVYEeOEiyMQA+br91JmlKqmBM
W7aVqbgD6IIfVUBxaVdfekv1ubVigv3g5tqJ/QZVJG6ZzAmX0GBMEcYdV4wLObdLmc96U7O+Afmp
INa2o44LsTucHVKFgA1/h5GGGcPDkhf0GviecukxeBdLmxVmoRxJVxyuU2OWlrNHsqVdLRZbLzhE
LBz5iGIcJW62uI3dAAchADR8NiDuGNrarqPM/jZKHwhoyd9GFOmw/MvSvze+Ol7yhdn4JL4QAgw2
jHrkLFFJOP6mVLIce5lcwR6Kuyuzv21p/WxkJjKmbBjMDnx0lXz8vui5tBcdUvBNzCySi0dyniRf
6kmTSezPayD9ae+Sm73XKe0rpvEWOgHZy0h6M30e/QcPAgqEikjb6DamSiOl+Fiyg/swlMuRCZYA
knZBXGwjO3YbRWHmPJUfDy92FVPhfvDEBt8uJ4Wd3ecsT81tWqAbVbniCMN3y2zVbQwRTzQzIkkc
CWKcBSLL7GPm7++ULoq4hDiTKqGXCFu29FjmA+08DaZltzJ7fn3Vh66DhmAlDRU6SG1oOS9eDbMY
KwoWGsG6LkIf4umoLVxqugo1oK5jNPng9b+wuss1tKcAynTguwxpEMcjvqpt2QQpJvdMqyEfMlGK
PnkYa7r6pMy4sNbU0M1kidtjdLHi3Dv6uIwcbQSkhK7gXsJh49KyEQX5Ocxf6+2VZbPSjiyufscn
QT4zwnVQT5fxSTZhAfT46h9FK9JErq+1hhqJJo4h4/rOzCyC6p3g3iK7e2IwPjTLgAGe+PM5/Kis
unXhpbD5KufqmI7My4obuaSeZ6AN6BYqMfv2LAdIbBe4RrnZb9eh3NVuRWr7oZrDadrwAlXg+LSR
hpPKBmAJjYHLxzDkMbh/vS1nIuMQpcKrEmyNXYkOBxP1Vekt+ayoo/ZK/JqUmupA3PHYRSo8gHLD
Ln+DNEkxCn0JJsv+6xGCaRnXMOqYe9c19zHlRre2jz2v1MuIfOhIJ8S5VHkxHkdHDhZ/t2dGpoHZ
GQmB2JoXBRbLGOvmLpuefzVw/qrhdf5z6F8SYP9BUcaJakzauNChEZ84INur+laJipq5j6ZirPlv
f1svnNHKEfVGj+4ITAePMfxuGWZpXiLVHZHs0lqNoDk1RqXcV04oc41k1Mcd+e7NyTHPxN+D3rTN
N4tuYEV/UtTnP1skm8y/ttc3XSGmG+B2UOJyhETx2gpzF4A3JD1PqrKEXoj9dMpqSjilfPEJtc8H
0aQGyNnXGvxD8i0FUYIhuFu7xeEKz/uWpBpC+qI7BVu/nksiKXoVbX1IhTXPN+zRlvWuGxmH0ujD
azlapLgPWly3MyQ4iyasDwLiUVawQshf8VZeayUANjNeeQxWS8PUdxjhc5iIOMyC2Ydf54tXxRpX
/SQlVwd1GXKogV1jsfW/idUaXakQ4et99DCdEKJF3ZAuusmd4RdsNvyV73oAVYjP2Nh03TM8zUJD
/nFBuG8AEsxjaY9FRWfcDmZWkRYs00NfyKgGTu2PZxd9fF9HJzYKuGl9BMzUGvzHoSDxxPEmzOPR
qnZh3KuosdgDr7nL/Vn22XlIl1UX+N5n6XxLfsHdIB6taqwm3yKP6MiLFW0D7yjpTkQSGvX0O6FF
QatJhSlp9papnbX9Ff80Y74Dqgj7p+NaNByaXd9aiRkN3FCO8QGm01rHnpkc5VlnvfQl+fhgNd75
LdM9Vj3Ev/gGY1EZkP3YF+IrxhipVpMSo+iLKykDRv9ALs4gkqpecHkSmqikEeNPYKobjOJpy9u5
V7TnXCORVrQAoBk6KgAoKOyx4j4TPw7oMOETGcw1agrDCH7tCbrKjf7RkiAjfVWx0WAxLzD7QEks
cXM2Rvkt1GoNNc7JqrGBFYlpvREWDQuGMfl1xZjuKYXhRF/3QYbAZEmFRINOl0NKNyxCdGTqUf9v
8r0i3Q0psmPowasa9ZdLDSIhX9a7rD3MhoU+CdlM8Hj26JzBybJ3Pft3HCjXXbqKu7E2nvLBCpz6
HC5DoM6TMRQR4e6k9nfSUXqvYZler3udPwHjwjViJq6MtHmzbdHPRl7FUO1ifjs14u4F/KfNLlgt
dN9anQkPGTK1oZgAqc4ymLxnLYbciVmeM2gcrIJq7jabyXjX+rEoDLmDhl7OYuvT0ZreGU7PWBjl
O4Q0NxGO+jVKZ95KbMslSLaRVnJdNN4rVPSfroDHqqnNTaNUqs9LIDo6iJDP51v4Gy20M0K8pBYs
yj5C1KBnK5eoAKyMlym32fh7EWNzOeODSYAp53c8e6KONxstdGpoubjMrzEeBNB7Ma3Q2Q/3B0rr
XsvJuPj70rtQUQ1qrkQRvYJrACFRAR7fP0GYMcP9OMsTrbzzotTJTLgy1DuGCwyrHEyQKRoUm1nN
L2IATE3vMGm79m5sizP/g3BWN0dPdYtdZHivyP03ntWtt09AjmGZ16aErOVq1j8V6TpVxzwZC2f3
y/T3w4jYLOcz8t1G27BCfDdsk34Q15SI86BRKv40Qrwkq4IddKo0J0LNktkkIvVpLLFAfcVL8PGZ
qGMpJTkB3O/KW6BEIGcg20R0Ldj7VyzIhfzxTgxKcn1KKTVApQl57Ui9zcYLjQ32UB69cAsH+s+O
EDBMLye+U6RlhLJ7as6RxHJpAxuvNl/mN3VIPG5wvGRER2h+QtcNr4psSt6nD/RCFsA7PIS8/o+H
4mTXZCgnVrwXcPHkmf+6Y9CrHqLPlfpHWhNRdsRm6oQ6zba4Akr/72OCbtVb8uF75B3XLCXFdV68
UWc/FEDHJ6u4F4rqyo5392RHtWjubmezfZ38psh64JLtrOE876rg/0VRxjA2Mmw29F4adHyFkumX
wtkX5P2V4fo5KZOCBxm5F0zxLGhcYwRkYaauf00lB+PcZUm+pLxJh64TvlKrgiQdStNveOF1h2Qw
6Pl15rkN8Sbbpr7N/1Y90Ec/22IIlVm4HB6sNDsBkM+2RCLgJD1Vlf78q6r58ZvVK/wY41+8TGTr
vAPDFQ4l15dMXPgopLmNRF7QTrF+2ve2LXB8VnxMp21g2EmxhFL4rAt2IXhHwOicMAvvEN8vvEaH
je6bO6JiBx/gc/IHRa0wHT4tME8j1f6u+0Aj6owB5O2AWzvlf8lUaH2/QwaRUMQInoZrol5wo/SR
Yu+FH/4qbzRK7HtNCLJ6Nm5xTY7auf95/1KhJBbQwbKTQm3dSiRmKTv3o71c1sXV9HBoRA6YA6oi
m7SQ9iDk4F2UVac8MAglNEfnWs/5rekR6U/OgTPsHoICbQWD//61M+VZv4BkUMhJX1c1vtK8hpHr
uJuUQSGztPDqVG3RfySZftJVKMhqE7rwWUf56OapCEOe70QgBubxAWlvcvIBj8fPD24e2510iaVD
LadDvtjvKnYsfmaPvj8i1algO+44+rqJoEXTrZ1Q9zosVA79C+0E/68qrW++a8UY/NPyCUOezQIF
318m0A8L+p+e1P8t+Yd6gTXw2xmpI+Kc87L4w0WlYH2TRm+I0DyjNfhaoPgDru8cJxbDZDjFUkOZ
Xr3ccyC/EbF3GXXaeraE6j09QA5hDsH1k3a2HZqHuwAEj29CpqzIHr9+YucttQ5NNHTKgtS7Po9C
jCmFBNmsE5npGBZLF2GchM5qV4p5ekBgY26/SVJwJkGgAEkihilipYfd89iBb8FZjEQBNOuh7uVo
wae+hNUsR2tOH7nzdvqjKqJW0XZISt/PaUG3yw4ZWJHwYR+htkxwpjoJKdx6FlCo7YgsmCRnV/8U
y4S7JQ3yZp5JzGIWWM9hDRBXiTntw81LWOHioV89JWbxXzNop2QLkUtOLIWvacax1/aK666+LTKn
LwyWCFwgK2EVijNNGYGf6cfxRdDc/rP9ytvQC43klIpxCzRHEYD7dkYe94OCNyJWdsPcjeDB1Md7
uX9uNad6++4nMVNiHY6KeWVTgqPvpQ3ZWIHbKChvIs1C5DhnreuLcuTwF1889lqrFC79ZaL6k/5m
WUGWIN4I++QfgdSbAOvGbHLn5p0pOaQ5kA7/de82iqN/D0pj/Y9RDskil7kcc9vlcnmv8hxfinxk
XbILr27EjohZaZDsTwX3xc5/MPOlooer4zcFc0sdKdqkJF+Mj7BQFiSOHS5iaqQpFEYKG53Uun6q
N/ZKCrowzEDnPrAbRD5ZV6nNNqRDQQ9M1+THmpuRIgYaxwGP19a7gdJZ+d6imjNAdYUxutqvNcuR
IOs1jAteYPfXL2YyPSp6akTa3oonFMQ3uTUzuyQDR52arKLh7/9vQ1HG+EyTDO1oHr/i9COZ1v4C
UtLxFJ6aEfQDJCV+HjhTWvj9uSpZPfVpecpqjt+99y289vnKVaqymHvZA9xQKr0627iPA3x8glwU
Mv0liCgNETwDoIV9ck47kDH4DC1aY8w+pESER35ZhJEL2XsvJU2kr0czW2NKCqiz1JqDae5Ef2/i
7gL6TLtBrAO+S5Uw0ua9uh6FYeRw0Ay8IWtnSFNj74VRB5mm8wSH2BioP8GVIM32mN68U4f+5L9N
T9a6lnXJc18PJmhCHbFofyC2F2WnwA60SMNrukaR0r/E/nA4tMbxVuYVuLLZ+6S3Cui6WZOfMiJE
qZdiZvbbRFd8dRnWauaUXSaLf9StHFe+f6l01RlOXYt5wrjYuSt0BeMt3+ojgPQ1Nd3kBC39UFIi
JQcL0E4I4/S2DDAQzlTRcK8OE9C50yALo/G3usr3YeU1x+7nE5de2E4IMUJlEJspxFJcXtNG3VL7
8mP4czHeFTAcei7Xa6VNc3sdJT381QsZiC7f0cVjTw7wmVKJpA1/q7a/KkEfKPuO3/nPZ5ZwIG3z
wCB0hjCNEXLBBB4iiBEASVLrE/2NryulOL86ylmPCIjH1QnPAuxjxEUpf93AM6pvxF35wrSHhkEq
PcFy2jPQkoJYeEzXxzXSqLmVEPXwQF8VhhrlVUHTxu+euiHn5NXkRASASd8qWFR0V2t7Dymy9Uld
52eM6i+dNGfb3dSV/h3jlxgr3X7RUGS/qs7z+gDmg/8BI/YdK6AgJj37LFxBCiEZj6O2ZlFi4MKn
fA5Eoln+TdjRuaKJOOx8VIPScoSxpecjJxYdSm9odgovFF1oTdFheroPpuEHQKY6LvRNqCkUY6Nd
8IeOeP7rf2RGbYKov7GztQ20CpHFv35X31ZT120Ssq96JYlkIWmh08+ToS/g1Le78E+A7D3uHWLu
3IvHj+3sCwFN71bDiEGGbpYtKb+rGQ0ABZ6VgrJETqJpZ+ZO5KZIVuu3efea0FPNqPIsbCaR0WP0
mCKNsd7ztjvQuX1Km2+0S+VF/8LxjQKgoLLJOjEdoQqfrVQ+53RLsUoJe3/XZtUE1hAZAiDvPWya
voLYyTr9OdtmNCBwE3/PAdv8qvdKXXMAB21RzeKOIgj0GKlg1vwF07c5G19yITVvdTrbdy9KYYed
LMXz0Qgt7R0q935oDmnlvkrTrunj/s95hVaLV3w9Y5jkc61i8KUqH4J+PpI8C9B5lDnUIGjGqVhK
S0dBuGCJxfQVfzK5FnLFN9+n2ZO3iWhyLR/TC4gvKgXEO+cN1jjyweHNC0uOmbeW2tZu+umLSF6Z
MNrIOG+tdm1iEtD3HeDK1whrY16E+6v5tJA7rFTL65d5jIIz8LQ6bOW/9vUizq2UV7U36DKOEBw0
B45N6htshWLsRFSdOV3qEZvoV/aiERoGjVRz+CTW3Tv9af7mncK/dNnj4YlxmdaoSOm0aBnJKaaT
qgRLaOUEzOvFXSsnNhE9x8BXwQ7bCRT5Yx1drCz49kHje/JDgpGlWC1aWP1qYwpi7hEWHYFsFgtO
q8BomkKGNU9iL53deDyccRIMkIlT6c7AMo7EujDEGHxsvMVfODh6Rzt9YWmJ2LTgfPDT2xqT9f3Z
PodGU8TYqSjSgq9IeDu8p6by9fFb/jsKEA7mJ83KpHRQMAXdzXmdpLQKmc4zzlJ1O2/zISCV1/QT
H+ngPmtXZnZtNvdVKYuVAQVXFn427Gk+O7HmwdqDm8IJ+YQPsoAAzqqxfh4J2RBX46SNQlZWWjKQ
Vg2ykUvsB/W4x2z04r+iFpzqZpBREqCpU6WU5eEJUBYow7f5N9L+yrWCh1nXRpM8FSPelAzyK800
5HIk7+9pOaDsttekog/N0K/d23aukpOAKyIn7xu9QJqfdrdoL88mjztqjG/aWMyIko7AhMjOP9gJ
xGpoId7Ir/JcSfI1J7dzCr1d6gBDuN7R8hWwN0AcwTORS8J0dbKFBOipUB0HlW1ErDl8NG5+pslB
n+j9FLNNou47xWnCn5dtp+ulRiNj4W4AR/vse//VpFYbpTh5TSB+sYgHd9RcV+1p1BVTa9eb1LD+
fchHcPOlkYeYAMh7w1CfUfxFZ4JvQG1ETkWqv1cWDghxr4i27mZPtKnOPOBENjsO3A154ZPhAD1c
6ouv495TxHl+J0FnhKu/KKV2bADwuQFfxreZLlSHoGQThbN8RjpPi2OVtCXMExd2JNVgLyHVMmmb
tlrB2KsLx24tK93api4k0dd+88tr/pg3gOjKJ0QPMkInjwWDtn3EBwlimWu8CmSTENH+sa2jB4UF
O6M9DxRg8e1iFsVBvPgcAzFhHdiDgVxgNyiqQPxYJbCceF0Nbq1moBdPgxEr3YCH0lrwE4AF1ZKL
O1IkBs05W/rkvxGlOrc7uCfywT3i2B6ILJ+RB6IfrhFSE/dkrXRci9S4KsgKoxPzHkbHdo0ZzVD/
69/oTMdFKj8MoEwXZDLuJf0bQivwtmh0EMy2aLuWEe1idDSOloYiC9qFL6jJGmD9sOEYxyByNkkq
iFlkWodGwvYxE74ip3ZDZiH0870dcNE9RkUX9KxS/gzxoJ2kAN0R7tSne1veu8nsca6N1PTqplNf
Bpqfg2KytXDo4pYC43plqy4AxxUGA/B6KbnTISRYVJTzY3gzQvGRE+zA3HYAGluztZ/PnGxWQE5S
12nTwYf9/N9WGM+C0obHFpCy9S8aubBeTY5b/3Tr7uOQN2PBR9ltsl7mh2adayDrs4ie3x3giyjq
eViWMB7MLq3ob4exX28ctcVU7WcUHHqfjGPoo+cA/Iyz8ZFJRh0xneQefdH/KSv1d5LRfo1MGP/E
XAhrHkFvKMrb+itgv0T9MLh/AyD9FkZekfx6xGd31d/w2v1/FWBaECKNhb8B7ISUZUy/BHT/8IVa
0a1u1F3KbZ7AR+ULst20Uol7epEKiicF5G2UmeYJOa5worghqow1IxLq2xWSo0WOHo4zVeD1529P
XXXZM4EHAJxyw/SzpKRhqN9JPpLOHi4r5BnhUgxrgGydaGyGe/3Ji4MM3JR4kEweuhy0NUgFEdTf
MYCAmjJeAjb0JTCAlBtEHpHodrL19TENOAs1sK9bC+A+J4PmOzOMoYlmKOqKmWY+5nu1gcMr3BtH
0xIFS4GGG3OhLyjm7Pt+wozLoQAlyGsf1rDKqotm1WeXA0TK/PMNxwMXqFkPosJ8Jd6yAeaC5SBw
7XTyOJo6jfCpFa00VZO2KQ+/SB5o3T8qMF2EhvvV/22cX7N81NKeh0KoF6uSuikJ5zOLTiM4FTTt
tHC/A5YWtUWnvIF7B0rrjSXSF/MzVG8vS/EXfxHi/Nv4cQ1iXhNiLGnw4NjF3WgRx4orogjyL2Su
4tV0Dpax88F5hVp8gB//kLa5RNtfn1cp6B8VXLgNm/WFj3naE/08BGKUDHZRc8mhr/fVH2spJCgU
8LjcH+XluR3Pc+Wpw65Kw881b5/BY2Z4h9ehb4XSPB/LYmekTpslN0oddQEVeAakjvzpCd1VBnb1
ytLsOqrnKRwYIuaqmDB8klj42twEumI9Ey5OULyxlzlHP5Wufv7epJxtWk5A1WQjAlvoYck3cbsP
hWKI2+w2hebP7p5GZv0JLmwEijpDgs0Rz1P4wOwNPp4X1ljbMUk5Y8ZTfA87/waV2L6zJmG1t6/t
I1vxd5ixUqGVkgzFRBnsD1rsAkOhFF28VbBFkGoa8xYCnuoJKBH79nUmtdSkb/hHcgqT7Fr4oS5m
5m/6J8FCMidKFE1a/9I/rrc7PDYFO7AAx0NO6E7hITenqUc41BptRbcHnMqhUA6xp0F9KZHiyUb2
jT0SRd1LbhvrQGLGx9QNePItZIL4WmZU30u68WqP3rtvhcTVrUBZdPD3sx3QN9d7vonH19ZJEAEU
7pVyZ7XQYhuWBBbX6DRzVxmshf5/KDfZs2N+zHfrug+5+GGQ2qzGbZUl9rZwlJ0N5Q2vHQ4ko1N2
wxT42grEySdBEjtokM0uGlBsLDS82YC6fXgMGndi6I4IOjKqjiQbGldAMeB8ACUIsaFtOCXtuvUs
PktNRS2kI2DnlcDkQ42KCIpb/3f4niClGtSHlOpyw5rPtL2Jmfm9JMT+1GaogbiadeGT0czfTzko
6aDm11ieZchyhw+UIWsHv4y7HBffjSAbJfvDtAN7Xr40To6tsSvmUlkwyd1PXCxSDm597by6U/D4
iPOLee7z/yWSmG0iqn8G9ukpzZ/cVMNybvP0XkBoZerXqKZKVU/sH8LmVF/WfpNZs1b/0IFAKQTI
OuNPrt9GSdbky7odGIMZHALpHWyb9k71vyclGskjqmlUeua5xR7jyG3k2MuCXqLZiBXsLfi0kWZV
FPERLZq3eEPEPdNf5TncJi7/fPENzu+9LB/CNtvXAIfoDSeIihmkzEHhNnYjevZBgb1D6lE9TdXG
/M+pVbmU/AA+tK7rexcWNg+Bq/oHJQtAhpqeDixiBYBdiTiLynb6EUEo0Aux93CLl2P3UhITwnIV
0gvnlHkSbyRFVejwVAAF0zBamFDCAX/Ve+5/V64+vs3z0Uno4RzkjiVeX97ZaV6P3MoI8OY9ksGp
JIE/4Kddct762A0ZUGeZJGG+nppMHNhtB0lAMrfhvhXejjT2ojAw/vxrfqTzjYobi9rDCKDN2y/z
JJ1w4BcfJSsVQ6ZWBsOnnUyc3WvLfhEN2ycGB2/Ib9cYzsYsi1suVJqf9kzywvSIf9Bmmnl/7ERv
pyIs1VvJMq44w51b0wFStaYN1vfgz0J9xRFp8JGSElasBBFlEcJ9eN6O8lsu6rRPvHImAhCfHbJq
0Z/zrVDVyhtSDmYI7nJ4xOnLjJFbsFmgGpT+3RgXIuGZWtroii9/ehOie85wlM5S8tFj7aNh7b4v
Lipf7qasi1W6nelp9cYWpkhqWMblX563BO5B21isW93mN5h4hpIfljCKneZqqaWLRKS1Re5I2b3S
LsezxoZqh+bghpc2mFnH0OPGf2ftol3DLhcF8blVpMXMZCMPqsKq4zNwnJdqQ+kyxEaWlb3j96qU
Qc+CGSwn0OpE/qPPGuJAhDIqpOE3xqGzyL/83uHHs4iySBUtrSt/O1QOl8RHrN9BCw6q4cuGj4An
a1LWFfD7JcGwRKM/vDtYQNCs/UuJ1rn8gNdi0+U0XeN72c9/TaIY8l5oa2wWvfDmAiaRCyUA+UT0
Xb3w7q2RiC7TthJTqmfMpwCkrqFsJ3097fpX/8rkprJ+uq67Rndm/bw4BI5xkb6/oQqdCsqGaqyw
ulFj67j95JJ5s+YQDI3RNh427si8xIQgudxkQY4IvrW/Ynm024X4Is5O/ej3tcCPi7mq4KzBLvwf
XRtln+x3aMlQlXwUwuBIzEOk3JYN/iSzlJuPZYkzTWw8II8gcXlI34PN+x9OheH2EUL3F1ap24C6
8zk8XXC+UKNNXH+DRYn85SqNivMSl2V8pngqLk5tVhHX//vM5Y1tYhLCL9P81W0CM3RsT/9OEWWF
GBOBYBJEyNTFpYhm48m6u3vyMBr6sOR4i/YG4CoFiONYomBqFRrM3nGRCq2DXvkT0H55VcQ9Ti8R
gyS/34QhTcmNc36H9NnzBCT9PYMdumABaFsI85/pdYdVnd7fDNyDRh1Y8BsL/phRyRTB9q/uFPM8
UeXbb9zVRnjQCYP4srbcvIiVUUMeD7qNnHsaxYJgXQGQKzSevEKJfKDCRpNe5FwWSu/AcUea665b
ARQ+JEz1iicF5IfmI320nEXfOZbD1SxDAAd8OEOZSFEAtv5gX9bsuySTQ6two77Dw/lc5UExjU7I
/OTN1UJ5I8iB/NUJdZIAsCPyFiOFfFtozhA+6ekABYlrtUL6wg5/06iownzaz9eYjenC994Fvmfk
Ij9xDydQdaXZ3LfPgXiExoKn10cY3U1oSSxyAHs5oCZyRae+mCLcsWST9wcLo4ffFUjEljwE+WPS
tJoc88ZAvrtPOQeYM0e/ARV2SY5xMN8d97d+dh+igqhE4iAbxPbridHdiNS46aT2ueSoLhHPpr2g
EQcc4RihSQh+Ls+5wyXR2YcnicunogggobNj+D2nbiu6AijYP63deP1o/sRgGqQUbnDraFvcQIoR
0UxUCd5hhzhK2GDFj0WQ2JCuXif9l/blgFaGxTLTRAgU+AviDA21JXRf9OqUHb1EOxq/50DL+3oe
RNZfLUoHXsZQ1RyM22n8ssb1uQWp2NGnVX+n3YnH//svPGSpJcSBHz//YnoYmcOrlkiDQNyvpYQi
xiiu8qdJTNr12eruNrmF49I20XG/TCpa9UMzKPpTqlDnvfe0XnP6Xr8OnhF4xblhB6WcLHk33soL
GKGpLXbc6SwqVCXhL96OjU4UiGrzXi/a/xDpCjP70dpRcUi2xOpI6w2iroWqvXRDvoANfKFczi3D
mG+kHXD29Tu3ur5V9q3e5UXiVrVxo3pe7uUn4J8dk31XSfFqcAhyyCnjUwWYEi82YUqRGAVVb2Fj
mSOrzZ4CcJ6jIgwCq+nInCCqNFRpHApkEFqq9pg218wWrxD3WBuomWaTy4SwSLOIbB+MQZlYUoc8
3EzJEuU4s0U4R3ySCR6Ohn/U9kTDE7N3x6DLI+sF6mm0q8/I1lZen4ZYbW4X9X7Z4Ze5RdQ80ANS
jRWPobR2tQrsmvQOw6T+fJtv9v8cylaGhs4YpjMnO6QCXbJdMXyopPWpkBb/3muYtn0hPfMmjCIX
3PRfKLg5R9ZVW/bx9qD91CNZRLr3Y3TwOBNh7fDd1Biskvduq9dmEzWDW41hG3x4qTPuvHI7rHAp
q9wExEBBQOE0t1NulDbWuB+WKh9mUkY4V9HkFHeMHmYGWdLMsrQ+yLmFg5eD9cM3TzEv/XDTAyXl
J808RUEawYF35VXxose0zHgwRgFtiH0/ZI6Wdn0vCiJBtctdXbzMJMg9r9dmb3S+ebx6QOxnL+hD
61OMEXkFOQLAQsV0f4B1qNBH7l716iyFjm6oE/4AaFNM5He6lcyrzxXymv6Sm5+A4hHMnN71WKV7
q1eJ0qQFl8pU6Pn2nZkItosSX8b9HNpxHpeoLxI1vS9FIOlM1jOp9yI5wG5ed2qSjExCLqvvQdxa
LXoFhkrJK0kg9RoPz/FtBV6o5hWO+GlquzDtfD1zX6oGvLg+lOa4EVOiUosM6TpYjeOpkxd6F0Qo
OESLVcyhdSy3beYSV6DMw1+pkN+DWK7SYlcA9eQelZjK3wDp7X5lArEEm52X5s2xYi2BErrSyWKb
r6n5meMqcnx5pWBaemBS4H3LGGzq7kdwk9RU1N/Cfs0LK7HpLayMwijNtmSwObE+Hc8UtwoxvRCf
v5rjudqh2LQ2jDd5XhCkWPeFh2ad1z2a6iP0h4CE1ca0EIjw8YEKEl5ItOlWdeIkzVs+mu9HcTec
K3WhLEtBQwBW9PvZ5vjxonkkiPBU5NEK1bdy22QsfjzQZPn8IB3S2cQZ4k10aLlit9Wt27m6rVRs
W86DS8o+0NJz9RvCCD18xanXHtcVJLd8GXxLkn1yTvyFLg5B2NT2HYGh3EkG1LrR4IljLmaIjE+0
DMLa3SLLeYLYSJNg31MXAYvUiiQNZ13vvaN1mjGpvGmXCcTIkzPLbokkepyx5qcDaibukOOMv8C+
aBOueLQ4h/hHQD+WmSGFZjCyQXuDNtkgE8L0gk1i9HXs8Kz4y98d5T9VOlyy/iwO1LJdt79gFU9w
XsZxT5Adz2Fgrh5eUgxfVFjLANjg5fb5oaD0JYQeatbtgbW2FBz3Uz76Ila768X2GPjbEy2e/+UP
mj4kszn6bNWaaFM0Aj++bCcl0oeTBE3ga1RaZZ83PSG/FYJGzw6seK7pkY0v/wPYqX+TJxCrMxEn
K4xo0WFQ3YBNrUPpaXlqGEKJ6k9jkurnngbD9k6KiK9jXjbN4cQACzvKDW2mYEZwy8wi3JRgsK4b
QbGyFWTjid8foMM6T+DPl+Sw1og+wV3md5vEpcJMyZRba/fAQhlq5GFiI1j8zxjjPGKqHLtqB3Ql
A3hKmx2C/PN+VZTv0wHw8BS27rXoxZB6iyfUfs3hc8ansWLneWgORnmRFb2jC2aIk6LNtwPbo2ko
/mQ4U7CNsk6W3PaDljSC08z/Snfw0v+MTQw4IXnm0mWgsMtNizy5PZ4qWrCb2CI9D+x8sHNtup98
viWAEqJM8j4As0zYfoZIPTeeF3M9pzNlIC9euglalRTr1PH2WJddDj7mD204Oy5FuvsXs3y/m2md
5SSVk8pS9Zfk6NuVPTuB/VojlwfCO3feUrhhy4A+7vha01neF6EfF3zINj+QeSldiFwkdcIrFsXG
fCVDeBKIwUg0eLzKV5kSMpgbzwMnbSFIj3ndloh2nICnOejpR3CWpU5YyXzPcHeB2iY/JG7AVNMh
sCYFbvG7jbc757o7qYEZQ7wp6PScB3ik0GqD/4tMDK0oTTzIOvNPBt8fNI3zNMvtxVDPlfLx6j72
Jn8DBVGkWWd7Q084v1w+zU7s+MJnPUn8E9XL3DY/HM3pTh5Ayfvt8Shca/GccpXZaVqXBQ+mVfWO
/Js897gwhAe6/BO0RbuKp9F4mas0fStx3lxGCxAB+nv2W/UOUPQylsw0krn4UMRUMY5o46YttwOO
rsd27ulX0rqHhJYDvJEN3mXTxmahAGvi8O8hj/RkaSnNvW2hBwmylDqNrpRCbYqncBph9KH1CdTX
UXead5/FGTojrlrdLN2JsLDnZNRfvsLqUrN53HjMn/JO+x8Gbsc+W/N1/lpsKEUuo07CS7JfI+06
KQeWLzyL6VPAzVgN3pwADoSgig9Ua6g+JO8zkf3BMuDrSGH+7HBpsXBY3Us+7f2ae9bx3Mo55JEy
Z7TSUeBhwubDhBlMPSSkwCLO3fiW6z5K/JT4jMVFKITlErK/CZFnm7jcAP2ut6Zsgesf8YUcf2o9
xZ8aSuM+RlfulREZ+bSK00cNtMe8antodtPB1hErz9QrE6zVyo9gl2IXcwgjSU/SuclDqX8tnj+K
fDhmAcXdZwMDyjHNiCvI1XnAfCS9SQ1W8i1HN2bdBXMthPyow+hxv+X6yAQWseRdSvSzsfHUCpLk
kmPSzBKt265LTRMrnXcTlJnaYIJPUtuBYUisWXwU1dfUs0M2ARRDFi3HlOm/ACmrS3rYO2pU9lF0
GUVVMsyQCBmTQYLpgLvARHUrEgGtjIZqV8DiviXKSpbc8aa/rFeNfJVBL8pyMgUQH3RO9hDncnzs
rF9BHSoFFdJAgqAekfGAzRUOpxOMEA1jOfZg/g1Xfmajx9SKZM9jgrR3gJppMweUkkjtvD9Sj7Py
EJ4zlvQ1NY2wwskvQo2x0LysXPFVln2pXL5U3kpEoy29Kv3NNQ24NvpJ4OQ0liUIXrwTy5jyRNd5
uO5q3c3t0/WpXwKhj+Ka6UfI93nn/b3BrZPEM3E0m6s19nRo8wQnmi8dOE9w/eGQX8kZz8VSWAEp
JlegrOc+/LNuB8AtC8hlp9FFA/7WeLlTucQoAQHfM0lRnICpGAevyqRdXv4UBcUyjc71RMijgn6G
tEj4v+Xr6pg/SyIRK4+HYAaW3trGsghxFOYhMlCqN5+iXoKEmUalOUN5Ygcl9kNOWoiZ/899S4Eg
761Q99vM+MziCKV5tvbgzT+PAduwgy9BCEr+WttFhncaEvLp7CLCdxxzU1d5ibFEFl7b1gqvoRSf
NsGFA0Hq9P+gSpkxhxQUSOAmrXOQJw0t/9iz5e0Bose6hxZ5ri1b2azjaHSfrlWvJTH58I2Weolr
m8UPC54wy40xKKnB0uJ2zPNm9sanz6SGi37XCmLy5q0ZFbFd+OKxh4NH6Nucag9BaKm5eeoWgYVr
Xsd/in0v4a2xbwDuKDazRpBgZlVFR/FzpyRF/FmElz3qj2Khbd5KhTkW+kTV72j7BYArSvksofCV
Cd5ncO8z5Dg95uf07UDCEzSy9gV1r7u12cRiXIHxzzA1F7NHNI63acysaq1CkpEf+IMa55Z3ai7d
quFemOgS/NZZh4HSSD4/NuZQ1CmKUCxsyX5tS+mm3Y9P5Pr3UEVOQoFbGvqjzVZlssij7sXNLsT9
kDOJ1sxFQIJfxSMKOJ+EsojWuphOm7sjpM6kjC4wSnOSv6vdz3ovkggzlOlhG1Ec2jtdqrDp2Wg8
TSmrCM2/FsTkKdGwIDQJJfL18ztvvC2dBx5h8KXkU9z28myHVEHxogziBUzlmmpqjsVPaZBPCQz8
mx9y9E6PDsCxhHHbXF1vxyXIbnkaTS8HhsorDiQyV+Wcdf/bqUuKERcUq2wjSHQOfJxVgpX75yeh
sZaXfFUchu7hJfLHeddmMUYfnCKiCpXbPnGLNfyM5/TPURlSMT4DcFrAiulleWAwFxoo5gkLBQDY
R2lA5nTZfHTuaGV3CQooAR2O1osjErWNbJx8ptSdV/8X5mzNGesM88AL6NCB7hJEDlYMT5+88AXF
JuWecGd14iTP4V39ZyiOWe+lW6pGpLhJs/XKOEKXnoVQRZkmdkrbvTc3+T1Il3a82jFx9dvz1e4/
GAIlPT3w3eilgfrGyDQgMRgCUYR7ZyG5vo/jS6Wn+ZnHhzjCxoTN6TbVmPQt0X/uDJS01VpKbxjO
s6RIkONmCR8W9J7QxKOnxlxx/5oLqiMqvlotylM6ssOjlC20mopPMTHbHmdvGAVn+2LcX9SPXufU
5ABrBRUgHqS9XOxXAVO9CWcU2a8rvZS3MYzjke7SOElmJ19K2ZCOnZp5UxYadDeu9Db7xGK88rEI
s/0Q0rklLnuOZ3u3hAuXzxmH7GELClCDmX21IGJGsRaVVCZm8VRDr1GpAcQq1Z5rvjI1ByDfwTf+
ZIzMgKcuRSk7SkkSPyWA1j9Xrx5DD/NUPKfydjcXIjclhwM2vPIHU3nertl9ziMIRtHgBn18xhyZ
U0WAe9uydoWBRSWC+IjWwgmfX0Go12K0AOufTcb87Vvw4cqxnnj6L+6OaLC8+48y83H+BSiyUQuf
Y8g+9TvZEwFegab7wNKD0qotW8BS3NBWz/5MF7o+G+/Yxt+vidVkxWoKXWeMfnZxxJwR0mg/5lwe
2yj5xVbaV5AzVRDfQtyMPYeEhy/O8wv3W89Ar4yp8r5YmARNcto9jC6v7+dUqh5f21q1lx0pCvxj
SX3UXEJaxBQiT7zaTtHceN5KI5tyL6q0Clrgp3y2u8w6c35/drj0jMNpSWMnDTrQaOM0kL7gGMkM
wo66aCMJsGSiTu8UYtm7syAqs6wqbnUpKVCPLAwPvz57+dopef59S8IF2ZlljXTaByJOwK0JRwgj
rXUn29ur7ma+p+nCwlVaWmcO8Wtgx4cEI0nfdZeHVIxRFOzGcw8RAcjMSzYgqsb7+BJQfnicjEy1
z0B3xFkpH+XWqyaqKEuNFX/H+q+LURhvGdt5digp6zT4WLjvAsA608TL0EQ5PvJgN8DYFLbSFe7J
UJRtfa55lbPTvsgVpn++4sIMicJWo/J8jcTYUwUnHKKi77wS/+1zKCjwQ0fUig9m+3El4LZQkYqK
S723MYDlcZtYeMl3jIqesKA9tvUIXwB0SrEeaPEWv2L2ILAAzgFsA5wd3nmNn3/ELjmp3g6gPoZh
iGjBunVf6/59ccU0nUHMBGdM5RDnx5YTIY9PcOh4gaGY1f8KvLqkqJY+Dv+Ph6MltT89+hkfTULM
/iCVGwt7FiG6tJX7AmTWtV1Ob1JXfc7le5ZOVESYJ/d9IsbdyQe+NfuNymENwA8RgLpXuEz33S+9
5Msdi8mo/jgMWkD0MoFsFncgDxbd/Y28IfP1y3IE578YGZnTZIXQT3Z/iL8AQ0lnIFY43jV0RW+h
ipaia3FlBZDvS1eoDuLvT7fdd2PQ2wWtdep1nBvyUL1pr78mFOqs01uXfHX85qnu3DccesZwKcdJ
kh1rOE89Mjdts9i96W3nrEv74x9mTHHItP+QbFhuWPZJeNVtlZFwOdn2Cg1TFo6OVdCpRsVqh36q
WG//rDBVqaj5gcvBDVNw3HQNzl4HMCj0hFQgGkF9lxGbDWHb2VDPgkz1XBqY4zhhODPDbmv1b+dV
yMY9EXOQkE9S8KEQkAF0njVnMCsODe48lhmjBaFkDj4eQsUw94pPiECciHHR0RsQtogWtJrjo/2M
/RxkG/zLqjnLVIkldMUZ5gGhPoJ5RSH8yZxaMC3Z9BXuYz3SBXgOMEk+ilYPikGdtR54ddEddwhx
Qu2Iltr+X7WXoZKVLn4aAXNDEaywvC/yrpy5mRrIUPSdgDm70PzT70I38oRhDqmNKpMfq73OvvDo
mNyDvyLYvXd0hTa8oWMMk9pxVOILFZQ/ahmrxBNFiiwxT822vBXUy2M2z+0okiELUclS1ujlQoMQ
4ZAnnEpTFP4Wpdh07/5fbbQ9ePX4JO4zjwlXO3ebQAlh+awd3tuXYVJi3Kphno0NKEpB98zcCF2j
B4VffdHyUxBrECQO+H2J2WmUT1mqj5du0iMrPCXgqD/tpCZeDd1K/fiNzHUiJlaC1uAzN5+qyUv7
jFfxDXz8zPXlFoIihzL4QdPUcTdcLLWrl/GQBexrtHsdOI+Dh7O0JhT3ocy5rRPXTJxT7exdwXAB
4QaRAbszWcwS4ZXwxNrLXw8yb4B0WkYkoq4SCUqC2zHkolSO4IUbXUa6ZLSo3lzrk7QaZlj4lnPu
sWqG0ftel8k0fPiupFHl1SGNPztNfzlWwFe3yn1XSYPfWA4KmyA1//LO76Ylyq+CgGT3+K46K8Xg
5EmG7aEEyZt0rFGHRkiSRb7UfZJ8Qxv7Di/7GPl9H3E8Fg1SfMdcufGmt217Q9/WO1JYp5SpkVaI
y5VJw7aVwWLuFE8jeLT4XXmPRN1MIS1hoTVgUInzG8Kc+B0VN+qOhlKmtED0ZOPwR5beEmpLWo4T
1pGmoLwEqRaAGIu9dY73OXIPpT+MTYwTdzPp4426g32Ba16D84zeqb2GoxG63txD1hkb68lAp/Ey
7HYyqMF+v9tABtZoYOiDzVqQkYISxigBJpfnbo5q0j+Q6yWZ6igdxwOiiYFSEMBJ81WWVqaJUxY2
1u7HPVykkSl5ophq4UOVp4xILAwTfhDGna1Obs5Ayx6xzCsZr5wYBdcGSa5CE668sU1W5ID47SmZ
u5ZCf8cWLbx1wOWaF3Jx1hBXkyKorSwcRB8dnh6ILnPBIy6reVyp3gEjBkokIGY5TDLzoPBLdGUQ
r6GfNEh8/TOLQbMItpmV+FhUaaNUxzymI2xX49nmk7oHXdwPMt1SEBWtA53BzsGZLzLLY88JLC9h
fgxxQZ9WyWy54lYiYaWesy+kXyr7nU6B5WSZ+dGsOcEU/jQAWZjFfpHgwu03HgHxYzXb/wZ9UuSO
RCsjO2VKSbBtKiFGlzrqP24lg2kkgBNLK8lkIG3DugHe/NG5XhABCbu4lqqWMvClcuI3tz6LTOzM
2GWJ0d7knL+4wY/Los4sspfnqI0jNZdefxo36P/gCfvWkkYY0PN1t8uHY0kgnGUSW/+EX3qm8Whf
Sovg4dFMoFHIIeKY2hkubERThL2jLeRbfV/R3+xD6NqCbB7HJp3TUTr50gckZ8Bp9Ga2n650pXKi
KKc885f0yQXwnPNuT9MxJV1Nv/mQPwzYPOmfIdNTxs4sbID1voSL/8dSbj9RrJhdsVo2vZ5ZyCVD
/UuNfic9OCKtRcaiLIFYVvYJy0HkmYvyeV4X10tvuvBD5EwtXWF106lgkfGry6vFIeAfXLISut49
VOFb6/dP6g+vaKGXdEEj1hDxPow6kPDgeKDz4AVmZTRzygXmqUdprtw6mNEcIElvZ1BWiXgdeKK0
dxU4hli0PsK+82WR3zT+QH66xoUlFA8RGh7ioi3oK2VkVpthOOh0ov+0htv980csADsc72pozhZ1
uvvDfyMCkNhx1U03hOyEbx9YG9AT4Gazae4RfJuHhUnnv84WUXWIowL6bA8BqeJczNhuU+4oOt2B
0ABSy0UilOgG9HzqwdtcMeavirYF2nrDbKnySeb3jS7un/Y/d+9aQ/GXpT0viSBhmdcNu1282rKG
7OiYFdz8xsZLCRPc3Cvvboz2v2+Q9Wv6rBQexBGMk2h7ADhm/YqtOB2JoossGjpsfUeiZccy1Lla
FQusS3fJq0QC9jrsZFM3cjC48rAJQ1DSOzs8MlW79IqLDZJXN/xRYXiwqj2oD1h1IFc1yjxJvfsw
/Dn1rItfbPY/Q+n2DgVTDy/7s3wgr1bQPvJJs/Eq3lykXk31JM9fm7Yuo0zf9SZLUGCRmlqGurIg
Are7+irQ7hDLxX/nn+g+rESN2LOvoqNRGVKJj0EoIhZjKXO75o7O4y2sbPaKAsgHRD7irJWGTaC4
BEGb4RmOcpc/jGLNoZJJFP0wJmOpU4o4V4pH0Gikk0JJee0MrlSvF7qVYvTbqdkh3hhezUOouflJ
PSvrsH1KCnFUsgyNA1YIBXYsQrY2SGUdg9NY5du1tvxwT5EtAOD7PLTqHxpZsKd22b9j3NwS5AMz
NUelI14wOHOy3SQzQO0ihlhojiziR2kZADBXvFUPQPrYFh1DqQADmlAvdfaSNi7WFWL4s8irAr0Y
RtUQq/9TqpcuqlqHoJrbY6KT7HQQ/LapPrwe+rF88goRhg6ELFuJBKsQ/jRTmRgs32RouiGc2MKQ
frKnLBQJR17BFulDrhIkdyuMSlh3N/V9idFxmIF61lijvWJoGtPu1UmeHjGgIOa4+MJguQzf9Ykk
hrwK1hP5gomwMdr5QIbLZxoUCWMamCjvTVbXQ/+4ckXLMO/DFVrggKpPTZnnwiEuWgSZhXN/EhQx
F4zRu26BECfXtA3RS+ACfIaxkjI7Uu9J7UjipWIyv7Dcnjk8P3CdYKWpGNwrqGCgmxi/PxW2z153
k3eOGuyNNFgOIZ8VTAzCns5rCkWbhOsxMyXzIqa1qy8HBNOWuCJ96XMZwLlYxcSCO/pyqcPisnJ9
5zy99rY6stgzNSLFeOnbuYWUkEUxW+T0vJSzbblPPMTdmZ42C6sfIvrwORONzMbyfdhJvUBNA2H2
6Pz0rUx05CAFmgLX5QUSfljbU/EZsBmcgYM1Sn9WsQMgjuvJwB0bOwNYHsrWKMHUBOyPwDDWwbYc
y4+8jTO85WpM8KvVDP6gjW8s8srH+d5Qx2oISg3Gu88IxqQ/H9rgERLbf1JZyHDOqslZ803yliI0
JqyOGcn1OX9Tp9S9pDIn/gGMjUBEm0zV3EOSgswIOXmBeNEQd55K/52F9bMIJk1TPSfIdceIjXDb
w3qVJN3SZr0MltAjiEVqU1k7iyUGfeSz4nq6iL6V94bPsros/8d07uIhzV/fywH947hISpMWu1X6
lWg6KQvs4aoQS3Fod6QdGove2oa779NKuW6tA/YwIMWr1IUgfGxThakQd62b8q9kLckGqHA8lEV9
OgC3EuK0tzNjeThinIZ95KDUCei6IX0MSfUmoGfK6nJMKyIWMHm+qdK0IU5ze/R74GZbUfJXgFT+
zItH0rzIDmwT3Wu05eOAzTSWPMa0dj/vo6J2xCFkgqZU8k3aupjCGY9Qg2VWWu7xlVZsxvvcFgQ9
Ojaw8mw9kd5ZGmGjmze/hcNdWZkYRwBrjuBbsNLtQSiYo2Cqqyyr3+tnlwz5VnmHGFNLXe9++nCA
qHJIGTIOrcadrF5NQZGPUbsgsI1xT8ANWikaRkHSY+23Pm0HyuIzOt4Ue8GLH0YGgTYf70YVYgcx
TTGBUHLxkNm6NtII1NncKsLS8Rdg/paqFIy8d7Pxh2zYq8V3+uek/z0kTU3qBaqQklugXrCCsA8D
yzQJ0tTQPvYuiMuTWlgpqcTZPDNjJlxU273bBSbxEAhuucALEp1FAMg76UI92KdcfNiqZbBFSTbM
6istBuxZ/xRuEvTEVSgWshrv67ud5v3Vv3Q4UKH/Db54Oec49MarwLJfFJsStsePBlAawqIE2/yk
6mSHue+7YPM7cYpX+TTpHy/rY9Ge9m+un8Px+wnAw82jg3pvgQ17CMgF0XA47ALd5Xzj3++7Pj8H
KW35GPMM59rYYBEK7uOYAMEAitW6heb+OD8RK5tRU1gVyb+gtaQTx2spCmFtird6d4xnuDg45RF9
vYtcrKD2zgiTMQcsZXAfS0cFH1hw/Hd6C4AWVAvRVxsQYon4R07NlrjcH1gcY1F/w9JtQSWKAwph
rL0C93xptKM4ZaGz0/hFZksIWoo1B18rXKKcKd9XvwluOQT8kiSYlcq5seu1TeGO8PduV72x2wqE
ug7FJQWXyEpdKeCpNbE5Agg+dr6+BnyKsrU24NW9/LvysRCBnRlwV+3ft3BlkfsjJI5Wrqq+gKLl
WGZmULTw01xCM+w6+GdG450zoRBaLCldvsxvayaLfFWhtZ6/ExkvxQo9Ui8OO3l2yWhwmbg1mhad
+yrvOczmKxqfKP+ASEdb/G2snmyjOEU3uXyanNUxfo148TCdgeei3ituamEQJATTA2Y0sBdaiynl
b4yRQxMDqkYCiLw/myRp55VOxfChPBV4Rmjualw/EO+p2htG16QElacHtzxG2ngF16Zmou8Q1ykI
pGk3HZTRblxAE+Z7Gg3Hnye2nqOBpft6uERDoYlYNsM4nj3guiU4O4Z9Yy9go+ZjikqcSBMrcqhN
xccoXt8N+zffn7n1bwWj33OMNd3LdssSfUDGGMBZuWK478P7y/89S2Y/Zd3npxZjnQQfTQJyxZt5
vNktLRMkbYR7N2xsP3D90JipGEbw3l4PJgfmEKJToLEUYpkdMnz1XM7BzCXogK3kV/zFlZsHXvJd
lxapp9WNuf2aGAHxDzh8VCQQaf8fjWpdNyK2GDQmezuyxWb/LmCG8U19Iyf65iO/defSzIXa/6WQ
PqUaWeZpaIKjZsGt1t29LeQQIQYbTE+WRMAcTyTvO97pG8yc7mYjkLnioAxLtVRjOtfuujaQkegF
uLkxsPrk31fXfEpD3j95DTNVokh8RHAJNETq2psw0h9qs+2hD62/yq7tdQTNGlEkGV01QGwsvilL
WkUGIf2YbxijPYMJNT6XZBJqoHS1cN5NCUJrVMQ5HRNJuAKB5sWAofwvhtXY9NDEyutWFamqfIIa
Vzcp9C1ls6uEa9gNrXczVtgnZziahWIxfbzpMSeAWhnbibAaB5PvQZHxlgSoQl2uF36TxNTjElgR
TqJYQxC78HrXiR5553Nd6/78x3rh2amR694Ak2Dgby1um/Jy0Ev/IxurREv5QZiB17VhF4miFWzq
jfLN6xbMbK8FMIMbsuxyjcZ1LROQTWmpAGm09CtAWuh3mZPVswlV6Fg0YRiZoLY43N5DK86gMEUu
+UYoApZUWaZTNJVTHp6ix5Ucu126KEnOnKNN0OSY3FWnyLxNt5UcqE2Q8S47hG63cyZ9KQvTzmDh
MzwCAjmza9BY/8A5UOK++GDnPcY7WP+8hw3o+oc8u7qwT4jTdlKGBx0c48ZFZYsXJglu63gFr/iw
PDufRz313Gc0Yfol7ced4dEEJa1cK0KLLwepwCIaZUkBz54daXyTU3x4VOHyueVauFkAqN1aHu21
n1ulcpS0T/RfihhNjuC9tGs6Cd1yCIvMplwBeqYUATwm7G9Td6+M9JSYOynmYUdrur0c3KXfZP0m
bIxFOxj2t1buCE91YjgjZJcofBvoUQnOmOWzqFKlcRAzr8VxKe/uEMAIoTUzuB8hH39hPrtc2Mki
Sn8qS+L5cvcaCtF3uud9QhP3zbGdRJbsMcq4wgQ4kSG4Civ6/J7YEbct1xTYCop4cxngrzdVwhTq
870Lw7NMv+B/jN4MwSZM46VgPs38QDe7zdAYTPDcRpQpq3MlTrz0oVUC78YG5G4kr7GPeBi512aV
8/chUkebzlmzZ5hcliWML5bChEftm6FH9SBNwwDppqMRQlSyQXe2RNb2s5rkJYUdCu0INOE8NW/G
8w/gEcMVo8a0jWRQLbG8aC0WIf8F8IAcDenYmr0kGrJtocpdBMaMC4pfYNyrz66wGAnLSWZeG6k0
FdIyvavB4lLsLG2SF7gFBeWEHKV6Evk3f1378ijA0N0JGaBqnMC5pKGtbDfcpZNr9JCo3fZsa6v8
u1CoTfNye0DYKvc4CygkS6+ph2ahQzzcyEiWL2j+kzmaK9JfNWzzxwDum9in+HE8s3g0VT9pmw1u
8W8FFp3R297rGb+BDGRsYvE8RFRWBzk2y3pCxf+lVszbB/i8bU+7FPRrJxn7KNGQmY7Ka0qt8Td+
fW/1H+efoNnHkwpVrOCErrMUYI7IzE93RjcT7AvfiImMW1nnie2lAV+1kRoQFNuHo63ONyLRB8X9
2rJJxsI8b62/j+r3ov34LwB+8U0rGe34a0SCBf5/xD4ekveev5rk9z8fhswtVyMNHpWzt3IEqC3M
pv4y8cppHXoc21RXPqUJtlPE4jpxDxO/GJOMIlHxVkh1pn2AFR0SI+Ve0m76xx2a+AfiolqXpXCK
RlStnCsIyqizNLgZCm0rAJ/MKdRrrBTARzk/G276K78F3seXZqNnk5oXdaoFt3bumHVwYcnTAX3L
eb5R6ZQm3HFN0oSlMQpCT9Bks7e7FojJnTOXOmBCRf7npEakijy4yjj+IIR7eayqNjF6OU9g7GT1
M386QHdSFKsqZtMUnLNOr8Fq5Jm78usf7QeJHPeLnKHSECY297oIjZqo3VCvmfuVynFVeYN/D/1x
yDOwwb8Wc2JQ0BTkEFDqbz8TjcaoIwB4JG6/O/8CWYLtiO9sJQqupoG4dpqloMeAVtSmhAO2fd+X
d1KbGEt5o0TPRNy+4RVEuQOes480+r5tU9VM8851vTcDHATfIsvlc4adGtHc0aWjq4uefE8jDcwQ
eeCH82ate6UYkBBt5jyF8uRYPlqOjCYh4Ej2fkLNlbmxr9dJOUew6X7rjfgUSGKUSI5DMIhBQWSx
HMpjI6FVnrYkRhcKQTqAv2LYfWOhmWgKEGypqODMmQkcXVi6mBdz+SU6Ms6/qe0jRV2I/cp+55qK
2R2un6ZjvweEJIzBqoCHKjOY4cpJpx92PvTJ6bnqxQL/zA0iKrST3Q4u9WNMg2QXX5eqzrushKI0
LP5toNgICuqSHA9zafIkcdIOmoY2+o1VB52bcimqgojbHz0itoBgSvE9+Ekob4PeCmLICsCQQ7hx
fICFM7IHvsMrMoTGKl92VZUs8BtEzhqmkJU2wQtW01G/8hdR7ZNR8rb42af9+sNnsTl8MvT2htrT
nL18N72YXJXjZJ2B3NffShZ7wNp/4oXZto1AW9/vasvJN/64xRv8XRPLYOpNvHPawGdVEG/YgdXX
WebH7rw1Xs7lKkVFHsCgegGXBzO3O8oKA8pGxlrp0i/OMGAR+rnUC1Tb64U2TcO+QQRYdN1Xvo6W
YlizZD28t2FipKjwzMuD3QyYtyRiR2gbPdgICuj60YMZyVt3qWS+Hs9q90Mi4nJDUD6Qy+j2Ha1u
cuJwG3dE824fdBA2lsZDvyD+xkjaOK3frA9a1o3lYR733tOa7fd/gxpxqaBkIVwtnBCgXL/K0Or4
dCrbzMP036QOvoQv8FM8bTQuYTQBztx+8fFEuXFSeFlZab7MLmybM6cvYzfK0cRL6H47nusUHB/n
GVtKDaqOzXLp6uqg36Lh/oAKdBy2Fytbd1NOGmjxHwkQOUWdz2O29e/4pUpR+WPgUmT1zKnVBUEW
8D+ryQxoMtFvwKgSkF5IK/qD5a6TTcwef22pxjLDe8F4qPT3lAwngm2WxvwHnld1vBGjKJ9JbKSl
IomMKvTaj72+mtbVYiA0cGcPTnkMtVhN3a7BKPBNVp6VDByzvUs99NEAShil+ZWsg6l/bRziAWBm
ZW/RalXihx3/W8mO8dQDSt5FNc2bkweoA/nXiPkWeTR7SV8Ci2+6gOFkp/YxMgJ35RGm8l/UpZ6v
Ir6is7l8IH7mFg/23kMAzwzyiDsn1hqVH7YosjJNHxnL9KPLhGTrxZFeDgSYHrumm/qVjd9gy3Dn
FIS3i/aLGJTuvyUF4JrjilnOHk9WFENh5J+/tFDaUH3BmoQQ8fO5E6u9FdM+YZxtGnGATu/QANVm
DcJTNQ3xhhmEunw+AnGbI3tr+cmuYewz6ql50TBE3hGCP5GKRkC8vZ2ObRfgxEgBWt2lEyAzJbuK
dSawmqIBqs9q+kmBABzWZfotnWCSFWHTLYQjPxePiPYkt8n1mlgykifp9qundHyhg/IGkh9pJVLT
/ZcRjFUwLiYhiTe4bFm1kAkhX6szEyz2Gt1TEEVidZHZEbLJvgUjcKtNIJfXoZ7ukBjwMYZA/3nK
QnQsU7L5s1arbjlsXVhthSoSYI6ZB5cQEzMRSZY7+i+TjhJCx4qi6Nu15fH9sNM/iH7oQU4PL46u
4PEpJYSx5hhnu8duC8ayYDjk6GBOcgi+B5stfKTv/Hp3xpGg3zfpmF5WNVHDI6kjXKJ+c/QqrsyD
r2aFIO4u/dlgaOV/s9J32v+6RHZkiLMTvs+B1b03yEMeGy/4jfKLExhpkdiDDMOi0GuUrO7omZCD
ILFpzO0ryfLb/IhQ5GHgRsMD9YoFkYDmnBA6HWYJkpDBp9eAtTvlP71FARIFOUQGo7eeHoSZdNpT
SDILKwPShK5Xi34PkvWZ2CEIPb4f1/YsQG5LDhwgidTDPzynNG5l7mNfVCAGx+7tmSyMPB+SvhQq
rH37JUOPcchAQgVcZSIeoSiQFOTZ5fAYPDphGCYAXw5QVhOtp1iefX7M3eutk20JdlkSPZ8UivWx
jf8gXKY0jv0Fpn4xxrSGRpcnqIOgozt0wzCBpS118VdHjbeFAmCmUmhgSK9yl+HqqfIZA7Uun54C
Bz3H5OqCH2/7TQsU4H4VsPsEJRavBft3lqKA/wJa5c0jcbnBZdkm/e4uPZRUCU9P4k1ULVOkrtdV
XBkaedNprWWPxiW8f8+oYgoepl2uw1kAoOaTvVPkP/EwcQcsZL9WuRuuwgRa1Qg4E88mLnPDBX3N
nTpd/BYA8sotJOOhx/c/ktiwTupjLaxFyVsxPDWlk3eZiaKKPEz2niH9RuDAUq4MBstIlr6CHu+q
3onMjKlyiKZgWGKemZuvC/kSKglCP65fDQROlOtcXTRqC5hrp+TH0IULGeTv99KGAvHFDoTd1x4u
1IAjKk4N6pcTiMgcPzw4cRjns4vu/Rx7fzepCMYY2uy7+70FfGyVTLJIz56soFk5qOXUp+pYX+1r
Mgbknu+mcqsdbWhqGUURkK/LAUQz3AxYxa0VHkcnqzKbUplg7n9tgTThAqVpnhVux43QmGH4Dg6v
f4/w7daRT1JchLTuHYmc7qFUx7WCrWlgzxz5yrSLOgBPMRPx2/uNUS9iyVbtE4nI0LLnQs2xpgR7
u1mCmxkmj+/uneFIqC6vEM6vqYDdHhTgAfQAOtMuvjYivpaLoW1LNq4f1/3LwZnv+wXCmbYNRLm7
J9NQjj3GabUuOa8uYr8pWbwyvBcAkoDGjH6QCBSfVCPcSJoJeABqXBZ28qsl/SwK0J2g9v5rQiEm
0cC9JbUJ0W60DxagFQ2wYAM9LIb7gepCz+H6fn2+7xUxjt/4E7q8l6v3G9YhG5DUBU2oQ6YVj/Cs
x7X5iG5rUdEIW8i0RGRlqPHJr9ZwrtAFwU57bTeQUfoVYCxDbLAiJwMr91l9oARukOA+2Prqyz4Y
PLxR47HzXV3Sbg/5MS3H1SrlIDAev2IPtb0rW0GuzbIdqxc+peLkfVIrkUKwgZhheHcMqLf2DJsr
7IZaiqBtGrtL7Ja9A+C+ngDTqiS4LcHTprowfft6rjfJrPs+fxagUM8K1SkGNUXPUbdOQUVhC8Lj
WekN9uMNXqmHEOHcvWw/jhZt72qAgd+r9YNSha5QD+12zbw9jEuiGDOdIFhSLS38OwLUkawXJYZj
lAPA1lUBOwUr/YxBnXnPI62hNMpHMNUMtoQbBYuXNjCIKZCvxpEGKrwtbYctPeuCGGLVLkx8Oj/2
+Qe9Jkh8AZ7nbsSOhiqH7c8bPsxSY0qxW0Vlt2rP00zryzxPnpPGs3cnOIfgJbwxo9iDXzd0btnm
fI2I+t0dDTN8j8gyWdFPYY0M0CqNVLUQYG5guQSoXjATyqhxFx0u1DT/HHxjgccFCMoh91pOaTkD
FVL4drBTplmd499hXvywMYctH3vuUcyzUc2myJivGLSerAdGHiYOKGzRzhyL135gEgYO/F4Mv33X
5dmDL6IvuipmVD28d11MvyjtAE75hU0n3+Akeg+lsSIrNzyImTGjHYs1hqUh6//mvXqPq1xGuCT3
3aJcNVuAoqd1EBECKWQOis0nSeLSww0bFS+NJfK99sS6HOccR/6O3Q5RsTqbPIUJe4DfFMM3GTcx
PvrL7I/3uyDWMxsrTipqyK7rpF/kLYrPfl4GeLCFme1LYgS2v26dPYM3To3aXo4yJQiEgnJPYQCY
MrvaY79Irbw99CElWvZkP/I3pjdls6gLGHh1GdFSF2pFTaWyoq9LBw3IIAAoLbB3Y2ugiHlvDdMZ
QMr+APsj61Zp2gFHNZ1c47YEiwL0HYuzP9G3WpQvIxGnTxRkHSFcQ8YSFiOpqh8xYScz8aujWcqR
7C8WtaZ9MjDYJplwr2xm/RbI6BXh/BJDwkKgQ2ZRMxkBHZ7nCuvyJQBcYiyiHLRqv0xDFFgcWGet
XtNfAHvxAaVmZ/siTmb1pvT1rJpt/Dbqf7LLDxXk9FeUFoa2PPyQYuMTigsBzFvoA7oBX2DGahwM
3QCWASGxrdMGyACMEqZO3FQdE1NmP8R5Vbj2RqD0z9s9E+ycZWWVg+Ta54qK0NMu2S2W8MlaZ11u
anjgJTA04sfbkZwZtFLtxlOugtXiBrbj0p8fdJIeA0+XjETTW6ojqWkjoqDoUvWjHL/Fvv4xIkHE
pOCQvjOYrP0J0QqWgsChiSI1R/gCsN+KOvCKi/sVFHWRBP+ACXmbEJZs4NkMuq2uiVErf+xUVMlH
rpiHR74iTQieAbmkdPEuN83UggCf42oUo+e/wOmWdd0FwwJ7m4006BqeM7z/XEdGgsrQQq15xJl2
rVlGoZqATmMSlGKwDHfqrV48CiFhTSnGdfikgQj6461hAQni4Cm7FTy/ff3gnmIXhXzQk/83xlDY
RvpxKA8CZN8/vaae2n6gsDOObkd72edy49HomKiH/gXY8d2/WOsR28srh/uaVZsUOyQSkEuSLvJE
zwXtf6lXDsF1RNVXFQ/cO8r3X6CTE7BtX5cW9QmaIwZa6kytoTuTBEIjr9acJmRspjgqED/gwrHA
z3Cxct5hA+Px9wY7GhrcebYRg5t3Cl6P4SvdWtdr0qMSq85GuAgRst8tP5oLcs2qDySMl0++jfks
1MHKlCmSihRfhMfpQKeYRJPZEA6W6czu+51Ub0wVcYHLZIwskSdLJhU8hVg4JEQc+Mhu24t2qIet
Gmbaa3eeACzKebXJvmaOr1ySquyLtmpLGsdcntUvm6SnjBSNHegTmIg8NLbNaQAFD6GgASBB5xmV
ierf6pFxrYmCbUwKLSW8pGX+tDVPtStU893UlIOqCWbJEnIqwNkKfT+Sr9yU9MHNyaG78Tqq1t/V
kfvKje0t7Js0piN0pV92DxkIrzdiVnYyDx2rV4RxiG1mIyeBJ8Lb4irPziaGP4iZaylIynDWtsf8
wBBYft4FyILd50u4QXdAH0jSWyYwK5hs0zW0FMZ3b0LZ+JpbWgwewP7eQcU1ny9D9YSrANaP8M3O
8B0kLCNW/sjqIguVWX6I50+X10rhGx4qRJYRW4d3EddZfzZfIAzGE2DXDweoQfxEBJ3acaDMxbel
FDQzd8aBvFR1vjjUQhgtjUVQxT0D7TDoJIhaK+vtNx1VbGd6b4SmUoAXgHdaoFMnYanakAdOaTVG
nZqwZQsxT7BGom9hjMawcGyxfdEDfhyHMffjRz58ew9IKar0X2IrkQGLVnXXXZbSpOQx+qixB2U5
cQzGiTz4+Us8LsxnVSr0uuosV5qT83pMI+DpZv3kfJib73me9JZkasHxhm27PhrdBGD/AOK2AaEd
pc4paCZtIECtkODNwWMifQhJbLR1g5r/ytFHIRGDJNz4oopxt/HW27evAQDHSRGhAA30byCc1deg
798AnJ3WpTaJunWiuvxzvG8RnCTSkFdkQGcMAmnUJ7wFCG8ZN3U330fchtC28OuL9qJs+8zblNWY
D51DhY709YRK4NG80J4ugqBAS6N6zvTOqjgYwemBgtwvLofkCV1zjkyiM2/E835DntZyeJGzVZl3
BTTFlb8wHbtgUFm/0d16W74ieqX+sJNwEr7VtCICi1MFmYuxRwqAcxMT6jTkgFWX/G0hYKOJRtwy
CuC1PdOMXXoKI/QmDUMAt1caRBgTNdzFOV5Qbg33/p0RdzxcVmVazxWHFq6h2aSFlrXZgDN1DHsR
FZsdtQWrBGQ1hnDcu7iU5RGKZ5XcyP5iRKys6ip7k8nVotqiEMGlyCEO+SR30ucyAwknddosySd7
MQirDRdr/2z/6VgsgsUyG9f3FFfQ/1CPFPJ7pNcyaQdg4cwQjwx2x3xirm2EIl39VIozT/dyoVsH
yPcwGdEn5LuwNLzGkl6oetcqV3FbIPnjv23v0BXM7ct4DMW5wS/wY5hBJeF+V6H570zzgo0ZVfwZ
D9YnzE8TokAE+qPOdbCfEBq4GFQ92RbpX6bPPwYZhzDmL4/LfHt4B7FWgBTP2nBXEVQ0V6YMcZTb
k50nPcZnJSFRtRijyt/dfH0w2iSV2Uai5pYYOcSMIpS4gLg3mNrcAC6KvorU5uF6XLZkgxm9Uxhv
az8tmHEQAt05fZvNGJ/HF0CnDaZu3xHGDqvART/mlXzQrhlXKOwaSPqsCSoDrXwhmtOKv/n8cuf8
4fhjCmdm+wT6IiEzPXPWeSRHR9DB9D8fyA8jSw7lXQoFATq6aPYFn1O+/OLZf5HiOMATSsmhX+KK
tV541CLmDnebcobBZnOvgrz4m/xl09tTlqgDRK1eyovPuAWdgkNPJRw5dpZsohT03071M2mDgcWF
dlkd2E8US+gA3FcY//lYUQDN0P/f5rE08nJMrebb5/jzB6yGvpxbD+s7F0PHMyVUla8gWQN0GRBf
yyEM6oRZjrQnQWwcY77/MiowdX80L4Wdusyo2GEQVPCkoyLuFHsWqET9dZAfPQXXQ/+bSBTGiYrV
JipUvuwXi7HPKWTH3dzmrpAKK1gdRV+BJKLZvSozC3RCiTldk+TSlIBme0LDjNFkR1JZ/GonxjHe
EH3V4jXRMswZHHXLY8TjWhbVt0v8FiWKAxVnLZ91/pYQxmi1OwuVvaCEjp7GHCRll9ge+Rn4/Gcf
MOe6cTbIGloEpoKm69fb7n+gWQj5HUs7JLEZkDzgMFyFV/q6xVNnALHJ/pM73u0BfGv7Gc/0qp+c
UI63fQO4YXzK0dur3qqFeV9Nxn2kTBYYoVxVHLgoqhXgskGu7LM6bXdFWLmNSzrdyTzBOzF9AueN
fK1exe92AJkDy1Ifgoy2Pd+4fTBpzDemX84/Lvd+jP8arOHmFBC76n7V7uSccdTksslKiUfpkeMG
36c9pivPA2weplgPDubwgotgUUt4L3uudBq6wT6Kr/p+Sd1Vgu/gtmnkQaR86wof1vyoFcQPD5vY
4ITJ8V2gk5feDTfMGV9CoRkcoXg3K81XITJnMWHP9Tn8fv3sacFFwE18W8FyavDOMOnFUW+xWX1b
9tAq8MV0RD7f0EKFxdyfmpXqVjXA0DCpiNtn77joU2LETZNiTblTCc+alLHUUPiN/mvZ1XJ9kL6E
fYlHsqtkSPnjjk4YCm6o6WKEjPSJc1cfGlGEBET1TvxgEtlWR9Z2exvKSRKb/Nw9jaUmTx6xQJrJ
SE4eIvU3WSfHwQ2UrSrYWw5lFpi8vr83WTV71LwdLYjYAj7tX4HYM3ng/huXiOOYgwSN3jraFru/
8FUXEv/tS7i5ec6plFyHbIQD7RwzcwWWhja7ZoVVLih6mOlw+xTYMUCuQSolD7f5Qa+fPflUWMC8
xXv+bxXuV+nNpIS3CmrUgCBei7xRZv08gcsgdBH10dYepeKUDXWtKBWs5o4F1dZDqIPw8NxkaFuK
IqW3xGiX7ISdJ4+iRH3XSkoL2GUn1KBnbEAneZqFuTnNQYZN8OT+7MaauU+REcsUHUQXQA4Xk3Nf
qe+UlTtNgA9WaFKKPGviLXBowGpGH3bFaXfuCA2uS9k8vzJ3n4bRkB5QOtZkXmzaxB9mOejCNKiB
IHqYXV2nDYjZ3wGCNDnTN5o1SUQTyXUEdN6xFqSpvs+ics0dQzgKvBMPy6Jr3wk0IC0ELWmlmvi8
x6086Da6yByaQ37ESgbzYEAIB9tE5FlBZc9hlDiI7/zVE/glJU4A+7xvuPtg6XWmjtmRbXyiUU6C
aU4jlfHVSkvbd8s0InKdhPN/ywCDmnA73PbR4cY3MBQ02hOttzT3NGvuXRsdyM2T9/5urbdrelxN
wMse/eo0Kcm8x5K1rWWhkroyUuKnWyDTqzY2YOBka64moZlHBSR6NfauF7bjrAzV0ZN8F2JGhhMQ
600SUmYF5eSKVuL86bftDYAlk2XN2/5hsWpljYDuSJK6fPEZNqCoPZD8w0FPbxrdmK0V7NA+h8Dx
8w2ri4ydy3xmxM4DvoUSbI24SSUDp716zAJ81D9KRJQoe4VuWIf9MYBUVVrMSB2oKrnYxMERh6/D
qAMC0AU0KPRlstXjPTi1ywE4zst71LypXsGoonmqiQDjkXdVu1K/daD/jF4tUy4avCOOqpuhdslD
sONRgBgp9rcRtKquGeZ6mZ2aeeHbxjVWZzAJKrCVNgfuYt7GD7pDIrfFof4hMPLXI9/PckBbTTqo
Kc5UtGGqCAtzv9HBMiWyUbFtWkLovMMGYigbkBvCfsLLNqWAvUHzglX4yzNGmggjgxA3FH9bwBTq
Cvyuv54q/uR7EBTESKu4aN8g2GUncmclyOITmBZBZ7kQz/lZiuw6vbPOM1ZVec66uj11JnDZqTou
0LLBkJsMJgVTxwEfnQq5lWsx7cV35IvtO0XOxHSOxDhE67Avi2W5e8KyPfAzG72LCRd9LRHXEelY
iZaccLVRHqGq6LAqBhyRXLgQx330EP4Knzbv3ff5l1sviXhOQQRfVB/DVObPKhW2NNICBX4sFaFy
QPx1LL09SNF09BKiy2VZrcCNM/xjTWq6n+lMLEkD7sMI5RxovNVDHJp6QEEhD52xZRJGuZcJbnBQ
AF4oiaVFSd4pFGkt7wrxjqI+Ip/IEPjJ0bzgwZK5eaA6BP/zTBysPatYzwYAlOG1MVesp1PpesXQ
QWdDfm5ZoVQ5E7IKhqkHQBlfW0RvmnvEu5aodCV6ZPjVyGtdNJr57C8+G9dg+JyzYQsB3QaepgnB
O6gi0S+r3IZ7Sd4J/m3RsHrdZrNnvLJpgcQGWJ3bpTLY0TJv3jnLMw4iUa820rzst7RS3z+Atujk
VBcwBtCcwsyNZDRlooTmKOto6whaV4yPJ7dkzSxHTVIxoupBMSPGB/p0mvzkbemFD0pUWs0nY98T
X40IQF9tPr4a5Vs2Xy+odqLxa8pQP0/ZzNdsD3kceMjF7U4MoPG15NjbYFpfUsIlv/XB902x+Mhc
mSiLcigQfT8HsabFSDN2acP9aPAV516gJ2XQBQA5PBMmNcJ2Eyt/x9SQNTsVMYSQhXhHtb9u6suk
ACwUZqt9qTG1uUfAgWVGaYAjtuBTgIBeDEKxbQ2WCBFxtXcpAJ6rt60Lwn8Cgpto7dEj6JiSMSD4
LcJItDahAXmiIivSjIKxKXqeno7YHDxcxxfetXfn1cgxvE9+yIV2w1WoBQoh2ZdZ4EnWsCpw2zaU
lsLpxkKqZbk/kpAL0qC+7Tq664kjh3Jfe4uSgQOb5pUke2c8e7GerusypJv1QczhgSI2QPAwF3QS
ky5jyvD4vt04Vd4avbmV4FsknJlJhPyaa8B5ZbKtcTf4T9wjct2A2lLrhYvmz5WeBMX04frLSh5l
yrduU4Zz41wp6Gd/7DPhHdbpxlxCBN6usGkPa+mReTqWIfhbbiCqfk28cmeJ5e0liAZjokXwfpjF
69Kdf4+ShpSF0MrimqsWxBTNur/jCBudd0Nv8WMY8HNIxfvwXCvROmVNFNa5oexIpzdcgrfeVq9n
CV6BdPB6RB75hdypC2qRxSElr8ZyW4Dp/lIzV8fWY/byBYITB1cgPF9adoxQnvFLKjnshEbGb7A3
LZVystbgjEQ15pta7t2Hrm4omoRgWcvCmoV+yMIzyNrKG3auEDzWTViQ5C6DyQmItG/FH/tcPkjY
i4DkXKUeazvB55URiBQuqwKp3AFjvvNbzyjVOTSMU3VUQqDlUNcqy6Q9ShHOSeXIBEIriORAMryg
iF0oXdlFHIH9EWkF5onN0HCjcbUdICwC1yUAeg8XI39vBPj9gJ6JoCkZOKAkmJ7fTedwFoPyQ4bP
Ewq1DvPUcm8CQ1xDdqnmmMucBykPm9AGV/sGJiSfeA+cOJE6U9lGEUyVOsmYNCmyym7N4X7oNGf6
z2YuhOU61Mz9AmzwxcqQ3SCHlEJAiJ9KGymRHZ2NmsOL8RbXtbru9Rv6M2xp6BUxUknYtGGmRUDq
6nxNTk7DPOilSoLgAYGyz61TC3gVv+VJo0bKPRkMEOAyvv1M2cyJvWYvulBfZ78OSPu4N5CB8iPz
HaKWj6RDkxiqXYEwlNEUv2BG28ZEIiLPiSs1HqBlU54/OCSUHQGXK4639JCtok76Ubafqe8hMo0u
hOXd/3u/100RV/YcHTLCcacmQjbuIo7cR2moZ/G3PqSE/FUL8jljbsshXhAviChUG1/H3fagqsH5
p6M/C0ag274+L46mu07gqKexQb4WqWocc2ORFMhGmPMrC5Fwm42uxxAksfsTMVjfwg1wtSYILYtI
QoQf7vTc9zQpfnojbLTWc7Ck6nlMSsVlRA2QL2Nu7pO8vYZsfzxPPi61+s7gOIdm5+A7j6+RQmE8
Ndz+O9hchEqT32AkNU5E5vmglBC5K0OtkXqvS2WA/+xrm8YTC5ND7VNlvCwMxW20qOyDXOR8Sbt/
tLmdMev35HuIPgMhQBR9NF1k+bYCTuP/u4rPET+gmR0VJs9tTRG9k/M8ImgJPobi5Jdinx8EAoTY
vPro/FlBeZZ72KSa0SUpwkYpwuFV/Zll5mbVuMfJDqYjPu/8Hqc92DffqK0woqYzyOhIoqnadpeg
LjdQzQaR+A+VGnS4bE/vz997nmMDbD3qyJqCdB+U0to/7K6v9ToLqNqVDDGruW+bKutflfs0MSX7
hLgIQ55KczQtyq2pCRij8nWYvVz+87ajqvbahSfOjJoANi0pTdAqB12TLubbFbybolMpNdzShj+j
BDkMHKurKjVF7hXCMHwjiBTxgik1T+y3eA0h8WqsDCwgwfmnFNa0WfcggpxzF6xJufs1HOUPiJHr
VYaOSAX5GzTxv96Lf30t4al4zPT8Y1dU9aCi8iwPR5dBSRqtYlKh/ZQLg9qb+nsbQTD+VM/iVnbO
YEEKWGiydO0uvAG06si8y9SxwbeHnTqM9FNLe8e3/poRvndzFoXhorkvJc+Ho8wduHVgJ5/1dlo1
qMxaSqOrXQ9TIlebHtSUS5YKCwQFGDeeqvefqdLhb3Fb4J1h5azxWo7qeGvCquJ4q7EDbH5Nc3GT
ZHif5Kcb1Y1L+qprwZFOtYu3tbqRN2U3LeLouFFVlgKrO3Duldj76A5hUbKXOWPH4M0QkpT08fkk
Mj/MKzqScRydkKDyjWSdDcMz+TtftIDw7Ur7PR8vRmCpa12wt6q/zQpCp1Z6YUirp2OnN6IU3yt1
wYhj3yC3TDCAC6nu1V4U5QnIlW1/11SqlXadoLbIpXZCNaMLlwDx9ReuGcUiU8fvVKYHfGV1Rh4e
/ddmtDqdslh20XAWxVfuQBR7/zVajAB/CK+KhfrKn54oV8pAdCvDgPiZv4yC1i0z18bD9Z4z+y1E
LMA42hyHBLn4JqVeI6kpKBM/TR6ztvAjzSLzUF/lGJsnLFhHQUToIDCWiLGQTxa1dv5XfXpaltT+
cmWWXV3Da+pbrgkyrWBBq2R7qDnLHE5CweAGAtu7VKmkV6/8MQn8dxPsMwRRZxVWwep5z8dccPp3
u1eaziin5n38ehjt6nmEKCxLgiJMQnxVgAfqCAshJNG4DElcCb6IDl0+QPCIIkxT1NfYNwshHLEF
O2od8Xs3psg3dG2lpNdXttutt4m+2SYYjKTyOezLONMWIs/bt04G5ZcHa3kightjMQIbNHIrf0sm
LozbFbahZZYcZrWl40Qag0liWSE4ZtqVAmxhT6Cwoh++scJxfmBnfqw+P/t9P9uke2D+kGhQgeCX
DTKA7sdzQ95v1n54tBEoWUG3ntsQ7jjKetYU6istYpCB3YCkGZnB5BN+JzsCKQg8qDfuqIdO44VP
/KggjLjSq3qr2gbN5sLgz866pdSZep1s853SfosdbHqfSUQKruXIr/asnJfZiGtJE4S5wygriRWK
j+yMMziDs552wHZQ/SqElVERshdOPl8fFtskwIEAniyHeCkTyJWnEMn6S9JE4x5wJeuwsMllv+8w
ECNcFWOP0lsX53Dm0xB8XEULCir/zwomfL566rRdfNbnFdNzWmU1Az92TbmEHpNEx9bcygsQhkNf
Xss0m4bShUeGJUdwGAsJ2ORNG52EDPrk698PRmBeQO4SQjDEYes4Q6CF+j+5AzM81ZVNjP168WKg
k8/NW8k/mbmfwOmw7BcoubkFBPRUiSBBuuvVeXrN1wCN/R6qL8pavFhs6wSiEhuapZz9i5fPjGD+
ya3NHRrTcwoI9buwB9L2AW19CcGlJZQZkyapgJPi3ed/79o226wC+8m96rzjHfeqZku4dB564KO3
T0+kbg4PSEu4qvueU+Hu1xTI6rp//MxjKoTXuvo/eTiVurVppwIvDUwTLL5fBRNnIZ7jWDxG29WH
ketEcHRp1szwvaCgcUjw+DopyNRNcHtB2xDSmD2NfpWgDDW0xRmNSCR8Xum1c3LI3J7A1KQXI1bR
UGHnaG3aWpM7KEeQRBwvCE0T9L7RghamXf/Ap4OJySOrGrjWbjpe2PC4Of5d989O4EZjc0wkjur3
dWzA5/A2kfSuw4+f0/f+svisEDtBfwNIYOgOaV09c1Qt7hjmRGrw8ZJedUZWhPqpIyfOhjUtWYKv
tgE8ZhL63hQXbESBeJ9rFkOFdHNab3SodMBqGqDmBGcI9nJD8ro4PaJxZybEo8E0XKsDaDb8axiV
Xe0GFSwGIN6J+GWWXnLYtu9chn1bi7vlK8vBTlOBfFpMPmC9VK5RXSNleBgatQlnsas3yHt78ABv
cILv+O60AHkl0/YvIQxEx1L5I/54pyXFsJJZCltQX/9len9hbDUxFUTlFs1hRZbA4kwYAb3yvNcS
AF3/WsIaKe685MMlS4fvVqYYmuj4dHd6sYa5k32xpRtPJU/qBg4Fmrzlhsw4nOqWe3Tq75oFKyH7
ndEzbaf16pmCs86M0DwtEiC63plrej92TOEsVQzGKIimvGwlOS18pA4jthK05MdvEcvMXm0fTo6W
gtR6yhF0GHqxK17tdGGXua1reGlagOoTdGTAaMLrHpMi4Q2Vo8jQDPTjVJi2wqg9wc2RRfMPqmPB
IwiY5YrjJHj8hpZX/TckP9Ls0TOtpTvL79QUXoyhWMw7S2MbUZGAdYDX07SmK9lDhgBr6zEqgp3J
VxCqvpqP3nZo891aU4Xx+s6HG8YgrmjyI7MIAGrAPmgvD15dUGwW48D0nqK/r9OKZ0SWndl6ZWNT
9OK9gznbjLrftm1NK5G01Oo9L3qzLlNYDbQAu5zuPN3mxiPVd1Gw4G9hsKvCRJl4NkyySU65dNYI
pHJNXnml3aHydBAFfDOyrbSqcbLXs+nJQzgWiyjCK2G7qWqIL47PAASpaWuf3C3wl/O16feFoWKD
NdQwnsSDSp6sr6aH6o7BB7tJTkodgIlAoZoC9XPqc+txH8y3mwmuyDsYFdSssxVM+1CXUy/NyBey
5bORt8Yjm1ba58xx8CuB3j4XB/lma+OGK4dMUnD5bpiZFbMAwy+8++J4xy0xaK4vbFUVP1cr69rW
J6qGG/obQ3UsaJVPgJfvaH9dCZjVC4F1K+GIe/0kIaZfu0KO++74CV1LH7CBQ9B7UYRwA5ugSb94
eXcA6oy5JPzAQFj1KABf6YHS2gXf7O0Sf7ZTqkXTVyixcZ9vTMNXp/M4g/30kW291j9NawoaOPBw
vQMR/YUipyE0UqQ5Z3K8dMWyfih6SkxJWu6nqQyJ7i7LPmLZfJtB6T2VoXOMotdCkcpqsxAtogmn
hh+X8hT2IxWMc33Ce1vD2pb1mjTSNZXkgtPTDbfIE+5OkYrGVXThbR3VKfSoGVttfFayGQz5l5XC
tXzjshHlMjELp+kc0CuTyDgrZg+BXbpqavgaa1URdIrM8gpKksTq244l7MjG2kZfVDC5pq+s7QOH
XxIgjL0AxorR+UNfEbanGrIk5w/zVisO2VriINB76QILK0sFz+onQVH1f7XZ8tEVpim0MhLEbF2s
+3aMyByNJQmKBS07YayofIurPgs3uZtGVXdLhSdbehh8EjoMWK8aMyDJbBBWyL58OhQ4Q7TSCjYY
kKSB+fUzNpSqutSUxwRo///I2cnOGNp6ox/77qFtfikwVsNIPvyLuYtsuNufTRKKb5A1FWafgUQj
IQqjGf5UCt1jJKllAXUvDiR0guOxRzSGMQGqhpR6106vUidBWxZ/D6VFywsigC4G1ubMrKCRSEMP
vgUVMosWGCy2Rd6BEdwqt7eFcU+IzBGK5f8uVrA98CdYwhjF3WQfAJklP+u3Yskn7lo6Mrq1a3dN
1bpRgFOrlbIxN+wUN3SscJxo6JofF8wLLc+ZiTdC/EoldOOSPQyDejRyYIXtObAkVfgtkWABcn7b
D+lBrRo7hZiIS4L6I+hJceiYWU7OC2v7FPqHdZtj9HVQb77NL4agvCev1BhT9458ClG96WyfMncW
pVMHzqMKeJSAKtkI9TjwxTeM5Og9672GAbQZvRK+8J+/j73bRtO/BSb80UY9sfFdcx/8W9ZUm5GO
vv929rgYXlfp7JK2STWm88CKPMRwSNAxu6Fu+82/5GqaPdPtVfN+n02f1zyMWQHgWul8gGMNw47k
Koz2Qlzw5MFWulNXUfrPaPCPwdU5u3UwzEx8lJp/t/bhXYrx5IUBtAXlrfo6E0zYhcotovHo0HDD
R/xuVCPIlVT6lgMOQsJU+QQa/iJrugSDpXvIOdZdjK/1Ppl77KSpBDtYb0fazhGI9/koxl8JHyl+
e9emEbhny0oKK4hXBPCey+0FAUNkqqniLN7Q+BWsyzIkMDzlXNUJtnMp8bTUQfJIq0ChtUvbZzVX
RbMTkrAL3WfNMrjkY+det+KpJw+X/KOLkuxhHPHgnt0MJkLRTlkQ7pOJOrErLbRcQCFwjjduhvuI
kRezFWAmG5Cc/uSHwPA2440D0qZxt4r4Q+qBK++rSOejiQaadttF0kTpUjQAAHY3kPa0FX+rGEoi
PVe/42D1LQzYp+rI0AF2I040sYhQ0E0r9W9nVMB/APzUYf4aZK80qI8vwa4z9WQjuPhLPAfoe8xn
Dv65pZl+Td38mVe/v0Wxcl1FUAhTexeztlKKGIFFlzMmaduXrRHb3owGSECy+7cnA9I2Upng8CFs
L9b4odWd7P+C4S/mDXdivZz8YYSiIs+8xsW1u7QN9S66ZgZEsRdKKMQ9tXO/68EdXSSGhdNAK0xD
5P9ZEjVpG2PdtpnR9hLho8eL2lTd93uVAqWVroTa0i5pRykc3DEAPWJ1+GLChTdGEYXRcKNe5NO3
Evf6t+0HmGDyrv4ph/kIBqsfKNWpsNJDpNdl5mFxwLCVE6xAN+N+7ISlXmNeBz7Co7KbvZRPzDsI
TODhtzGkq+9sJETADGZq9bDa+JQkxomRd04pQv35YzcFLwUwqxmskQ68UkvZ397LvS6eVxd8JMAt
tnx2ZZmH0/dWqbRsBdyNiyhGgVCMfXIfPyksCGLNipZ+YHjT0omTBlzQORUidxBF3iq8aVRe8vxF
LxGQ2CO/FwcpbL1ICKVKUrSCZdvXba26OpGhwih8SX+difbO+uePIAD23nZ+tnjVJK+AsaFeatRg
Ll3HVmv9JScczPa+ByLQD2uBy5uUxNEE0vnETqOriW4967CbJX8xD0wzpp46AJHSGpBPVARI7rZC
Zcs5BHOLMsNeSn83fqaQjlfyAY+aysVoq2vFb/Uhv+ZvfxX9H4q8X0wZbDhIoa5AS66uS7SMa3Um
bVCL/fWpUAD+7OWxPD1N/4yQ9yaTU+Jpv/F9grWjk/hfJJUdmJZsohvTvWg4ne1xKMTn7LfIsM/I
3TjoaaYCaXjjH7IK6ODOm9rtA66d9EpHcW6aoet3CPN48LgO6nuCHZN8s2Ca3uIfL/ZUr8OXexWF
t0kVxoTkqf2QkHtGpg1zQgDYBnfYCwc5RxnOHPl5TGBmuztVECAITQ/ix/Wv/LLwUymF0hxeqR9E
8yEk288uzgp537mhDxYFyhXlanKXBon94HM32dYxkmar/qT1YxddKlKrMVPpv/+OntduUBKQB0gD
5v30LkVE313RusBXPkzveXOuNBNO8HxKGwb12iUoarDJqLScpS6qDB4DyQodwL25NPT3h4X+ufHr
DCR55hLX7khNBx08yCFN+wWyD6UFT1AVRJh4twx301LnJVAbleUdCJcXF7/DXteOUv+/lPDunURU
UBo/UGSC+1Ytlb97dROPyVSfNC2e70WnBO21ID6oUTJIGZDXeJtmGUKobUClb8WRH5igJQ5ErcrP
SxRt2zGVc1bMFbwuI6/g2g9Uc6JnZ58tYX6jYywmfzWx7BYH5cT1wbamCruqsIirFV6b68YsEsyb
WESi8W/1h8SqI85R2TlLlyYJzufE7BmddIEO78kqMFTtIPbtXeo6wuaY0eszPl9/8FT/bAy5wKBf
e06fSjo55ZxurdOt9PAf1eXg8RK/TccqCe1qycxjaMIRyOo9KiWAKPur9Wlldz4UQTIU7VoL0BdF
1s7cyJB+CsxUe2a9TJL9oJjhV4BZtUc+ITSjFkJAQsn/qFFViCZIEa+Wb4EfNrIsjaRHvrt57qW3
jYZEj+hciIK68+BK2z4KME7kHWo3y1Ua+wqycGLdaJGgqeCoFYqjx4laf1mMUPAXwC35yU4JmAq7
ObHoM/Z8p+FE42wjwC3IvSziprqM8KEjSsE2RYs0HbbUJSWVBS1u4Oy/51u0ex9yssKDy+D5w52M
SD0Cac8zB+8+bJrcoBhpcwaZHODW5xZKegnETC+bilFxx6yU6YVlMpeEMt52t285x562TzyexYdJ
BVzbmgUX3SJVbxj/5YlhSIB/ad/PVHaD8U+0X4jWPzPZAqrVkZZ5HMeW5kBTptZn3Ssz6H8PKXc6
p06nDHw5gU3TCuXmpLCloK+Ukx/IcMc8xG2cFet3IOzPbA+nLdDKexz4iy65O07+ke/mW8Gg+i06
b9ta0+l2KAU97/BaFVxe9aUKhh4Utqr1QoNxsbtGw8ayXuaLooZ55jr7Fdg8LyyScbt1a4hORZkD
8BNGZUZXNRFuibTL1Dn3u5vbiqtGrpzXW9nOGHuL+ukP1SCvyixQgQx4/YyL6RIbmts4f4Y3OFEh
jSRlGSPh4nO/tdmQBb5UCcrZCaaTvVoxtimrHku/DIfn3MNLT/165MkYhVDxz6nQou6RVQszV8Jc
ltBSg85Qt3jW//U2F9/B3Q2V0kRL/fDQ1FyyewtAH68u1+1JroKQH3OcpevKKOvvNx8XwX6iPKsv
xzgEWc0Wf0aGXevySctNvLx2zEzBLEKNBpyuTzSG/9OTJLlmyJ9SCPlHWjsX6S6SaTw/oU7DDVDp
Ooru+ehPwvTG1EIpDqbNNber3yM9C+wCMRv0uEfYU9Q+8no4yztYfTu40EZbZPV7G8rIEvT1jvHO
qPs7GWlmA3NS10U7LEgZkbChgfJqIB3CSGorhBlaGv57TMEF0oGx387u/rGy0iVtESNdBAQySHPx
PuNFUxcpbaxzhdkCPC0ef+dOlhXeWgY0fEZ37X49Lco+bZahsIavpzm1g91tDvRA7IMtobgpyqxd
wKwh8Txnoo5jmlFMimbZoZkpr3QyyqTfTqvLAHmL7lDg7b5zB959Qy2y6ecM3+lxwo7enwOHW9mq
p1IsZ/H46hAj9W0GhGnNriLEK0qpfoinLZgGqIKMueL/1yNtWL0AzrkPWlB9IqaTlqqVV/PdWc6e
5PG3dQgfe32LdyOEOeotVNXUk8jURFt2ahXQ4Q2MfmD7VmYkgtvPlUPFDxu/moh7a7xpSKPAhjV4
XeybKJIcR/fhaeVPiaZeTTiAHnfjB1woSfNOKgtFSdd3lXfRtaf5+vOPXwIZO5EkUHgzhiyTIkqR
26t/QFyNayNKmNnCed7R2uoKeeES2TN8Yc8dK2qurMVwGrFvviMDyX+qqEJom3ASmxiMOIzYprz8
mC9KPhBZWKRTmYTBe8nUo+Os6p8f/TvFqkY0h1Vi9LK3qCRurKeNOpjQxdp05Pt/R+CbYoVdtX4e
zw68OlsIfugcRm/rG9Vr1mkhHRlXNIHBjGriRhrQ9+vEFjTffOuSsNo6nXkMwzFfVbAKHJ02wEJ6
yhE+1a301ZUrhYjHX8hWbU9+R4a56TUO2QUliH5TJWCJ6xGBsgtid+Bm/ic/DLQn4ds3c18Qb8zE
EB5XnJJ8AKds5rgEQURlutGx4kPdtntW6PZkiU4ZCGv1eSxv6bG/QKAOU8oqoD0d/PDyKmJKQhVF
zHgWsKwSYCcsjweEmdesScH9j46SGZq3MhRkRPugC4e0R7SuaAusL3qvrhgZgKh65uwbe1tJKYq+
UvvgxfJ/mHgN/v3v7rpcBfv+b+SkNoSr6n+XRrdj4Uf3DL/PhbUSLJdPM3JkeAijI5oiKCQQGReN
LvIXMBBWOU+wIij9MZF1DO5N58Ywap+KcRjWAlssX2nC6kuh1ApFw421zH9RDDaQ0krKFToGIoLG
DmJbq0xuH0BqRjxJx43PuJF39QZO9ldW2o7pfCcBiW73mAe28arxI4SJzuc2AIGJNmUYFU3imXiU
ZGYB2tu0V48x+grfnGFpsZQllYYddENLB+UVgZG5JBugjcZorm8Id0oBEsflgkSNdKMrQJn5Yh3D
mIMSR5SYyOX5G8hX/2FxZxYstMJEG+kLAr3NbWXfIixg3owfgwufFm3EoykCFs8bDeZb/SMw59CU
VkfZsVwdvolQr50b9hy1AKYp80UeRtRhjri49jxdwjP6+SCuHwG581sFQsgXNch/p7EJ+0RF0OVz
rvI6FCltnkzUb4Qj+ur/pl5ma5Q1d8zMtmiYuo+YLD2Sm9oULcKqLkt/e3+OctE7SElklT7zdud3
K/iAzXaEmfFwudDfFf9rXYyf7WHkt6T5VmTqg5g3RuqFHwb+rm+3BGONU+PKQNUGQ3GA4SJyhhbD
a9N8IcNw8jRqNvPxvGvF3SNtyGvINTyL9aN6ImeOXno3XnRnMVc5qDt+8SU66WKsZJ4SHRvHxIAg
7ZGuEAhNh3s8ZUUNnUY0ywteo6DPJT/5QaGppU3U8gg8QHD/9EXdbahOkIuFy0Prs4+eafy8ie3F
ZIqdBx9fwOUEYBHO/SUeSmI/JL3ym8D+SrnGxmwUisPMm0WhPMwhOm6r1gz0O4vdTfWXGKyG3+pU
IU6y2HlQJSZf9nS9p8RdjkTCZwbrS9fc1YWCHYm9vuOhQOJ8ffkDIEbITlS1MOJf7D/qjsCGmOTR
N2bquyFjsZQVlu9frMdVgDeszSQscurkkPsY0nFuOV4TclGR2wa1defDINxSSFRWm2Dl22pfsrby
Y4P4A5KI+LXhGt/UNV4q/oWkuBl9CE9MkCd1HtbTNk+9DGUnhucqeuAT02/7I8wvbniSd5VJJwBz
sDbEcQZA7AoQebvqefGMFM4rY3KGNku09ge6j/dWMB++vjDdsyRJ/eJpsT0nU+vd1LAZ0rje/Rvo
OwxgDndSrvH2yJfo26UeXEADoaUwu7DtZd/YporDqHEKfF90M08BK7+lTCg45nhw7ZS29unSxQgL
PnM6btAYFdQOTjCyPaF9VdcRUUlI3XsEcXA0moHME94Zuyixlh38zzAt8ep9KLwApFBgDAgWCWvl
DQ24rs4ICcW0ukxpyRgkzba7DFx2a+jPIQLuFx3ccXoqeeyg2ckvF8yEdDL8fBfR/dJ6PoHIHXyR
aI/gmmBCZT48Kr69/xOA5WSQDJlAnjy2iOj0lYbvRtnJdcwpfrOc9t/Al4BDKHeahlxDfpLwJXuO
uBZFUW4bec9ahk7oj5Uct0ciI9cDqpOoUcMBwNBCnwGmY6JkXjLJCj9YJAu7HMw/HmW0B8Mn0nMT
nyRs9EHYKkQkIIXIpmzNjkFhMxAe67++1Ms9IDBNvKC70Ojc0KmVfPNEiEp2E/MKsWJ45a34ncfi
5QbTUrcQE4J+QoaTx9ZciR+e2z1bf4+I+TKMedQ2q2ZTVvYLkmLfxocsAfY4jSSt4/e8f01I5m6/
aRF04S0IeS+/kuxYV4lqeS5CBegdnV/qXswe6bPVl6XOn6x6lqJRNj4bAB/xTuKkWb9Nf99lEMUb
i6ldv0iLadKIJzfWJEI8+sHEl5c92RlVh6KlagyTTWErLvLM18w+yJYeerw5nf71dwVmiwyy9tmH
QxLZ0Tkyva6G/Js2Wn0Ar4OCCINYrJ8WTgEv4gVb1oDHi4FYq4HfSxw9UODJ87z3Z0cILk6qegep
88hqpzx8Qlckxb6UyjVGnWKrM0Tv8e281P/U3Ye+bb4I5frL5qVkffhMC3pvondo6AMIVwEIZ+Wc
JOgm0+uqrnCMjwOe5jIV5F5EQokpweQ9rUopj1SJc13+Mwnuuth6ZnUXQHF6AtWZ7a1UDGkZSfps
a8fdZpFRp6zBpJWeMKJAqwVgpoMwEjEZ51zoRWSI8p7zFd65Vez7kw07CTMXUimXsCxSCK1C1Re8
1GaDEfkh9T5Ko3ohWlOwPX5UwU9MKEWOYvvP4CblimNHFEWZe22k9qBZ9xEkomlLaHYNzJetYiFA
HKTbxoMqtC5B7UOkDQkWbuRbspCBnu/P/C2O+7mShf/2lDhGYgexTUk9i4UstPkad3RRfb/bbLIs
M7Ee/g5b5p7+zPvLRQcnGN12PMimjA5r0H+AzmRTKtP/7rIqfcb0sKAKBKjVuyZ/XBR91J4TBt8c
HdExow8edHEJVBoEvfr/f6PSDcotzeNpRBudZ+idRg4BZzNqrtqYU3k/VX+oTvyhJX5pfw+G02S8
8xn03QS7z0A3K4P2tzVboWemYRRaP0uWxTFWntDZWUK4fxSVzbEDueORGY40MNUFe63Xt6/0PJd3
rl59Uy4N7m7oV4l2gkU6AfgMhm+DcRBy46hOjE9FXx2xZHRhps0qJbktKLMf8JhtsFqqKhVlRDYN
uhFU4VnC0YJnlASx6e14YDvxsB0w0jAK95Id8QQLIaHzOZ2p84kAFlL8Wi15WS9zGQQUKa8vwy2m
8t580IavSENMDGd1zMb8V6ExWdDiJaMuIeBoDBatUMEFTdFPSjsQ1tmlEKqqOEyE8JE20XLzMYgY
IsJhKVGZrb1EcO7YF8rQeo2A8CgPsfCDJBgLUl5auSUxmec3Jr+BcW4DjtuyT+qIini1IZBrkkcp
Y75R2C63ftLGxtIK38Jv6o+CWVPi+2D/eWdHdJxWrMa6Z/ok0erL9Pj3JRYdn1LNkHj+kOKJLRdj
S93+rJOYNK1/cIHuZjZ9tqz9195TpVIar49bIb28t9YOLc0boJpGTA3AqyyfPOtxOdm0jgnLNo1g
jh5sY8PKpWFjUBOPq6VJ8V5/zxNUfT0VI1QDmdchrpshnK5POVdniEKheCGYGuE92T81hCBfQy5W
CzjiQJiwyboQm9nzCTofvxKmlbVMoYlXTRylhCdYRem2vJOiQWhn5jqIWbYKC2q5oAUoh0VNPAqq
axuxSPlg5dbWAqsw9OrWibf6FlRTzb/XyZ5Qd+IkSE4Z82pWk4Ip8LDXRwhyG1vadPM7gP7mvHu9
iqA6hY+mXmg2MYxWUMo+xXMmqpfTui5GWjYkUwq4eljBLHagXh93Fxbsub5+szDgfHwHThN84tmn
1tdk+ZNfvd87FyRqW3Yupqo3H9zu3/71C+kykHTmBpCASvOhs2ZeGQ8noodobjBDsyWqfNQtOh9c
uOGXznnBRagN7FN37e2s0s/q0EGLHF9hRFjo6mc6enyMi+L5BcZRSi8jNXhJ9zxr7UraR9l6hkjo
mfQv3vS+kMSsMTC5WOLhjYhBoRN5h91UBOLZj71A0tYoTNfbWKeAD/W8Qu7HhsWFlXzHxr6GB7G/
QKbWvkMtjv9auW1iP0CZZyXnZtlvL923hFYBxplI51wfgiU2ncRDZb/OPNg5OHhFv7brpV7fsi1I
RMhvMeyhHU+ND7diGEBs0qhy4lMzUwRk+SiEYXC56wzs2ZqMP3/BmRrfdGJ3rall8xRuDIQBJw1w
9RX1XMsPWTmDny0RtWYkDXloW2kLTp8ualiqDkWiHyToKNDG7zXY20ygfD9gKjAHyHHUTbI7pqMc
12WNuHnV3SHpYjBg3gmVdHDtLI7G12fwSyblaDciWmfs+anZiySow6w7dYYqNg3IA8qM6ALsNBzi
1FyhTY7OXj0I3mPsWkxDZxAUt4iechBvABvC3gMY4DCPE3BnOX6T5hzduSIbuRed9X7mzm4F1Gbc
7sdvPw8g7Umbsxo43iDelV6eUf802mQC91Hfq+1URUPvN24T1XtYOf2icDVdNPjeaJBdr0ikyG8n
+WgJyyQJfglXL7t4OFStQDnQcWV9v7ln7CSv+YCHxuB/wjOTAN/gdgllK9bcUZjpRTT514QU6+lJ
eHvKdPdvYPSD4Tu/0jSlVrVJHp/UWBR+xobpwAjXgvH7DM/m8PLep5qUGi0qT5YuGsrxPqBMNJ7K
8429Z1Dy6tHMox7+05ycwsWZCIoCn2+DYc4BjGTvgzHUzdBaWWzVxN0aEd5z60KU2qRVWzjjcYiK
PdtVwp2VPz2KhRiJg5coUMikX/o6/EW8XcharXdJ14i13SOgO52hJcvVBxYj8AwWeOJDeOhFs6Oi
GYbo5QiCyTKhpRhudZ3S9aYnPrUiA1D7FNxC2WbqtLA1pkCbwdV6cf9/HDnwwBKryyVvHGTdt9Pq
/b1L4I2952wdF5KCWdixj00nSZ0tYrIJI0eVN4FdM49B1oUK5YgqNl0nmvNAoYAAMPAeGRuhMtQ1
at9sb7sRRoZRdZWh5Q+Uqsjx8bj1WdwkJXmKL8sT6i4L7x7Bgws4gZFeFbrCN9Ast9IG6ShR2RQ5
NGjlM7DLc9VcrDAZXc8kPuaTyS1wz2oXb73xKwOspESllIp4grTqYq2i7CRHPlMlHxDnlALN6Z8w
I2AJe/GUI2WYgxRH/bOrrKPyeZnOGlJNDVZjV6M9MsRahzmwwsr5uX4l1k8VH30iWpP7uOYKCY9n
fGaH86jcNiOsLmDlvKeAr+ObX/gOTq+ZjVLsOnI3I1vxqDj0nQkSFjhiQVXaUY19+dHx5vFC3Xh4
JW0lbJ9r62znKW+LdIdM5T7hxuATxJ7jjjSucAn+OfwWJci7aX5oFgnJk2mqwfjzzDis+4BzDwfg
AU0Ti0Cf2Wgexd3OPUYi7LYR4lu6Pwdq9jjrSd40Ph9M2k9RmQOwOmY5NJrm/CrhMMwwbEPaT7f+
hfpotRuvqUahIYkKlA4mLr0fUWTQkLTObBFfV7MVgpMOvBkSXGcDmsYH4Qg5zSzn/GLKBiS48mbF
4MVM3cdwPQNEozcjnR9+tAT5XNXu9+OXLt8HIMK/zXjBV978m7bjKqkpDwyQXXPX4Brq9JutDVWA
/I12j30XuQE8UhjxywM2oPvHgMD/c/d7mxDZ6JyWV9A77eh5iRkt0MmO5A/3lQ/90ro2p7nZgUrX
bC2dTSMK7TaYmlDBckRvIjo1Hzd/lTBlSUPexX6pJs1dfLqkr1ReaLzrKtO/lPV2H/YEIuap+AaV
9X++r9oUulGW08vY+HGxRsNhTkhQuBTeuCn7xJ/F57J9T6BYgzI6Mn0A1J8R3vpmdcfebw3eMAay
Zek7651J8KGSpxBDfVFkh/Z/z9yYoJ2b1tdKok3f7uNdVvHse4GsEuiK+YKeAKbkYz/rwce5o9j4
wCnYFRVAdK2Q4y7nPR6FhFbNQ1ImYUL2g22oyDuDBs4xq0tALilTCDQgP/khk9/vGZSJvzS6z+wE
gWC6mh1sMXgjIBoy000grLxjm6KEk5T/N+19JLe7cSRZ0V4vTAUwixIlxFiXCNqEmH4ICXbZPRnn
NtMrbskC5C11of8s5Q1FXhmebEqtXpde1RLIjN6aKN1e9IDCqInZW8gg9C86nSl/2kunVh6BZ8wB
mZrbq9ikwCn/IbNpnpS1CmaXVKh/0nIfatLD3BtWxSATO7CcLWjFeiR1QDlMNWhtugqhdrjH1r4W
Jt5pboi7bju2Sbe3PqWWIv2UoZyUezbileF1UvK75u53BZoidmGnMlLtTYn1rFkZuxcve9mDiMKX
p1XiDTq016U5ezBEQPBDHgt7+A8kOAh1xPE6SXmrvj9PTNIA8K5cQvDPZCI23LbGBHx1dyxPTOGB
UphYG4Gh7ZiMtdLghwR52zuulH8g08qiDZh2oRgLUNnuw2WyaspKLcilxd7PKHNr/7a8ZUaoLVsB
TWIWIR1RkT68l585IFhLo7+X20vqFgoI9GXwJqD2oe3W3hp6IjcKjwQBNczL4nKPmpr7kZ08D80a
dX6kU5zaiM0a+CebTu7M8P4OPxPn+KaZg/Noe/aqmdMygb5UwuaHHDGmng+65zrUtq+TpXzjj5a8
A6ujkQXVV3NSu+RGDN/V3xd91Sl8iYv28rTkmI/3xQCcQoJvQIarvRMfKZvi6M+Pb8m2/LWej9O+
9fSbMaO1m916hcPiLN9mlPT1NP/zcIKkkHgd6KFVzteQc2Tm1fa1eT5Ftsqa6eCmJYBkB090JsXf
+9zbfl7t8Q2BOeWkjuVilqCfB4gLC3mq/NmTapMjima8Q8mAzJDglNVFlpPoSPsXVV4IF5UbK2Ap
EeH/R4WfytRJJa2DYZT+uMM+XLvgzTvQSNkd2Ij3Ror2tpoTFC0kb+ppu0opDr5AmVWvqen7O04H
OOV10Do/5cw0WZgSpiZZuOz562j9X02Vikl4gTP6CsleaIWZKHXx7Gh7MJsxSALdGSdgMzYhiGlg
gyJjTdkImecwwNNz5OxHRR4p5FcfTVsD3LWYkWoB8Tt0uM6greAFoAklLxKxruF9cE3itusVEJ/o
0TvfeuANunHWm/QRXhwTV7nHL5j5p/rRkgNBBWUg+T6YG5zeH4LXNVSUBKSx/aga/0f45NI9Wemf
JGehYZQ0IxnZD6YwIH8S2WMVIZuYSOqaFDeraPjhkNfA4lPi27jRKtB/4rNlRSF2DAdGvJngo6vd
DCZGOIlIxbo8Cz9V8PJaobhbGyVOJ7i9XPUfnIABjzJaILClD0NII/KdRE6OOMz1t7jUalagGzww
I2PKjWyNUF4SpNedL2OoTWF0xyiRdNYlB0w42telR89+XrdVGwXSpliRmnZnMw71RAsg1XGAOu1u
3trmh8Yvqji12xG5E9uK+ZdTFM5S2zvxJn6FRNySigKzlqqzSRoEQy6pQahOglrYAlHsbCc5Z8Kc
dVtIEoy2gSZCeCvVHivqgPDHEFUkNc88QiLqDT8OaToFZYKl5xM44Gxzu5fhCaP48KigXfcdvUHi
7pXmLnsEaSQOKKg9ThJoyepSUvbNCyD5vFgHNfFrjQpgU/b3Q8aPknSQ1Qd+MsK/9Wq/IA0QQwYn
9rCfgfa0GkIWoYHBXfoSMagRxzAJoEwPwBsv4n2+/dQ0vqw4/WzbEmP54BQl6+sbHol0OPto69rt
j2vV8lSvi/Rsb2hqDffjLnIdN1HmrpRnyT63LfEg7PpfTE6ePkofcOo5VGb9AlNYvUtAk8dQMOsh
ukp+ffao5IE76teLfgJFXEaia6A+gE9oKjvgKGoTUfS25NAq9COBKBMq36RclHDWlkVMn8oCdg1Z
cJNLVr3YxFA2g2Uu2qgMS9KWiJY17d4VUxhmvMEhOfAdd3AgZC98RgGxKTVA6Ex23Xdg10j4pER+
iBAh+QCwSLYmQVL0BO7Plj6aRwWmHbLMVEeN13W1jqKlV5F7eIO9YOIf2ozIch+qquSTp3aXVUr8
6x095aSNNsZyFnqbKhbE+xDDZgfcz5tlHOY1CGDTmSxXly8OP8+B12smGqu+0YZs7FOyAB9iEjF2
iZbQV/IWVOjOuEg3Kzrwm6lZgmWvq0M/ZMCjDebMF/ObdLROFi52biTiSWlnuCTjM6S4RlTpgsec
VU1yjQUvG68tNeptcUg2U8SvyKFCvPM684bNSaqQq3ljedLD3/QYz1wtJ/dJYhzX8GhOYw38pgbK
4vHyiM3BawCtCbAQntxDLdJReMdsX6WSr9I+qzmOd7ks3FZHSKh5eUzef0o4R9fr+TpDwiLLE/5e
7MvnN0QEXMUoKNkVghg0WSRWgx/uyxpbP3oS4cBRp25A2aprmJtD2VpJr+gmTsyuG1d3oh8RhYad
ysSynwctdwW+AxshkDsAJ7b5jk8xWLXeSp/QT7vCZ7Vuxv9PpmQsomWMESgBli0g7+SYlWHrnojH
KeI8lMQhGn+yfNE84p1ssUqHbe6YBY9ZndqJeAu8+P0W1w8GoA2eME4Vb2oG/zKag26FGLki8cFu
imjBFvPkMHPxHT/0zxYkjoPYfCsw2jGEOLzKq9oUT8y+WsjZudzwC4fY2c6xWkJffEaMVXgwCTqr
lSEOSSEGY5K2Qw2oy8hQd+vggx1LzxbhnGW6Bwy24Js6TpyC/I0N8624hKmx5GIKLU0yyEvz49g1
T69MzZb6V5NnYjeW/rQN1k3n8kxJg/0/8lptRdVV7j94PtF8qYvTsk1DdFXAzQioMZI1T/hRAn8u
990h1N5G+uNM/WorVunsAacGLoFZmhuFIF+LZW3qfscAf+sLKr3tulwt31DSbxAtGlWRy9tCOIJX
PpHLytF3uc8a0yPH2dXOjM/U4udilZvioC1tRhdYwkfEQI/7eNs8hB5ZE/D2kuCXGHWEVRy2Gr1p
/44vBdQpGeqEw1Buv4vQBhri3xUkS++Xrdv0qI8QghkyI30bJBhY8rU2baF6/sK6DqYUbQ2sG6qP
gn1u8/ayhuXKMUqDPUQgW4W6/yv3sLHZMfTWJmwsfQ2niCW49C39ICNYasETA73uuh7tx06Gtfgl
ZXVprGMRVzFWztgdTNzMzBxGl01MQfSae0alaPsV61ndPVf+UnIR634pfyDduu6G/wzGMhiZO1zu
ZHLi1g2rzZQ5S3yfyZrpFriuh2tJhtcMVtChgEL1pvT29scg5JbdYYYUxvquwh3WWWOsLcdjcnJ3
VkFJz6IQainf5+hghW+hQH3r+VhzZFoy8RQ9AGjOEb+Z5RLcKGWnezb7/SvZD7v1mwBc0BNNUQmZ
mRSpzkSi/zoPEM7YOCRgI/JWaCeDKNYC5Qy2gFi0DwwX2RmR+nVVqRXDpTXHbWhFmCmb6Njw9uIh
HevWqT/4zfEpL5V5h0jh4awAdBhkGQzviPwSSaEOQPbWPS43u8QD0WDY3lsvI5PR9UVOPCniAcd1
rh6rf9dpAinB7U3dn++ny9HXd+nVmuQzpshvnsGVo43av5woPqZ3DPEJT6ltmk0mhKr4BWQb+KfG
itOVQflkBGInKfehnjWnnu22Joajm5koXR8Dm1sNrgTOwe6fXw/LS1aFIvWPdJ3y0CbrCCjuBieO
OM8uN1Qn0uaTlw60j5hovBcou1LxmDEncv75Zbb6MhY8xPpYHrk38oB1lY1AWuInJcKax0t/TEWI
csqyAxYWALNrME1+TRQ7JpyuXwq1NoFORnYPQ77JCip0bVuJa5KkbAZy/fgMjAhlvHx5RVC/vB3z
wjBgzaZXCLIZ7MVWwX81ii3Aa+ywJ0BBIXp3ex6Q7GfyGGbaRn46+iHIJmx98YWyYw/D66o8vtFH
A4xZHEBbrOlEETrFmDTYxSTxWAksBMYhI+kHRV7KsCFMaBr7ad7HrAXUGmB/ONBxV6jNiA0SYZ9E
FezaALJV5uHQxMbqtMIAKHXrJhRg8CL4qQI22gXrppGYDmSTHf0YGmZqPfu/s0NhG82EHR1iEQGA
nWHb4j3AJDh9U3esonxw+TfzYrDXnSDaUzKqbl5XjXBwKtRQOYmIBnI9Lf5k7rk2LlAvgFXcsbsb
xLoh9fCmR9aF+tSU/DlYkbG5kddEAntyS+Cc9V+4VMLPIbSj4LmCC7rGY3hoerg5y35IB84c9O1M
JV2xRodh1Cx+ttsZmItxFr4FoVL+he5JrvdgwItCpkZFckKADnEItAV+GbJGK9C2wysS6OJc31tk
OEru721MiQ4mZPUWppldlasf7UKfKdEZk8MJ711tTF+ZLgBgrvQ6/shUT22U+riKASnFfEiWaANd
XMcSSYLkF+NPWiuUvGxk8gXo0B2fS7VpEclVSLolVer0b6LowlojmOx45/xx5Wu42sZUEqgeXtZu
MFtjIsmIjPhoKu3opieWpXvD8rZwLzswI4wU4TAznE8OMIXNJZDljHh+ZDVVIYhDXCfpw8pFr3mM
mnlIEaa0dsIggACMZHqVzYh8MBngu/JTc8UYZOntpJKed6bkyDZMPq69H1616HVzrWpZ5weYFZ7R
kW7J4viqiUeSnm+QvzQE2XP6rsLWczmejEsLW1osvrYu7XBnbU1EvuxPz1NjWq3lI7eptTUtCyTN
bcAJOBGz57h6qovLQOEwc6E/7NN+RngEr2XjlZ4nPaGBfvy3d69pWc/eQqu6byRlti6owohUJ08J
7UmcxecASo/tz87hBIxMiAED84CI1gY4VOwZNyhMfv2FkLmV9tmm8ZCwqTneVoReLXzB7JQ2CPqr
b1KLAt7ATCkAnsiIlQdc1w5mh3yGLT23suKFaVlcSyVtbVZ6oY6F9fGTBYEmdGoMwMckKqwXBVGN
vDkCAUlY1QQeUodOEK8/lAb654P1PoA0YU3NUxnt++jIQlMnAIiJCRN+1itHRWF0g76FVq6tBM6I
w1kEGG54BJqrl05av7DGpbr8qA2hzKUNlinJUOUAuIxUEAAyyB+G1hxZEbPeNEo5AOOZZvP+8l5B
vyGSpfBzFWA3QoF3zd6UChzAAk4esUMwCySpzPlOzJU8zJSDVzJi1IgK58tMrQEuakjmb8goMp4C
CCtuJL7brMMzU4Z6pYwfyim1qvpEWWxe49YUhrd6JAn4aUrYWjRnUBTk34Hl2dlrDNK1hJDgEvIU
d4dCYn0X2CRVwUIRH2UdbuwJ7af1gYQ4Vtu+lWcLSWjeUKfmibxZ+sqp5WJd8I+wcSGcQnGVKAO0
IL/XOP3FKR7nxvf9juyNhn/OtY0Z3rkQg/OnkhvjdzV80LEZxT68UOJSEJAV3rW94mADnT2hIVxk
M77Q3IyKpjHTHILlg0o611cSmdt2nsv5BPDHW8i8wRF8niWeqCIbiubusIPagocOow6q7BFfJeoE
PGD7h+hzePEmzANLaq5CQa07UaRDtKQpzClwcGjzOWoyqS+8Z7B/Z1Ql70/TysmSXf/aofr/PyMV
p/t6HSznww+yXFzECEQIu4cqs1RZVr9DV7cUeqhsruhp7L030I3QhrbSchVvIau9sA6Pku3STexa
8mDzyY0GyapBGuPTeiUhj92kG0DBiBvRQOdxWyKBXfDGRpjoW46v6iW4oNMJHxSy4xPjbNv3hkY6
g1Mmh5UzxggA07FMZ6R1yCS8ms041KnKdQHlcZeRm8rs3BAPr1QrDIgiSLmJ2LRWkBxDG/jIWM9v
MHfVQrm/KJ33qDxeO0IF9Xfmf4BmnIlTXTdHwYg/rJ0S/JaEKgYcn1pcIcrUaL3WfuFi3P715Cj9
W+GVx6NYun5mO8pOED6+t+Tob2KrRMuOYRDLHwKJUSE3MpxsZMPv9MtHlY6i7Ucoa+6gNr7Fw6OE
CwTz0pweV+ajwxevKk3WgvwVhD/FZADnGqV7qMMA6zbcm+Ul8KQ2/jGHuqNPwUGDookqds4CzGDQ
ish0emLIg1Nzu84KRJCzXjgMlhJA1Ln89kvzdrKkHlVcD/oSbdeQz9VqK8BTWtKoM5Cdxeqkl2hP
pKNrq6U5CiUAXlps55NxXqOO8KY8MVvd01wt5fZZauFxoYr6B416K8Hi389XhB0j0EcupSSmpIUC
tLFyotktxCwvgPiK9rJ2RzLJZI2T7upbTS2ooao4ezPBOZ+ZbXifuxbjZdsGir5MDkAzGrwQ4YML
ZKu2EjKOVNp582A7T+w9rmx6gueLnGlDBoD4nVp+wXNDyg3iU20ok5/wz6wpJjXprrYU8mlOvnPp
2M57+b8DIg+b/RcoiCmZ+kZk2nW49XsIl4CmqkCogjmiWCWNHKkmXaLvxbvIImBQbO/kgVF3QaVW
2XepGCB2LicR1KFz9PG5Y/bCpkU60QLfz0e+2dkSaPNJ2VLbt6YKlAscDh7eStnnDxR+AcX/oUf7
/2baktiY5LL8cwMU1SVC0AAt1AjyLN7JewrljpOF7BJPs307QYQzICZvgRwXaQgzNjZJc9z2c9yS
mpwIE+HztPO3vYIpioDFgJh/uPJl9p1gHqR9lPO0yzQ3Bc/lx14AGi3eXzBklwXucOmjDZCHgOCT
91Uw2FGn9oGYB03BGa3XvOw3eBRcBvRsZtAhxhm2rARcxkqfSMDA9cRv7w88VA6fdoYMw7vaMcDa
2OCfAQXE3WU7+u9167EXQ1xccrKpccpSQltP31zhLkvpH9/qovfmlimZHp3EVv1FbNU6CLkQd11a
TEf79orJLbuuwPHucB9Lkh67JqWFLmahlxLAIWUgcr4awBY8oet5ZIUSDirVLVzPN+/PlHZhP+Gi
aZopGwZQfFVxIclP9B+T8C/oGxvs2hfZLBTzaq7NUHs1vcqpv76Tk/q1hYnhWlf1VcSAToNDcpAA
65Ph4rjiOJrdTbFBBgQ1HRFqHsmzoUxuqw2CwvhhqKfhqrrVdYSwKg3RlkbCvFaPyQ4GAHcwnkbc
wqTKUXhA1b7BQs8Hv5huf2C/HObLGAptAijLlYb7iPy9gZOsVRneuWm50XBtiQomZYcu8AGQQR9r
Vfpf36Ej84MXlrp/N3YTUxcJRbxD1EG8WBFhdZdVKdneOEwTZfS63fbVR5Fs9zT+sQZHbylM9qJV
ywOq6bLmGGdU9yAw9iYwCJL3BoG+ddLQBUtJIsZctxBDKAZ+4zSiKqcf0rnDwnRYrbxZ9yD5/+Zm
AzTPu+obMIOzfSiDLkApA6jddyq2bKM1y4W0+TIXhqbNA6c+SGS9CXP70fmdcCU3Lw77x3ttHeWd
tbxOmolSfIy9n3s2eatOvvtXmL1LKRS41J0tNsY4ygJZkASx+yPTctvE28yOZUJGxFLVfLHYkVCS
sWKq8MNRecnREn9yXg5uXYpK1qgsg7ZjaF9sh6wArnvox9VMLFQpLMzeWBCqcOT7uN+Wt4A3dbKf
+YTUrTdVsgsfkWoxoKiAHJ6hoYFIbuDNV1XUPUWLlp/ZDHgqPcZ+ZgItSNEFMDmP5+6M6sV2OyEm
AGN3noRcKe9c+qys9YgtNOx9lNL6sw7+dFMjYU3hftv6Kdz1tgGzf/liYgFrajilKu7ICOx33S5u
RmDyQ3RYTPakPSD7WOCAF+Lq/o54htEQXtsKFG4OfXKZ4arEyv78Q57tzb4n15QmgjVSIRfcVlqq
RCx5CKf1L0l75L/874ts9Y2emhmWC1btjTZ8OWldxgJx6qGwPhoK85vUAHrdd2/8i38Ef7XXGTAH
sUkcvodAHeNRtYe1j2/YM/9OukNsXA7vjlBGz3WQZtE1JXh+H4Jxbh0wPPTdWGX/Vigg6ZEQw0pr
5OxwFonGKvqxTTzNo+Vd57daJprkALQMBHssxzcddehEOa83eiIJTwg67HwflQeRrPPf2tkiAtXC
ibZO7rAdxo8kyhw5iz9P1WP3aaXWNxokvy0cJ5ALYVw3+QWTanzt/YWJEZtjJv/cAr+jO48b5IBa
VR96jrN6AeGw+dAIt1xBHL3zKzNDQ2vdSLl/FNpz3NzkJ+vEsxeseVyPoro9Yafm3CmuQ/RoWtgG
b1wndqUaTYsKRi7jD4dn4FWmmyBP+4bWFmPDVINmXL88NDqq/T3U7HA/QWO6oy/nGRk809TfsQYx
N2ngYBn7F93XKA1NLR2KgkCju/5cnt+R52ikfCwy+svqfOxeT+cvhMPEl+toN+w0kLG5BJxuF90W
kv3SG0IuKkMaU2YWyvuvelMjVLe//5Iu7TvF2TDfE5tJX3/6/S16ElD2nl6VE0dK/QJKLKMrH33T
ihIaqyRHUaQwsXKjD/UV+mdRzPo65Svxml0D2naNKtMhWOFx5wzyAAm+1y08B8Wn6HlPXBn3SVQw
+ZuWDanGrRAjW5ZrJVkue7qZOudlWqHHvMvDPtSBC51nJQbU6buX6KuK42obYHCkNFCgOpuS9j2E
xKS+Dfd6/FdRcXZJ9fy72ZzMwY90572ESWOs3hfhbQ/4Yk8iyYA7he/kPZ39H8/N2x2TttYApVOq
uTvUkLScg7+CwdjabREQBA5dP/c1Zd3oCB+K7qGg96HwjYUXonlPPDzYAt1VA0O8YEDmuESTah/+
zN7H9yKK6lG/I3n63CmBUjNv4xCdGWdFiHTRAM32e/fCmrs+p3OGK8d7N8pZeeIw4jLmoKQvR2g7
I/zjijRzxenXYaURUz6erdVwAg0WuJcavoYpL5iazWaDQW3Ts3FCuF48ag8SeWTfAdUB0V9QmHlx
P7AzBQwAUmWThneOdn/V0UuxBuiv7m9d11tXMqse+wUQjX/tDVI+x7rfHbc+U6hpb0X5nuiiLL0V
dY/7Ag40lr0mJ1BvYIfGDoz44phj9YvGo+3EojTDuHW88zl8rlrqEa8Yy+tD8PdASvea2duBROW4
JIuQOjeKtbLnD5dkqI00mrDCqsi7zoy73YxOLZU9hRYchZ7FNtEp5eUDfCsQ9l8N+fQG9CTvUHfw
HyFDdi/P1yE81oBjlMTS3LDXt7/BIpGTH2EAFb0jgHLARqPZCZ8bd5BDjnr80QnJ6xw5p27AbN5V
MGJJXiXzK5+e2fLzSFVn6UKzoSlzxHwZLaX94EAgSOGV/RC3PjKqs4eCg4t5qHx0Cyh+vawQb9TQ
tDiKMVdWWsvZpqHLfcKw6qF00DOUkOLlqwKQ2ycabHnTgq4WCVEmVTO5RH3qN5l6sg5VLO2Yeboc
lda14JJ4LMvJ28eWqCGSoqrN8eFyNcUMIisR1PudyUCiU0bEjprCm/0pnULZElhntGyrAH//sv0w
BAR/paDloYzcC+iVZB3CbNK4RNAFLvFMROB9Be08dH5FMHZcjIiX+h6e5hGu4dWZMc4ZpXpv5WAO
bj4CzQptP6LOOW/ZdOTv4rVcPvws3TjmENTDuiz2VseQ49vYR/votgn+uBgyLQohtQmhjgvyJMQX
twHtzqu1BvcFfw3+4YTN04KncrAQpLgnPmIYV6i2wG2MOTAiukm8DsWaHS1hj6boZedYdb1CboyT
3+ey1RCAUB0DVwZNDQhZ/ZENfnye1S0dg5YlathwcdoBrWAgdt6cXy0NauUHUAKsffc6rw5M3879
mcCm6zRdnN9vl/+8kIz7ELZTE3DSP/No7IzK4aw8YLRbP4QALPXbIVmfBi1q8D0rOFdI+9+vOTMK
CoS+4boELbqg7Vk6I+UoYDgbpM1aus184GYkltr8mlMUesBhwbew4n0/HTnE8yjlx5pDJ9meOI2q
IEcV6Yh3sQ6kgm2fqPldMsxByWHov+/H8dC+jZvF1J3pPdnCkvL9UdClQWp6vnabe0it2Au2Uoqi
83nmUotzaXUcceE4xqcxKf22zOJLWw4+woV+c5cZ8kWINKikQDa4G/yTMLlzhAReTeDqdAL4K4Dw
qFfGvfdSJS+Wr4Kkueoknq06vP6yTP2l7HJQz3fX2A9sKabMJzkQB7S7qpHroE1HBwBVuWrdPPt6
ho55rxta2e8UAw9xKKTnOeLLfuPchzKkOyb3aNkevVrE2AXXztnMrWbgOzJo/D7+wYPiplJjz2La
kxCOF/iSw2VflsZbuuvEWKGj9ioBxX6ux0gZPHCN/QcWfm36MhWo1UnEz93P7rUuqagod5V5aba4
GgCP4Xj++/o0KRuobdkBW5gkknjPrthrdTQyboHhPkADHS7nrMavuHCVWhpYWxTzGXw4KGZEfLiP
wDwBT6HjGEwrTZlvco0Y0oncDGtFPjCs3QkZXmk3ViLFZ5oF7o9cvu6f+/QrFUeqMszLyl6YZZxY
YuyP0uZzQrXdp/fli3+FUXpnsVSfw61fJBOWK1w45RZnGPpu3LVxJEvJqYvP+SCYnWgmw9rSv5R1
Ig1JE9NgWMBhxR5WODOMqgP16FRvD/e2BYVIddFjOppMOzzAfiIpNwoFw/kAzulKuoWRqmsYpn3X
5mQBFL9uAwvqpt9Hv4VOxPN9+i1OW1WZzdzWfGm76i+/HbT02EQeh5mFzH4DcP7Zg4n+flXG2BDH
M9JQ6Wj4gqhAH9ZFQRG7IqSEaV6MdO3WHOB7PFcihjvjnzM661wB5ivZ7B4Jl06GFsQRzYDlAX5Y
7xH2Jj4w9fgnP56d8hJeGAoStBsdOR3R8Z0JhXer7LTcNPs8tPz7Mn/jgpVOBHPQEXjJZCtxsIvz
eYcof48HPQLl/Nxsk9CB5sLTftK/8Sh4qx5W3PGCu2pklNDzbpB/gxy07BqAl1UOEjle7FrRKwA2
ePVfCzO3YYB8rLDgIyREp4fi1iezi/+4QzpZP3OuwOm5O1qXEVTqIdT47VgcwFXbnl4vdrROQv25
SEPmbuSpQCcWd4m9p4gXYz1+CWwWhzelquhEcqZEOf4v8xTw3ogGFmGYq/rkDJ1o+DlV7WDbYQnR
1qp0pbevKcOUs2xC0tbIwWfPPfqSsrZZakOHGc5IlocAdm/gey31WeFu9saJ9bvHQdVYquAcSc0B
B59wD88LXZQTfs31gZWTr2gv9ChCGUDMU5DscEr1b/u3NOMrxe3NO5Cql2i8dskkYlgn8HLonlim
9HWsarPA13xSyjTls61Qr/+i6WuMT/VyHrL3+6sWPSKqNZm/jMOGHmONTrd1UpQT8o3kdEdMpT/N
kMHgEL+jqyeBG5jXa+YWkcM17A1Rd1B5LeOPHI333/ssIqvI1fbCkxud+dTwnvXw+KQ3F5H1i5y3
85VYXQekHtGv8iG+91PfTQdWBmKR+ZfiKX7McrKqStnXny/L+/qG0uNEuPBkILP2Iiaj7aMYxDIh
UpQSW80TxfOoy1kbn7ZyVXMGDF2M6UTMDwGp2LoMv5ae3xeU0EKlIdx45Wh2ra77iPtwLSv07tET
1Sr0TIku8uuXFNTe7Q0QGTY0AtH98Dg4qxYkIyYFHtUNGZ52suTb/Kclmncgy9kBacwOuLErzMdd
eE1uNYnhi306Mn8Jw12xwL7s1LfOwr3RM7eKySQ7TGmx4qQFYmzB9ZYbH2ZXi9B1qIdCr57wkwpO
N/iTo1kaY8W8QTz4Jt2/9vDPLQ0l72GwkiKdJwu/Bypfst5eZjvEU2ZSbj2qDEws7joySbKCXhCV
GEHBOfPmoSMNNsoXr/Til71FLw7+pl7W9t4Ek83AWpjaz+LFTMpAA+bdiEq6gCrdHc+LbWQwKqsj
1KOxZ+OpgvfkFp+hLVsjUB8oN0A0ynC522/faZNBSw1EfHwtf/wI3qHPYXl3GvoG72j27cUbqG4F
2P/s2vABnIqLviW7HLfOi1Xz7ufGuHylk+t7MvmnJDidbuzMI3PUIdaEzzEgAxq0IFyvavXdnivW
ZEf3k193d2iXroTFGZ4hzxZYlTJBAZJdwovri85lhzglQsAcuoV7iclxhagBEz/14Yd1dRwwlZ+P
ogazj3u4jnQoc/1Eg0Q4eQbrm8faAzDt2Dsp62bjXmDy0WLu5wmXRvTdOlvWrYMKz6J+P4exVj19
mQK+RK1h6aBKCUvAYHbId9kNkrbP4cSggNQfs3JPy/UBnUvIVx5MaVk+viIFL++hTQptLV9nMh5s
H1oCsawrohlbcAFz8ovFpVK9qpz/ep2I/lmUSafuFlgjoJDVH0GCydQ4phLzVFw2VQBYGTMD0qXO
Ay4pn6NkAcSeNh3l1gV0F/MSFDxFyMUUpFWMlu8fPsdfeCZb24SBkw5UbAiZus6gllvxacIaE9oc
3r39lssUHXkAx1C50go7iRDRr8gBMy6EoovoNo2oy3HwDljoywWjR/DmmULSI2hCiyizpLqUZ074
x9FZWbkHGoA43BhB2qxmCu+hAqdZjUGaNxaZkcRxPNyBUbBR+sMvvyiDNiVXpCeSoZlOypx+MKOt
h5cJ7HSW9eEr5sdivzOdxM1rXpC5ZbmGaR/KDPpLSBfIJYSZNhvJzbe0Wo0MBEb465dUgFG3Ix+U
S+XNhCOgtZFmS9lJyNJJVCzunCxtPAiitp4OWetyC+kfLsKZErdxuayn0JuE7HDsvqGA+lKMExV2
yT+Pe1O2nJHGN0/hGXuoIzmc840h8wTxHntzWRVBv27OmEotkafqUpnpykI4owWF9WxOeaoUPrLY
/f3c/1xZWnDwCylxHl2eDPTe97CvL0KcsIR8NVApwgn9adkiE2xsLbi3/n2+aBF5fdwLI7mbctLR
FMAGrSySWutp2AOpzU6BF8IhZKxhfP+ug0OLJwXFY675s37QRO8SU3yBYA6ETFAndOr5o/pV9g0p
T/iIzBd3ucIzj3rqCA1xJUApQu/oBOcsFkbHK5MpLDF+bcQpBH6ts5+r2Bd6GNRUlHRtnag/0mXF
WZJ2G+CPmY5/OcPz0On+dUcrYnxtbT8ZEPQ8dLr9jKdOf//SVmUMa0FHDJMz7a3dEVsr6AxEi4VO
tCF6HU0ncLggHzmKRZkJGEQeKo808MHrtlk6dfjs/ds/AJvTNCLPYk49SJYLeXOQt+x6qhQ9jwKe
HUGOjSA8GzRVfJGMasvnWUUc9ViBqraWFG7ins27us4NNx2F8SWRu9HAwLsVFFkXOM3gtc9ZTBKb
+kdkDIhPFK3DOsTgbo4T8NltVH6WVAcl4lfSa8GMZsSB8qXjKmAwMXQoHBNSYLP1xjQBadsFqEj+
BTCoQdL/vf9AMm7qSjkVzmbg5G6iItxmmT+Pxho+yGG/eycmRM1ROstKXqCitgG10jwHWEsqr5Am
IRLLEvdN2HjOydvUajLFCkrnexSsLM6KuChr/8IqbxINCczEzXgiMa1uot7ozN90n0n+wPbPLek3
UpGEYqzbYiF/TD+aJ3OTqMnf+CYabWDSFPy4eRln8m9oNnuci4fd1BGxmsZgyC6KV4q7fhTOitfG
jDaOgdj5Xf/FxaIo+EY//a5sYkcOmXXuqOvTo7J7TECZWBXuTyZIPEAwnL5YF7QAyvzZMQVqNPqc
S97Nm8tPJ/+h4JzDnkq4Rv/LQfXZOnXjTGc8RpCO1fY6qnK51r5c7QARC5mYnyM7utZfV50xc+is
qbM45SZ+rgh14o6mbQdNbbzXdBfItdfwe/JNYHtN4ymlNYoLpYxWCLhO7Lgf1O+QT5LMCBKCpjZy
RUZ+sJnGSclx6cJVi2aI1U3FY4rj5ox6t7RD804QSJFupjmeQPsjbv7w+QN21Lq92wrohAE/CRw5
8FRqQhg6GI1VEpW0SYbXQqlAuuFdz5DkUFxZwPXrK1S1fEXTwbTqQLIE9kHmOx3osL9aPW5hZNY5
rDA8jF71rVrM6DSjE819ga9dNJThAnkFpHVlG2OU7SkrW7Fcj5JHqflOxUZAzS4cExLss9RONbHy
hEUsfrDIxKEcXltoa84eeXVN/D2iurUL642GMsbi0EKovo1ZV55NGEuvaHtIqq95t4w45uFpgedY
IdYRCJxqpcUPo5gwWc5ow21Gh6Vb04mI4lkeOBTI8UnqkzmSOS8e1o7K2X1n+IF6cBTDlw9c8v9r
91oaxvxS/y+0uCik7lzi2KAQ0gKSL4zN8TZWoV0uXJt8ilNNpwJ2ESGvXHikqtBJDBZlpWCe3Xuc
HueJV3W2L93Aw8K3P6Xzo2j1pUe86NOHeNlNaIo4sNjudBV/aNDuGmYeKWRfa2yBKKdZWz6/V+Oq
xrfmQgK7rQoAX16QP35lD2tpwIJf5NUolc5iGa9S4616GzDzHiF9Ft7qP2VcPNJj8GxVNDTERBrr
jecNQfbMVNKI0boe/MTznanMFDa2dyMRQoKuj/Y+eGVFo3ohbNVgl69TNnHBwMcyGrWtbrBZpUoV
IIqGXwPKK/X06gxefkOulBIyOOLCOLgyFvxjzqYqPC5DPSMyXRjpWDA2wBcq0oVCu8UwUOenbPON
KuRLH9ymqx8E33nbwZp9aKuz8wpB7tM+fv4d5ti8EjbhmHgf05XSo1ytRuQiN3s6kg41CbIPROva
dViWOdqCC0Yapbg1d1AlcGvpWpGO2pAGPJFfkNpanPjWEx8NwbVmb+1+h+WhGxXOiBKpmZjfShhr
6N5lHmYwJ/EICZjgUZWPBhPYEh960BpTKFmzzNAwGHJUp+bAZ4cLr9hyv84yKIge1XF9D0ibjkT/
TPPki6BWF6d1NH/yK3C9G6mk75xWY8UHqNIWdQBgLTmEtqEIHVvMqrFNaL2Y4ga9GlWCKSDBpMQo
j7a0vULA5sKQPttD4U6frGExpLfpzEIjuPCNeIMwEXtaZpqouC92ybgbtXXg5oWLTnmgVv95Le6O
KqD5g3to34E6VxYZDpsY2acXaNsNyo6QfeuYbG/958/qlOKjzkj3NgL5IUxnXVQXuIHWpbAGkJvr
CoBPROUA4kFJurjkZLp5Qm6gi6QlF6GmxgjCVk3RVLZNi5Nyu92HE/iuj7GLtb4+q8MCdtKzVMB/
M9h4/dY6qf56hoKFqtRoB3uhSPpC7DFbUD5mtZi8x6Ml6DDX+uxuQoNvCJ31yyltO8yYzf1/2i/F
HYNkWMlXyP+zn7oDd58K9vHk+/RuMW9mE95MY9D5Fpa097eLjo8/ugObjzqyWzvB+xsuUFfN5iJF
UtGUM9mNwyw1bUiCgtjNTnEYFUuf8l6BFMnIpRiU09U+bTJ8xGEgmFrJ/PoyBuUk6oc3FVYwhEqX
EXRvRzS0hUuvBdjJpta9H5yAPiYzgTTyQjxDZ1qSBz5xmrxeo1bDPnNMwiMXN+3Gq4q7031KzOwO
gzRB1oLQ4h9PtDdpXQY9DQhDFmWaPVnIQ0uFYUmOJ2ot1w4ZTNQ10osKwXHpA1occ37kzzhiJ0RP
54yi65vL8iEvSwvmUu+PF9IMfX1FueQ8Xm3WVP5qZU/gYNIJwRtqnCvGT/93msJPWfsaBl0mGwN1
U/xa7WctfgOKaowHF8ymHqIOzgRIyBw6UK8AT1qCkhUzbguH/nG3wx0SD2XZSrHxt9i7w3gLZUfl
7R70/hVfQPQmHI1vTNzTq3hKdRZ40NDGCA6VvKYrRcQpJtOfGfRKA0hGznWDWX1puj1NQD4cxqV8
b62ItSffHLmzkF4W6dJru0VHTkYCOt70pOts9Voo3+p7MejnrcQDe4EStP7v4EQoe88/Z86SsQd1
eEnymc6Wr7rVGWBvwk8LYFParJHUC0GidUtMKFNkDJ/4VJ0cerFyzPAPW7Baicm0Z9cn4KgrqDs5
B7g7oSwp0pP3ZaXq3jZSZBnUzMJHapOW1ItuEhMu6PKKPhq8PZsmcfcCNZ2ATRK+WfuPWHr29vuV
e5/TmaXReRH4T5LQCutFn4w7rFjx5UCoHFanpMmD9vpwkKlyMeGpmIpAM0qbiX6zc+1S3N/8KYaZ
ADVlM8wn/OwKMwny0Ax/2/7qpGGpDoRZLGM7yBTTurydPoAr/D2xPQeb9i1SPcT+7otVtNBKjytd
tNvd86/jepdOV+baMkN4eK5Jokg30pBg5Rty47qwsRJaA4O/kJCFZ7Wngy2E6CraCJu48GXIOS2l
Ha4fIB0YeS6GxlHS7mTbCQr58Q/mLeDdZnHPm3TKSsS66thXHQ4LXqBYrqcwb5W81NrvM7H2mx7f
vMamS1ryc8tsqDtaMBT/lBLfF6c1H0sHDIXGBliyDULTaWqZgYg0XGeLDKoAoiyptFz+0RmIbzBS
OriS5r5jC28viRk+M+PGyjBZrMBdK0jVAb2f4QB1JwM5ywMT6NMeLrimfruU5fPtZWzxYbrTJMCn
cXgIERJ0l2woh4Q7F19Bwys8qJUYbbih3lTLApinjcVk2/qKPkWZmJN1zfK/kbsEelPTjk7C1Z8/
pVaGa9LM1hDW/Ugbo2zAvAcs73jF57z9vLU5Uvr/3laP6vKT31SL2bxTy1HXLfnOa2kjKcFxv1MQ
HXigp0iFweMbhyb9mwQn4VIZb44zRWNNO7+OuILDjFroym+MH8FdhuQOhjuDpwgnbMc7b80c4I6V
mWRUuKzFa6x4y+CHfyBA2N1PoY0nvA9QNpwoseopQO7Rre6TeJX0qjTEseDUqXnOVoUm7q/sSrgo
pMJpAssVGXx2v5LVXEgZALRI+NGqPSmF8cbU5zECiJjIAhg+Rv2RueC/LlGDCG2d6sB5NlZ3flt1
RSrrXEzTpSioHncI7Dt1gOWSyjuC077j09VZzBSgTk2s2iQTianpswLCfXqoPfMqPuZT7k53FMLC
LJQxl4pFWz12+qcNWYjo7uDPIaqkIxQt6RnTow70xo6VqEg/A6luojBkm7dyN9bErYD3Ht3h7nij
qjV2JNwkJ/9rw1wE4xd2q7cFVUHwwql20Jyy+eHAzD/+IETn4HT8pZUcF8/l0vdkWX+p5taOGQJv
uLSRWGsQm1/SL97CaYGs0VWFC+n+pbWyKe5joE8BIQ62Jw5DDzgc6RNUOM5q3wqIPnYVBH1GfkF7
zGQ/T0XP7neAiqJQqo7WawmFgtIGJ51Fp96RA8ov+SfewgWqlDqQihxb4L8U7v14N89Um0/Ok5aQ
QmWHtqhOQ+MAa5r3nWBp8DyZLdeDmaC24QEO1I+hXa+XCdYYa9itioSaxDyidD/kmQ5zsTS5hFH6
eEsJ5CqyLIf2qnfXBkALmcv6mAbItW0oNY6AELrlf0rWYPqbfDMCxWY8w2r5p20PAMqoZGwqw56q
IZgpBULT4clouL0mZWlny0fMyI+OF7yv6bm0c8pSICKBN/D5i2SMVB5V2YbMUiwL1adtYGms2IFh
y3uzPT+KGNb2cB/eNkGzsySK6nSDx6Kk79A9D2grmHap0/fe00Vi5nliwoVYNBlwLhq8CLWbmXeA
WcGBbi1BwBQYB2GTN+gR236VdCTmjaSN+O6R8Et9MmuhgHsL4HwQyqFx3jTdbDGfwUzXWMFp1TPQ
lvqLEITBSII2HbvJqUBi88ra2WBHv4RG+MAxjQvbfRfYoOPHfwwR7vKnyZcmoqTxH9iX9U+gnxj2
YG0SKlvMACQTxmUkfgYB5ratrA6YYEDYgwG5KQBgrT/7w0TZaKt6xnQ6SUJ4l02zZK8AdDtZ9JQB
DZhta2NVysMPmLrQoVc3GtNWe/FooWen2HZA7q5K5TEmth9TUiAQ1rnwGzkqwgtmKt5S8I+IiW+x
fDJiIzXFirKAdqriyT2oVba7gk5WHajaybD50QxGmBI+m7IAZM2T/eGeN8FqSdTXXYri0iCQxT0M
y0ejETEK+RDJzSB8iSRQyck8bbkS7uiXXdPAOCEeb03t657pjyguyzhPl9y1Mhs46MBWhd5b47e4
p1ZeQ8xVkP1uklV9jPSxWsCCX7Hj6nnNuTbp7k3EaP+r1iDepBbrkgtosV8ZGWMDh3oHdcon4fA7
nq8YWsqNrOiC2nGlGMEmLqsOuScIVEjtMBSldla+uakWWtHBKiEYkKJy/K+moMotBVTmzAvaudW3
srKHFXzNaPngBjfwQ4CNTRE6CVDhoX9wOoFdPpLqGga/mvkh9cRHi3kqfHTrFJPQXdoaYH5hP60a
ps3G6dL2X03bcBrd4OhSUWWY5lW4G8GGMoF+Y7G0FzuS+ybOnM4RniEPALXEqOKr67LxK5J82NJr
YEDoRUeIkmptD07tiHxvrkyf0C8HR4fqQdQ5oHZEauHFBWc9uKX4WJa4X6ngjenJ1v75LjXDBnm6
3Mg6H+tQcQuhdFZyWALozYejpCESK/D3C5PrxIUdb6L9s4OZUwGffPUywkPK2MZoNan46fSNJIYC
btqBGEQ3PuoNKna41UDeXq3HGx/D2MKtxP0GlVr8SLWpFpA4BZ+tGAMtLgGF0V/JOfdJciMrPTod
IkEj5APM+hsAEw6qLVlKXeeZ+6z6dcSklUj8cTFCsF7FFcocQQzr3D0CneeCGB5yDJ3wC3rF2Ovy
idRtqQvXkH0AwGROdICoCFMmtpmvL8FrjUwiefnBcBvdAuGdZ0cEld+QV/6gZYwazn8fRKnT/Nvl
trL7zkWmK4SKqlDQ7QdUEe9Zc0WIUg7BYNfkxqwLi6ILqKY6R9eel3yMUeqpbe4ca528Tid0FJ1f
z8fNuJWZpv+MrYV9VWZ30TRFDgr70rWX1xQzMjoL+3BZT+j2p/fWqsFtPUM9VQ0mLaupv7adlm6x
6njtRD0s/4UJMJEODn/9OEd4/1Vp9uDlNl3dNMRE5BYJQB/oy+PP/wvwFSvjavI3mfeEExtPIUl+
Rst9Y+vIbvBOk/lEfscvkDDZYMTVhlLH4WEBknVO0ei4//aLKDi03li1nkGRTOlVXVv8wwSY7uqf
vyAFbTQj8VYGTlVClIOTZmTol9XDenZM3Eh9fnJxZ7aMtaVH2U/F/O1J773VnrYY34i4X+8+e2Y7
oC1jRE+N5PIlKOmsi0AGV/E5rrirQgW3rm1Memu4L0j5lptC8UR3cS46Vz65Yaxzz6GabdVsLF82
tSIEbbHwqMQ6gVts4YYy7RD3IA5YF58zLb7dcXGDYGU9VV8XUSLzF+6SNvPjNt7rEzlGatUVITGL
6hRyeLqPMjSzhik846FdmwxgOnsQTzfj6Zf/Lp33ogM6TYHFtqgpOf+ou1Uc8K/YF5ERcPZ8ZU7+
Ny0wnaR6E81mRvbN5QDcU66KoWgm/glVXSCuVlR9tr/IpmkR3m1l2r0c0rIKxzBu7zjBSLdij57a
LFPfrZVP6jbBeIQqQxGOLxj/MKkB1Xki7G4ttLWc9Ubkx2P2UCcLNw7bBBQmce0qokEe9QH9axCb
sA4YzIVRnKj4OLXuTrJmZzCN/0Bhe+hK5aL+ATTcwljA1unIOoaVRbc+I0K0n9hhG/JRyB7001W9
9kDUb+POCt3ezf8OP44qT0Trft2LKf5b3IrDKdAxVFbM6g0cJV53XUfCaRKuGnmtrUlF3Mp00ID+
yh/ntxfwhXuNWmG0uSpg4bxsIKoOzZpKYWslpAZxorV/qJk7yiVAq5slVrFizZ0JXzfbLrMvunlk
VuoNviRyhXa9CiLD8UaHarAMxGuyp02NeZkzmoDlPYLTOZtvpK3Lb22PxVkq48GdbjPBwgVb7NkV
wRVc8VnQpUZH9LW0nyoOiJS7YG9GC7sTqarOgqrAImLohfxlegUTRGJUTo9QDk0SF+lQgsP0LC7C
INs25F0oAZdXduos/0Oy4H2kMCzSh+IRoS2mt7H2NDvkoAoN5wCnHMosz3patCOxxIUnsoma12rd
70OT44k/zcg04gXNjJtFnudzexSKXkrQB9ZnEZONDvPqLriwhpqCrVkLZ/mmn4loB3RMNyC3qxuu
XY/zNFEGgvcxrnU2qDJ2ENqj4PTL73fUe5o7maaU4XniY7i8echafuDYqJrgoNBq0tmJ0G/w+6BD
9A4Me1K9t7wpKeASm554dBKAHi3Vj86iQyOUzwMaw5TxhqpSB9R9siB8VnwyRqGU5D2EZ2c+glTN
NVoGyvRvXIPSy9NvuAj38hRdm3nVdSK+WuuGCa6HymLsEh6oLS6Ag5jN6R2ROWiJ+fZGNSgUyp12
2IWEfprKaWrFSFf2tzaYFuMVWVPgg+b4JiiQp2ffPIsYcuRkGmoFrmWiJJte3nMHti+ojJiqdMU9
5MUjOHOwLbNOn5eID70lTVzgVezZSxcP5RpOd6h6Kf5qt4oP3cxZ5zmoDKETElZOBpYqchRhQo5G
7c/k0ZgWkqxvxNBR8x+UnixcKdE4SePxXnCtIy791lgmQ5BixxMwIiXuYgaE94d6HG5KxOIYaRKM
EN2U4g5E+Q3U4sDxpEpy5yH2eQjRxR6ZwI//aNLdu7pyYyExoHeKFeKflRzCVhNC4xrp4A3W9wqO
5BjxSiBPtWgm1GMlwfELeWeDth18WtOanKkMf6OkMT4+nhD3WI/vLe6EYsTJlPJWcOA4uphFg7Bf
Iu3pYAJ4EJFzKx3Lbj35iD4mVSAc0Xv9PIRIH15ltDEllR1U0PRZf4GTh2pgRT2Q5VQZa7C1FCM9
iZv8QCpe6e39eB/WmHy9V47sOznTjB6iTCwbt90cYfqkJkhUA43Vr4pyY3CThXvZ+/jY8X+1rRio
a7y4Yj8X/GLY6qsv25XWA4RWABgFJKgII8mEQQF0YeUcdsLTKiARKG8cZbLxDQnnMu7rVsEXNbPe
HzVsV71Dn1Ga25xnVXlHmfUJ87gQBM8VfAXvJWrIkd0KrWqQYRDP0Oel7ykTTch48POs6QT/RT/H
5tM8xhJrn/yN/h9hSTrLAXHhGInCoy2jHRaBydDSlsIM8sDUPd6UkG8O2gED0nJJVGSeLA3wtSV7
KQ+UbKGwVoo7AqYMPhRU8Y0sjW9ItYeHAeQLbmbEDsKB/TZdjh28sTkLbsxQNyBaSzOxkhvwshGR
wKbUDshcGtSiH+TWs3I+Me00LqAfSez18u3PbYgMnm1E4mZ4x7X7INrm6dHuTB43Zey0ysNYdyMo
muS3GMbjYwMhh9QGh4QyTCavONFL8POWuH9JZjtIl97CIVEVCx/PwNSvshb/c88yGbBESZqbUex8
rTMBSTMzV7EUPSihqz7qZOytXRJOJqLZDZ5ivLxhaw4+b0PEYsuz8Cajmw7xIB4GP5NXKJ6g8tdd
7R+7Qzu+Dadg6a9hZEQdvHlxsOuxtnGLc0pCMjFx/UdQ9QwGPZm0jgz6K21GG21B4V9MZsglf9p2
QCH83ckQ5ibY7YL3T4osSCXjjbHnfu99K2ddHEkaGwHImxvQoa4Fv3OQth/gnleBJVhMnQAbyRYD
Qfq4Q2iPbUVSJuV29tSGQwn44ttp2AB3KHyX82DFrM/x/9uxOC0mUrFPKfYhrNHKTZD0fgT6Owus
+cd1/EJ6YFP+nCG49eDFEjMKz1YnxDZuNMkd7hgDq04hRX17UA7GGzUmMkWTiCzjVQmRX9kfz2zQ
zLeyQgMYtkFB8TJyBDImrCtCdi9xo/lKzJlOJ2oDIe7dJyi0w3eej1M/SsTvt9eBdxa9GHOjYBat
K9fwHKvlX/RXmEWZJO8lPRFSpTmtu9s9VzyRjJCFIz0bbO7J2ychbiKsnrxSVcheWCByFRVh3Akn
VEtTub7GQ9JDb3qefPTvUuFMObhCtWORmQp8WEjWZWWV4dBKlZWzMeoSy9mSi5Sw3g1+6VKsHZJE
FSmPpYeCz/4w/4fa4DmifCBDZ2eowWEoHFeyNgsvcE0tQpUDBDzpBpmFu57nRZSG2XE+QILmRqtV
xvOK15pllgaLxNVkB3QKzkcrQYtyIzbuasZkP5K210f53In5c+uFv67Wn+UCwAL5GiYUOXStECuk
2ZkaVHG2xu3nRtgFE5UFaSD+eB44zqvh1STjXzNf6+OFdHXcJfJE27w9RIB5qJco51i9VnQm8UUP
4JAJ8/BQlvGrV3vtGzEvyuVDwfRrk6dg1rReS+J5mgCJM/flqQfoUB0W2iq9fMBZ2p5J6ObBqf4h
NOBlVe78j3UNX0vSVe8W7rPaDiJLkYge8lrwqvGfZxdp74y8r2cVz+rMxmLvmKz3/TaUjqxsFjfU
Kx36qQsJ0ZejRftNOi/EfnEbFZM1Ld+p091xlBL+PzZNtZDA0L41YLMrOl/BIoZiM/Caa04KifJU
wDiFSRB9PYzJWX7LYKWjkO2cS3xzfccRDnc/1fF6QZQr4im2TxNM0kZmKiYUW95B7Qho6gyl8wS5
Xlf8GRN7RsJfCp7agILt9xwew1cQn0GvPqI96wmZTXkvpHmpctjnY74QGkqChl5e5L4UAQoY7Fip
CDfdq9xYOEDKCiosU/Kfzy7vH4cxmQBhbhYA84uw7g5z5XTjFjki9cTnKGhorMfWDP173Y4WbH8Z
uVwzWZFDKxf5OJCIT5Kn6c893j+cPHEwMllj4xMX0F1Vdkax4XuqiXp979h25qiP7s97Q9tu08g7
2trwR3QshONo4WVeQbPwM1saUI6iNnEcClvs9hyFbVt4o3C5RRiFXXJCCx+RgFOgr8V3ei1ow+2A
jwce5+57i99ztZ5Om4wqXQY4tABxEXAJ+x//Gt2rS0vPjVDNQJXUfgRcGScj6DdXKBTZ//7odgpW
xUQ29K5TulM0BdGedEFaucPmqnbviqNsWEi6vaqFQJh9JYHlqfBDy0cSDntEp9LziTGGiWWD5VCa
6gf4s1e7JxbwiqZR1XG1orI0x2KlUpVDykqataRoWkEZd83c4nNbjoHmAsvDqG0N6QrLsMsSrG4H
qG3l03A06SkkX12l3r2g7BxO1xc9pqhUZmhkTdIkQjR8yECBpDSkVBqfeN0/xLM74Or8KpmUNEDD
izAfZ+snunsnet7xGy0+yKxS7VoX+E2AodLIMTDF4pNu1q6vaGwICZYuWZ0YAvY/2Ok/rkiFLVnp
9w38dSlkyUggjetG7XG5qonJXq1lpWUBIRvUj5yzVLcVzW6LPNaZO2FVUuQwLFbwIf1TmhjDi+0E
7uYqzO8Hn2RO88TkSgH9aZtF9hhP86CV4qg/GhKMlEIOKdxIZ8J0JpAEDga4ZfGBOxxT6yZ9aiKM
RoO2VjpdN2uetqWnWU5v53V9Nep4QRrlP59zEYoNIWZWyLNNr0mbbEt3jQLEIeikJekIfHoTVZtw
Dqv3V2thMa6FNsIbJR3QTFHR+dqp95n/n8XR4REz04kXVTp2mq/LC2cP+iOi0GAW3I6mG8FYAatK
0IBR90FvdqmhDbOcyJQNgyzeMUnjeLGMpIHhisyRz1UuHqnxUr8Lwg5Ahx+ugLbiGKcS1L8lgMZK
bcabpnIZ2iWm2vt3wdLdqU6CXcXz6Q5Etft8NAKZKlIFieoZ4rjbXZMr/MavwB9F0GN7C7dW7CAQ
Gn/+ARzi87hqHJQ/75W/egkGbAk+TCzyHPd9MpTiyfBURoVRZl3HTHb/sOEwm0fdbd9EYv3c4YKV
B5mGbgcsdbHZCCFnWlGh15nniJ8d22QofpdyJLQk7GfCF8kqAFFDUIXtQL6GryZz19hBHaYsdwds
Oyec8iIpDBw9UQp+IuC0FGYWWUn3uTOJUxcCfX+0v5h/x2s+11S4dOSuuWZUj10j2igOIeOwzJ82
jor+Z4b8EbtV+kbcyKhIHInbCvKDdBKbaDJmnAc3qUQq23Q6SX0UJcYWydd0W5WcovfDq0YXvhuD
lXNv8CK6ux3bBlYzHI776PjcWjk3HvQH37yEQWA9ML1mcvaFIIPqZodwjdBrMYqM10i4Eqri6ZpH
KvrHHXCKUvp6bcSTKiMm49ei0JBcyPOEFAoUHjKdcZ+zMK5x304/oMp09XUkBN5R/9GigleuXM+2
YxDIk2tYZ0ai9TavSE9C/V9lQqnEa9YkSKbR2BI4VyAz3HHyKeLXtiYiUp2xkVVqtQaL+FnQyN8E
J/2Bd8uOTq1p+ufMgjyX/E+L0dP0roWyhDfyCoL8m4/TUgGQUyAHxVdh+1+BLhpnArJQieOA0s8T
J/pcWl0Jj4VtMDXYv0WxWXo/USYwpykjAbrrUq080bQ7bL0se1fzwioeh50k0/QumPXTNSt6SImF
V3EYc3FY9VZks4O3v+2n2uuxOm6ydV4I6IZFHmpkyzGD4+GbSPdqzt3tpOJv941JGTfyZknsAU0H
L9JUQShAC6eVnZvQ2lfns/I9XXSWKNLFhLUx4hln1ukksp65liCbg4FRlwpxfrBtE5wEkx+chG5S
iG+UtcbHEUREFxsKIEKtIgXoyaShYGaTIYufjlZXMDGLXEX8trqLjcXXLrxS30+I2Bjek1ANkDG1
Ow8dNlWl9x/4a3YxZmckcMwFe+5SXAETTUw+jFWB5iGFBqDlEgjEe5E3q+xo3WKOxgQ0iPLF/YiX
G3CLi2EE86K5L1Jun70ZSqzCyQfO/JZOTs79+Woru0LAsj5OkCJ3aVM5ZLGwsouBhuaG0xJTrXJq
uyWD37rlN9GSqh1GvwVvk/QJ+OIsYsRk86W5J250JLDzoZMmu8Z+xM8dINY6D5m8aH6nPysfVT6F
slx5/fIK0i0d91/5hcJmirzEFr/pRMzve1zA7rxs2Lw8D/5Fxp2ZLcJZEO5/62WVFdlRvbgh6wbR
pDjhbkDQjGPskQ7OO7emvFiGaRjDqaEzifnFJ+x45fIOZhd9Fqsln3BjDVEpiscwvg6Id22EZsna
Rt9D3mp838PGpcnaSRXg4iJLhykVHreiinHaW7EM0e+FYQy82K0hUC4RWVipP9kfrmx9SfJmr9OW
L0Pkqwgzq080CVDm2F4CKGwooytR3YZxaNoD2GA1Z84O6NduWxdQ1GmQAARxktmNcHRP4Cqi4r8B
SPilSJ13ezvKBXZlCOu7sNvS06ZSKm0XYnpVsU77tyq877yKhh/FXR3WZowNzfWzagaTAqz9AD7M
/pf//6MQPe0IFr/d4zxuMyqfVkcuAYVvx5QG8kv+aO9Nuj0mqr7ItzY7L9CGt2xDPX/0GU87ZQsc
hCYjMOY8fPCb65vDKEsBVcb5LZ0OR+FENfqKvR8Ksmw6+BYmw0QPQdi886nBLv9S391oyKIkmRi8
roDTiaZe3IRD1sF8YPYYvTAYhMmlp7pUaIxTTTissBqx/a0eEvbpsqYIbzEQaj7EqMAtP/Y9DBM4
63hfH2stzS+SK1nAN/EKK/+duzzxsBoBKshpwcw+rCi7Icp9MrbcRtrDe+Zn/yAC7l0EFH47v7x4
SYh6ZMAT93wTn234E01VxjtVIXbos3BPGt2xi+KEcetcqrgY7Ka511gP774A8GDUzYT2VtMZGpPS
GqezCDDvVOokm4bAJTpd8+MkRlgwi5VUlwNchxjtwqKaqLpvOt2uYzjNY73Y2eOKx8TqfnpE/WNa
TKHQlGpoj765Cjg0V+PsUE7LJQ0yXRfj8r69Y4CSrjZAges0TxW2enR0u5JCbeuv3RCQo6zPNLPR
0znNkwuVWJxtSMllkOZiSuE55476tYGQAh8JCzCanB3pQKk0WyPLFQ0HVAWsHlsVeWdma4hI6PXf
4L5lzPHgcOwtUdLGqCFGfvuucpT09/0NSMTZhJA1b//b9TEnwUd9JhGsTr56MKnnp8dGCXfTHsrT
fC8b6Na3ZOpZGXDtTc5IsljJzu7YruiSAolfieP9Rojv+NceZKskZZnrZAk23ceAGrVoOJ9zgbsJ
UkRHji9Y2EYKfiktp738PnmLKUAoRnpcCRQPyqKbyc1suaNn4xggE2JCQXDbp10B+0j9vRW9yvAN
N4X2dYsaRjNagPW9HtmPvsSlKeegO0oOyfdapt2PE4ylIxnQVTfewqYqH9xA5gfWTmLoz/Dp07SP
WMCeJqm2FaYJrHigP7BFlfs0Xhk7nPr4ONPwexa+tP5i73E+Ipvbki8aHKMxzWNQuq8wkr6ToR6C
AYKf8oPqosN1wXPRdAq/n8GJjsoPwAjwOJc4SGWKpn62cwirEOu1eWxGRRxHUU4VEH9ee6p21zH5
lXqnMDlH1X/fHRkioMy2KAVUluWeJvrbKBx3KlwoiobuwLmgMz5q28H6VeBuV6h5n6m11WDaGifM
PKZeuBVr7qxpG8H/ZONv5gbLsDCmCdY7dHfgj0+qxuGV5+FAOR3X05SI3QsuDcBJ15C6wycfP/GZ
/40CREgD4AhBudUbnF5BKDGeMibVv1P+1nDq3fkdjFCn6nc3PXIL0MHI1YtqGoBkaXt/1eH7oDeU
FDi7hERehp9Z3kDPn+wCb82NBLaGYfEPG51sPygPQquaDtiYKhwDvAeuRGt0pGkGXT/1qMhx4tb7
/pfUex2Tw+M1DdsOtbQoecnMGXjRmVXOKHygDQLmId6TXqARxYZGPj0rVm0SXw03UzD4sfzpVWYt
ICxojM+ST6M1EKoBkjzlRXyok4YpP3J8JH335lNhJhmzOMmpVbp2dBO90rDR8xPjBib6bZk/Rp4T
190TxFm77/LGqU+Gk/JpCtd+VQqrETWE42wrreKbZUUdz0mZFk489FotY4uOE5BhkwhB4uhHcpVf
cmcVhB4nKheU/crrUmbr0B6cfblj6mbdW6XtJ6F/ZZ4sJBLoZRpM8IAboR18blbCMpQkeHHQaBtX
dlkdwSqYLgbvIY+UoYA1YdmofNwCMxVzt5Yf7eBz/rP64XVhAj7Kdab+tOPZYgcoy5Vw2w3PXd7H
nmcVJqKvMUSnjQaRkU6phEuId8NGjnKInyqxNi8T+9eTuO01KLCF0E09KAZ0IY1+JtZOWR5xSH4z
Bp09ZpPcvtklYgrjWnRvoefypzovXXwhryoQ6G5u74WuBFB39KFF1A3V9lttaXO45gv/Uy3Nn3hV
M+y/8PwTp+YiTYOfoipDtBLUZQo5pFTcvlG/t+o/Kglmn5z39iHiwpqm5iSfSYoLNj3JyM4FIn6J
ApqWJwho9SA/S+nKc+ZtaxYyLHa0V1d+ebQ4l1dY+J/qGlB3QmxR3LjO+wYVf1WQLGjcAEGbnOPx
CjxrNRS+PX/oFrnNKtiiYeIJQJr7TBldHKKjTDoM4Wv5MzcfpUsAHDFNOMJsA1BKpkyBc7gSpCpC
05W6PEs/vj7a6E7fP7E0Ad3P8OtER5bxTlSLKjHSdHrCeMR/rEXeJ5Vk3e64ZOsI+tRDSPJQOx2a
14sSSql0CBwxEHH6RcBD9DNdiuQ8xUr8d4uBpaoOi96FgABv7elj9QVXHNup5D0D6H4FB1J0KyTb
4PPJ3qZpkl3F9XSaeuKdf8pBidCsAE4tAVEfk0gmtlxwr5A3mVWER7XAu9S47lXbmaCc2G7galDW
Ec1M6IJiip+H4LJVQdNXHizK2McR2OxNP0K+1Vg5s5HV/+IutTH9AQnkqb8onWEKw7VXYU9yc9ga
Bo+eIPoDL65V3rJkK13kDkfGMkYlK+scwH1vd5CCgOQME8tY4EhiuEq0MR+GrFdfX5SEriLAzEky
NK2xg6IVWuDPi5HOgxcUOQyUMYw+wTwkzzCwEstw9hORWKClmufO1RRvaO3pS4H8fFVrWIayZ/p0
ZsYffHe8gv8AW6T0Rj4K5H8t6FjyzAA2zuUGKBT1+OxFrQBBIqwnNkXZ185Lzhw62tjtAKhNg+TT
dy8a1ZQDrKzM1GNMb/+NKxebIa1qiZMm7As+w3xcn+r69/FcxDp/D7WBWy8w7cJBvMhG3jtLJK/j
tMgnQGhXerrQs7tNiKUb5lFc+CVkocELzH7ooN6mnDpZRilAYY/C29ccr+at675SdMIQsri0zeYV
GZHKFa72G5AO0Ws0Zc8IyAEEub/ZfcyktG0bBfIYMQC5idUSjPsOYya9Qkc9m5JyY28sbJp4ZGao
NxRi81EGhXXD6/8EV2pbsGkbLH5zsX2zwHeGpxNCAguBs+vsfk2zCl6s3mZ3kssfr2lPnknZaE//
z0FYOQEZCzpTdQNUcKyr/HRTaZeFKJv0Yw6r7vl9uWKsBHqui4LxJMDNx2udzDnu0wjTDLuShWF9
TipmP6RWJ6enAufwieFe4s9jBRZ2/ZJxwFKwTV769ZJHGBpl5FH5UFGpZ1j4JNL1324SJV7+V4gJ
WGiuiQNKu4jB6ARL6zItQf3H2pPURR8oMWjoomTW0yZHSf8y3qm1Fi9ihr1FlwCZ2JZmk7wypKGq
YASE/oCMdHAWFwf3+mguGJaPZAIn5bjPJs9+bP5Vdnl7lvS2nOAIqBEqubBtkJBPjddfop5okMbM
/dMf6QY5sGEBHsU0+0IB5+phix+/4YhsoXgMP+EkosykJ/lPI1OXrZSyq4tYFCMMCAnzKUE6V7Rm
fVQbd2Pjl+kBqWp0GF4yLS8Xg+CuI711+3H/jckpBWN88a2i1+XKQS30Wpl6Cg8oBh1TKr1dHiOZ
/kR+IdvFvDOKIv3/nI4GRUjP9jHp/4sVvSTXbLypSy6li6/KOlKrjWEiuxuuvuIDh0QMsJhA5ucy
lXcqsHGh4O6duvhy7YzJAKGZd8oZiZb71BcoVpqPfL9ZNENyBkCSZyErabDf14H3d5q8vmPJsDSF
1c9noW0R6kiCOObGluYo8IWfLy0n/dW+1SV+9ihpA5wYdL6ScZ28DdNniXXufarwiyFKVymZqBrV
KHwxYoTy6qMvZggyOb+TJwRMGz6rc5CKuw8iflB1pSza3uzv5uk0cEXmymoIeNy8W6EJSXgY2eza
ynGP8wosr4fFVZnw/0OzQLMPKEbMbF3h7hxjPv1WrbyypFLFnHEK3/SxGezhlcVdpbc0/vITBlcQ
vKuLTwNprvnTJ+fIZfAm7Vf3Fj72bKv6x1AV8CE/LTelhdX+Agq6h2uH+Sw4h0+dg8FjtafNOE4X
myWlFMS63lK/e4kr3rOjsPpnDD6Ea/KuYkkTNOHNGJjyQmMe6X/PNBZPRAeKhNpA/AKuc/MAJvK1
qapsKZvk+mfZKHkAKarNKFcW6wvlUFMm8i2Jb1tGbuUxT9FqbjGEDZ9O83eTIJshLOSJob/s05gU
ELf2/h5DTmeBBl9mKmN1ROkyo1UgWm7jGN6Z4PYQpOuS0FWIioXtDu1P4bQSioH8myOatQISOb2V
ypg4TzoV8F5ZgyiRIV5owz4plGyjacVdc0otzSIxneWadb3ZPnVKog702GIq0ZVUrT3wyUT67RPa
Ki4hanv/EXH/B9w1Ksj7bjYt6wWJb4PmpJGooYvuHANQGgRGg3p5BcoGlbLp2QMpTaplPBymopww
eyeq3FfNIIa9pqGibz+IXQfltM2wvdl0zi4P87N7AfQGn4l7mWTupaFiUe3mXfXi7nSBOJGn55SW
LAKKX5BfEpd0gGJkJXMLppVkkSJfDOlf+o8U4qXef1TFTkMIXue96nbznZbSjoWBKZe8dnQ6XxNN
2/H3FlXyWYLpR2AqKtFuGaCt6E8G3qFTFWr/JXEu08Hrzltk3VW8RwmufNp45G+5mlzX260YrKm/
X0j6p7E+eEKaJHJLtFrV3gM2nb8YU29S5rqkmXUWESrwC8BaRRn0HV7FvDV7gsoFHOl0zQaQgT9P
NaoEw4emJAulrE9WspyTzLQMhx+qwFHm3sorl6Arc9eD8rlPw8WCMN9QGaQKa6Gh/CAEIxyZlcNo
+LjvDmdN5MhHIUoC8GaBcq51qTaUQ1hp3QvclMhYFATr9+DnJjMt1TljoeMKZ80lTpnoFBXPnHhk
3F7HOqWjhJYVhKKCFL7IQ9Infyb0aiuJ6Ee0n38bfZ/4B1LfKn4U14i9W9AKhlkbRJ3fk7d0JpBH
bggRn+nFWGkuHa/eskm656xVvZs596RadtWKAOkUmnPXCpvPkNhP9g6511tBUqYCu6DEW+QQhKml
1zl0xZn+jp41RcIqFNFaklslEww2Hg+i4LexZSu6ymen7oyR7a1iVbPbAlaWxT50KXiL33CZNVsG
+Kli5tNjg7KmIE1m2ttoLpmT5WO1PzX0dJkxPMp42utOnCf3G2ywySqp+nfDJRPKIKEm5Y+qEOV3
2IvrjWD7XYYgNHGE/i4GQKyg9ZQh2lzzmEBFBe4ib/LWc4bnDpJv0u0AKXqqu10KApz0X1Tn0T7y
2P1eJiotD4qLCnVd45NlR+8f88rcOoCUIO8B4RT1TD0uv5oaAx35BHbd4qfrq1nEIoOvrsK1paZs
ZZmMJq7sWruufdanR95+tLg+6/qmeidHLMhdbz0uSKQpEjl04bfHG6y0bFODMXGIFxj4olO0cUqk
FM95Kk1ovfL2FRiKad41hRrrOnwXjcoGMzfomqsNv57YipyaFX6w5eWLHZGulza4co3TMeACnIBb
42fTFTuN64L6vI0Lb8aA9OAuIIg9cg1Y39R4HQTMg4kLxsXt2OH8x1TAO3Jkifz3d9Qffd/SceWj
4b76yowrWTsY8Nb6sAezxK4zX7XOFolCG+c9qwdoyTcGOQAMoPcQM5UaKadYFCIAvIwWcNNfgHGy
WxAXkRGFpWJ0UnPg/jMVpVDh/YOgCc/RmRNY3G0r5uqxpV2I0BsaiWw2DGhEnuIM1C6VuLwMIItW
6brMrqyv3us10dZ4mJ/p32O3zbfWn8e6iDnRtI/zAxfVryB75Rrj57LDd1MPifR2tX21hKYNPIxB
mfIZHqOiKzsIf/mb9hFh9tXQ/nAPZV7yxf9pdm4n81WJVDUAZo5jkloBnksZjEmE6hFPANphhiH3
EILhFe22VbMkK4cIF2XmWKnFoxEXN3C/t1EUIH8C7hV7vZPoAclb9Glm+7UmVoyjum8u9p5xvgUK
szb1pWWJavQv4IvbjM99vlmjMKrtay90QRKisVNrulUp3koL0FsjIrfQVT6rAA0mdTIs59mPy3hs
KIca5o39/eZ3sUNdm+XGxVr7Mtl7vOp94FV9uUrw68o4ou5bj8qaAARC9TOEGxKiKLJUAI9EiyCs
pQu4zIeUjMnLD7+CTzjVzyNeYOBDUDZWRewiEb+Nwp3+nU03fZ92C5KU8WPO+fd4w/Dp7O8KCrg/
zE4E38jNC09Lpmwdg5qOsXPNZl3qvzGvezP0rOUJs2oro5OHXHtF7QY3xNYeh3ex9Fj2esDmxlbK
TSUz5zvg6B40hOjkp4Nfo3kHV5toq7hzALvOoqXu6K8QPePxbEumyTOyfM3AdgVYunooX3Dploj8
zEDvInez7ZYSivy1EJNUVcZg74rwTb7PU//kmKLYECE0417j6yvI6mr2xKfwVMUgVgMJUBvVv4EY
aHXv1OYkoTDc8It8/i8cTl9HROV4hv1vcgJMNsDFRiWkKf2LeISpXVEEKxsUrVHYRlUkdpbaJK+h
G64sm4Z7HTPb6FsNRFknzu/3EBcncvbnBIdR3TyIQyavT5ZSa3HNJXjXbmrYzOUGe0n/+rFXlkk5
wqsw5xlYFlpIunXDV/JCXyG3s0t5QLVcs/vCcV0JoIFHhh657TECcRgqPe3O/xk2mm29FiPd/xDZ
kRgLrWOXTGYzDeLDk4LJzwVWgaCoL0ulnhHkzQD3ZeBWQDNoYVeTxpSiE29mC5EK5228InofY/XQ
gpBjZxsJrUv8FPtNuRCoGIE9AQDgQKEcfqWsiX2fPXka8wJQ6uHV3y8Q52JqdGYb9yPO+HXvYft6
4BNN4SizGy8SUljVCT69TXUc7JB+w79XKc3EoCXJwlti0EyMGRhKmIWPABqkeSTt4j9u5Fqe5ih1
b/jX6oLjsnAbT7XKFJEICsnw4DBpwOethb8eJhtj+C89jEdMfPfBXYaIwhk5DIxImnN6I4YYYN6N
Q1wrOnQFwBq5I3Cwk54p005jYfaJDcWzMrMayKUXeBvsK1UGsHRtTrmPeV7rhe8QYZ4Q8cBMgM+u
kQkwTRyvOG7wH3mCplKfWXDDKWu1DBSUiymzJLPt5uNtflhcnaS6v3KMBmNR6Ae5B+VKSxlBbDi9
MVS9Mg9KbNUhK+fnLFsYmXZ0znrY1XOPfucG20aoFpPf+ODeTbhTIs1MOXuvoEQO2meJpQHkAPjN
hB2TMlKOU8jX1khaz9H5VTgREw4zMe0GVm0e/z5Mxl6h64T/OoILZQrrAMzo8QFxS45i4/m04ZPZ
UqMVZANAXKuJLjdg2+W02pkkrPB6vt3NnYYb/2c3XfdVZidWIy3LbgtYowZ3qrn9dvPtC5Yqp8dX
M8wis7mgBXr3iSifeVJhjF1XpbfjSI6NMVW54dlbFMaoXFqO2ztQK11vTlAjRQAY2hPLWhzxmKec
UHOhrdjmL2fK8Cbm36c0Lad+J7DWFVOo8GRI+6lH08ol4aG2pqUkFQbdWaBvvRTghM+PlThqArxQ
1LqFEQP+a+SfnO3NtjRLijGHigzznPl7B4JYhkFRG4pcsJ8oh/KjkOznkZoFyOykV+i5fw6jCgNv
C2hgiJ1Xou5YxdwOE6yHhuC2PEu8zagxxB87POKN+RHBry+li2GtHRN6zTpGLLg2mTtTAy40Gkw4
g6su8U3BoaDaj0KhjCkYozU2fYeRNhuyIH8G2eNMKxRHAp/G4MXHK9Kt4WrnLiL1lD9wAPaLoF/m
/zHa5KphwZfAlmuT52Gp9LEiG74EWIwhSS2L+JrcAORrTnS15vD/gzL+AdEivtYoa0ZdxtQbiJoq
RNWQWla8pBrEYo15qmWAzxFd+POAlm5JpROqoLf7uLNiBi/8yU7RSfEWpR1EFJQT8UOG+A29ODKZ
fadSUOQVPtLW5YGS1CSBa7l5+DjJ6HReFM7Pbjqt2cEcMQBKwb5GduGmV+J3nTUryq7NAyfhxTVF
Uy2eecwrnvck8C3l35IMWgdoWuomo9RP5IV2z+oxeERFsAX4view7pWCsqCcxhvOlcCP5gzorKEP
Xu4/latqS6euRAwgNc/Gk9/gTv+8VhVGpYHmYVAiLNs4+lRuIZT6EYur3HxUKOBMmQ5lBm++OPj9
Xl23D76sDu22Z73HeJhsLe4qBXAhHhDElWdAeDOb1KpjWGT/Xg9fyrTrqlCPh/GXsety26xSPGM7
2ARRq9+8KqSFoZ+bgeKBgvZZy3SyPI9OhFP1oeG0ZnP5ORtncKqm/azsDWDNSoLAhV7CcVsV8Awa
X5aywmLApsTFPuud/mBHXWUP9y7E4yjdPcROWW6P7n6vWv4lpmScTBFDU/RNKlGSXJP72+vcP7od
RzUBid1hjliXXcX8m4ajgs5ICP0Hg5coWWa4gAEnm9pq+CcVwPnGaWttEXUgwoITL8fBeT2eWUyB
eIkwwbnWU9d5IvLlai0e9Cegl/jofoynmVx45qtnYhaS1nLX3nbQ7wosJ7gXIUQxqJauKA+Z2KS6
bicF1wz7Wt3tNEcwjM8bJiFVzCEEBiPWXbNm3Axgz9gbSIgXvCJ9fmaeHBtcPeIo98Dd/XTj4A/H
hCFTSAfWfH0CWUNRrcrgDgwUwkohb0U0SAMP8gAqs1TTgY+QCk5Pyu0Hy5fb4dOqisk5Z6dqqkeR
YL70uAEiDD2z0ObgCf6LsvS4y7hfZHmId0Dxp8qqXApnriZdvN1nZpcLPxwaF2HWC9Pw+JjAez1M
v80eDGUe755jegOSSVlZbT5Em1TfWClp+H0flYp7kplEFuM2y1GHkQWU2HgaHDsqUIGaJk0q8UrJ
vI1jPqMS2AymbPxd/En235cSYgpN4ezvkouJeNjbrlf5xcuJk25QWEWxzpmOrgmroIZpWeiXMGCC
CS1bagjD95fQVurLEjNzCwMPLtHptiPml6RCHH+Bkhi/AMrxRX7Z0IrTuuPCxY6g1lFo0vjSvsQB
OJceAhnEebK5wT/9AJmK6TV08aQ0AXiY7rJlv+4Dl2FAJCnPn2UIUsU9hIvCxlt35C/qGs8hO5Am
mKQIj6qH4ezfJfpqa5txACg+ovmzX9FogwaGjNOGoaaLoeyH7b1N+tClhzms7+WbeLrQYXX0OkS/
kP9tWaXVCpgWBAosNAHdk/y9i+R6oVSH1C20SAxqIZpIR2CqVDx6fAbJOI9kA4EQyZIXMAxB5e+k
UIAt6I4QwoDKWitbrpS33zjgZZqaAe7lrnU1TFAzwsbssGiChZFdgZhSBy7JSBhrac3qf/3ycrts
qcHJTmk7BBH+LUolgsvAzVkZrlMv2o6u70GxaZ2h77YJlbILIy1pVzPVlHu5iUDtuO0MYgH0tGHS
yyS2CIobjtqtWT77nppU3bHq0J+Gra/tPB30qSagn0ResohYe7ABK3XsvCzPEZA4m7k6vF3LynII
JKrtnlX+nrqmib66xtlWWVbRc9z0OrdhR1EVfUF5+Yn/LSStumJxRcqlT5F9jBH8ZkEmZ/aQpSFt
zTcrPHb5JpIbwutG2+dBwSWsb9ivGguDNwM+HuUBCF0YO2pQT9BnxYg1uPeIuzmIrUd84kjFIrlX
9s1+5MG+sNai/ma/maCrvNDktqCDd6sFfu6HObMUQbBk/0IaP4E/B4dXYuZ7Wo+EsgWveM2C0/nW
uh6EpXcmx6mttJlAwhHXTFerIkbn81DpzptLo6VbiQloD6Gc3R/TNB4EeSNCcyvI5PyPOzMKrTx0
DIZ1HRY1erM845YN4lVaSOX3mRqxUTeGN2+UDwzwu01gGFLg6H7s+KndU43uH37t7LVH9EPVE1N4
XnPNIxJ/SIJVzveE4W8Due3xznUUGK7umJyakysQtIImoz6vmMQ1SK4rAFsU85oUu80Xna+rNWm0
zOyJ8ECZx+fNKsWkaQsoq6uTW5VSPXONSW//1jAuDLCNhpSakhRM2mjZjozZQyb+by1MMVIMkB3o
Vd1izqwuREPMBrkQSxXcHzbdXSfRku7zrMx4XbrNpe3YL1PoDsU4pw4xFN7Wd/BA80s8hcZrIff6
AzDI16GZ05x0XU+WSTcaeRoboFniVitmdrSmUTlMSCD6nSOnpP8nBrlweKOUCz6S9n9G9iRCByJL
/b/hwcQXTrKsOgrxB33ahIg7tS7CYA0Eks4jpzoIK0Rv/aLQJGKd+bcCrJCUrrgH8Yl2yA7t/smg
Am1BoQZUfgF+wxaJsGzT987iN9l4FY2uAuEH28cX72M0wIDWXaFVBdkyf5RDfCUxW6uLoAedNBoK
In68FOt/N0B10u09aj8w9N9pxkfeV/Xb/JJmDnKGHMQcxZQSDZtGpteEcydq+RSnNqJLGJfaSZdw
LcQBVxPj3qUKNFHU3nbxbWhsjfAaUgmZVXYifRO06dc48qmzF8DbBegMVcEQQuy+3c/MToWOL0se
joMpPD95+wI3l2HKbztT609g1qjXagCVMlaQmk3vBv8kPejiknog7kTnGA8JxDdWDHnKMPplUcko
IqSKHNc85oUJtp9b1wFOX6MH3XOGyrFv6Hv+8cT4iulxy9SFcTyzA9Z6n0STJzZEmsqx3ftvoNgk
geeIjreAcPsa8CUjDsJefncPhFvCp2kipLYzH2BKdS2MVcsuKdQycc56Rq8uZh0ptZ+BTyWGG13x
ykxGZkq7sQKzcW3c+m8O/1TY+PDeXw7VwUCACaf2ssL4jQ+FvH5ojj3/tAbLJWKlABqWjR8zOE09
OT60cb6UOqK7AgEFd3iASgz7w8cl2brA7rhzJ1hc6QuWGxIGQEny7BW+E0+1qDJWZGslojkPzurA
V2+VXUK8O+veYZ/b2XSPolmY3rH11SKfl8Jh/xj/e/FExm4wYyuW4KQzmFDqTzDB/ax96CCQToOu
SgmwtMtdso7Rx69thni0YwYEjpRICcv2OlubMq8xz+FLDB9CFKkEUpYDi5VM41lgPQuxI+7/WtNT
ibf3TTTTVF5det/IyCMvPNki4CGy0MIKoOjEsnPruQI7uohvSLfUNAxGYGkuKIjdT3qQyixPXzsw
zEZ0qi7LQ1wu1BKwRKhgsbdoi82DnbxzjRBkW/pT26P4tiy/a8Co5HAsn10+UumVpGTYpv82AXaf
VHWWZLGBfRCnABJFeI4f1nFxJXlg11tXY6OTY0VSCcIwQwRVwxy15n1UUGIV75JUxn4CgwlX5Bea
9/o0huNHKtLidm5bbgCr4ePMa7Vft87e+8nmrjjL+tk7HKmwMfS78LGvXIU5g42i1M/hV1bao7T4
Rid3t/pfwZ3kpWdIkLguI1QeMSNqFF9MFeRE3iSRbnJxx34w2zoB1nETLDUbRy0/uKnuzg5Uam6J
yvubMjrhi8kP5U1NdTMtVRhYfD3qp4mI//ACgSJcTpBJGgSqNa/acMoEKF+o8fVRsom29M0KchLt
FbtASKIs4csOdfaO1bpb0C4EDAtN9pRIxiKA9it5uZcpK5NunOU7IjmURzc/xRWM3d78AK2HIznW
INRgpkHUw1pMX7tP9J5Liz8qTEtDZ82bbxt06NSjh+fAV42XjtJRmC3aphmxvN6GiF9a097NHA98
2QMiI6o6frCL1L0XGcU8mFTn72jHUPrE4lrunaCdZSDLDTFpnmlxCq3Q5x7dbM08/7iTtHp/e/zx
bIWJwSJaKbjRjPJ+VtOv/5DgDMA5+GHG5rgMMCm4wMgDOC6Uxx5OfHukPMopsFsjs4g1gHPmlqqS
gDvRhSglaWEbg7TgvFkiImyA6jQDYWV4jQlBkzvted6LeMHGtmVd8R38jbmY6ByEnszD5BGF5XQo
x1aWYCHdNBlbze6+PE1hHufWJZ+JnEa0CnOp3VP652wQ7fDRTvA+r+vDFhU/UKFRfIsQMhVWZ/it
H4EA101OJjYg075bOyDZPJfVJMljCpMl1rBt89z8mW7M5Zw1iMTlaHoI8tbXt7BzAZwxLmji3Tz0
Pz3bi9li5bVWx+DiQpdztk5P1d2lQK+/BNiv6+3HM3YNfWDSjZjXjVE0/Wtb8NbHcSBuMeecai8N
e72Y6v65X/UZCBjorLy57C6hblTP+ktunvo6ZbDEQ+64KFGh+3MRV7ABClKZK+83kHQQZw2yFB1t
aZUrZkjFM+imoS486I3oSfq5i7h94kbrLEo5RNrlx/IHK0ksOALd1/dXbvAT4ayt0sDU0R7DQeEt
BNOItTwy06RAh4p/OYnL7aJsw8PyXatA+CLfhvEmd+f6T/Jp99ae9v9X4oqq/xi5Bt2tKN8bZ2MA
rFk1cy1imho0Sbk86ZiuAQFIL7r1HXI/xyNXYNDRdYTAqFvtMS18YAKg7E47iDGcnFToI9Wq/kpt
AW4azUs4C64LmBB5M8IrJbrHQau8/fpcXLFpBqHWyNSy1k0OQeYWk6yOjCa8mZlfP6ylwvQXGYtB
vWopKSy3OYy7TNJQ3/ytT6DHF3/ATCxYVBmEORoRzrocIWUug8I3AxYnirrfc4EJ9y9iRbSApA85
Knf/XLAr9UeVFGBcMH0kLmDGDb5C1amnjMK4UPV9E1pINXjqjWwvrenWvey41tB9WbCj2owK69gM
/CaI4N4jLvsDTxE+yOfr4Kfo1zx3XRz2M1eg0KnR77Fm/Olc8gUwkFalvejKW2UKlv40e0tHZpNm
2y577vnEvFr5jCSABDbz63KvOioXuULDX+G7FzPJLorCwh9br0e6gvqnin3sdiCc2z0+JE6KabDy
m67YZtoouhd4ISdNk9J3wMVvwhftQTeZEtJKexTOEqZdja52FF4NLVPE/ZS7bSjeqS1Su2aF8umY
qEYcTYsNbGiJN4QJXdfpZkb3NId7xnFfRfrxrBaZQ1nxSUqSP/8F/4OY7c7Co2ADcFv6gSWUNw95
//68dzf3zzCnWGZ/QMq3nGwLXUy6GY5NqzP9hWbya46jFt81rG5Meyda3Ql0XmlvJsLD2WPXVmD3
wM6PhFfOM7L83QIYGzdWFKZTxh+fUXjq51l5Q7wl9IYWzhJv3weVhqCJbNU4Os3McvnOw30yxf6f
fE43tmjxG1NR/oobo0/yLKbYVQbPz73uVV/XVcMJCUplp20eJODmWpHSEsa8VT6wgM1y5y1l81DU
S13ZR5pYqQJsKoKyxyGUcFUD34WWuBO3pKlIzTDVIsW+ynRqGJ06lLy3d/bZ6RV+ND51Tc5DdKDL
w0LWI/ql+lNp8yRLgwIWcAvUwSkciukPvswyEOm0ByEkN2V5HgoNwIBPkbtSIXqEfh2EqyrobdVP
qnCpt/9526MTD71XAuwgpORGTACsjl9ZMDCQSxXMgFIqWILjo84mwEuiVy3Y1+r388z3lZXhZDYQ
uxdZmwE+suVOtMRP62Ye8BHCyXXQRSbJjCbVimtveELw+9rvX3XhG2K9RmkF/5SsvhuUtHKMC92s
ngXDbD+z9sfsLc0nF+0kio0iKX/lmN9Hwk13LV7xuCCAT2EQ/PquKP16EexeOvPzdrQ4TabmfBn0
3XiNy3Y7Pxf4YlXRaoVhGYRU9RrnQB86lCZEtnCn9W47+pqHx41MwABK7NVFlAfMabMo41LjH173
J+jjw1RsZH7ozd15i7jMEgfei2k0jmE0U+G7lU6PxAlauShdv5Was9LGQwsf7c96U7y1MJCJ63pA
pHD/A5dSnL4vU9SQnburiYPMhWBF0lOmNeJE3QhekrMZiOYnKiu09ng1Hs2qnWCDOvip+76pd3td
3lIoQPu0gcIafiS29rWJAtbvj4WJGbKBIv6cotXrjUJPFyBoRcPdnIilin1EIcSzkOc1VT9YQvca
CumS2tMaNnaAi/sSeHEQ2Fdh6h7OeW6niUS40pmyAgs8ooCrXFW1fe8THoLp1D6p0Dl8yJpVpDpl
qV6fg3QZFwTDWXxYK6lxOzEdLtrR+Xg/yhomq9UxpmTk1Cz5Ol0mDNpwk+i69o9y2upSAVuXJDhs
Pxs7CUkMC6Do2ntkSTYPYXpITuvTHAuazhD+ZxYegrLlPz8sxgh+UVPYfNVK9a/Zaw/T9igqGpEe
mhj8WB5MU/Xf3pBhTdX9asXm6fD8SVEoMLV0GDZP3jrEvgrzDH6Fp6HB3w7sZTzuHLKa3hwHqA8j
pIfurW92VTqj5bkc+WG2I9icQdet3APwd7ynwUmEDcrhmJHaSifLP5onItP7MtvI04wX9GOm7klv
IJHEOVE0eE/cbQ0AWVWvlFIPvvsYn4tcAXEcff1ruqclZu3sI9Ul9DRzFqJxa9ZUXZaJu8pF8g8C
no58BTi0e9jPFSRZ7+VinTdo2g0q5tsFIeFdZBv2XceQyeg5ZJmsl/5NKfHSsP8wB2mfjTRkcVFq
Idw9wBN3+3CUEa+yMBXr1nEMlVt970RbbshRV1kD4a2QRRHdg2Al1Q9FnI+zSLMUQDYTzkHUzjDa
zBebDasUcMWRiCQUBBaIvnRIk0asBtw9JXj9pKbamFKzr5WP6oGlU/dwfb+rfm4YfvGLEi/F28Ri
WL8BhJHQn+6t1IDfWA1XNOsx8SodgIuPd6KOSS1aa9KXBbs0zm2OBoabnJBfRjNiBIALxa0SSVG0
rzUZ/Fg1gw2e0ACX0NDjFOdqZU1JT9dr4K/p2mMAgyb6x3mOoqicLtGjvtHSnMxMBUuk0h0NYoXr
p3fKB3dM3Fh1QjLfsMF7Y/pTF6buTC2+EykZz4WAFgwigXLQqdVjrPJmo7BnB5XKsOr1GiA4YEeY
E+22Etk4bSMptEf4mUe8d6LoUZcD48pL8eZLjSG0GFLkaCEw787srx0a2ZggzHaRuJ3Z05AF5zW8
iPQ1b3y04PLYwNmyyf9ReNGA27/SUaIrLPDgPayrSvLrU7oYtETgka1BuGQxbA1w7rJHj1pbOvOY
cMvkKzIKeTz/7PVvnwvzeQEacihOFB2uHH0lvQ+yiYSe2P7KOH+Pgu9e/TpjB2vXtScPbcyd7NZU
EcYgt3KWKYKU6jR6u8t+8sFgPMMg7EHX7lHYx01ZMkXu1PxfIdPkyDZ3v55Yo09Mvj/IFZ/Edkr/
z169HgiV8KCrlbdQVDhC7j4p6v+CxKNLERrxS6YxqrRw6dupk3wn8J53OO/YBlcGm3vU7AQSouCT
BahWgcgUSFvYKO9dQphltEBcx52CE9bgCBRN2aviOiLxZhCY/li26luz/0evnjKxT1U/7xmyVta9
4BFhNIhKsYDUX8B8HsmRoqfrBIAGDNqr2YJXW65xg+3DGQ+VRqbf8dwjSU1iSwIxbrviszObgg+1
A+1QVpYz9CwoSpxGUV8vmjDyqTAoJjMxpVbScdO7QpnHA/AWhe+wu2CiJxOVBJSWpL7PipRMxPbo
XFKoU629vIc8XD/nFfY4E0eeYcKbAgpwdq3ZYA+9AFNLy5mSIt810gBbSfM/Ybxv9QWKdx+5UoGm
WHq3k04oZ7hYdAp2ms58u4Edc/nWHuCErlv36y+6RCvy1SyexpWO+uXq2yN9Lm7LDQBqkEGYUV/S
SJsaZBv2STRQktewyQdJgWVbP8bC/K0AjGhiVJUeYs+JNC2FBpeT+unt9b5YzQ74pZCOF406IiRr
ynL1bSY6jcLPw12uaRkVuciKMaqEVlVO0/ngmdnq6vk2f11zrXhFkL7tFRAe7GPopXNY7U3RaCt0
fR1re352KGxyo4t3iWgz6s+WAx5+qybpPMZ3bQeM18OKYz9TEAYbIUnYnVGzrVK7lzDzGujlkT5a
zsoN1rrfy3Nk9vpCZcd+DpfWPXQM4jfQWWUvoZT8sLszfSqm+7ZOG1zLr4GSy1ogBhwW+ehQ6a0l
9cmwhJBnoSF7iMihs+a4Lee0mUDIY0WOZeby85IlFln/SN4my+9Lt0ICftmbYkXPWcHRgr2fR/K9
5ZRwaoNyr2yUVXxjh/vuoy72d1gaZgybGKefAJd+/mW4JCYYpCbygjqK14RilWt1BNWzseFaHVXZ
9d1h8kIqyVxMZYOw3iAXpf4u8B7OOzAVJWtq9gsKJAhToAb20TgWno6FifyTeVsGj1mGgd4kHYB2
3p15w/Ng2h37wcEj08GJNyzaOUaavp0px6RfXvPJJp4wkwNYDxB0JXicrx6e4plxN+1YonE3eGsI
l9bVMxH/fgo7I19n3avmlYIeXzDbzOrJBeiydF6Y9Jwjs+wxpQBVmHaWWczpr6N7eIHb5qiFWrb8
ypaIEmXyOUEI8KFZqlKkmyoAMJ/XD+igO9JSLqYB+5dLWlC9HY0rPBUHeqnY13aY8NM+3nCU1CzC
pwzuugk8NJfa8wDgJv508qY/L6qWHbhVap8KG852yhxniaA6M/J3x7mvaLj8cs0OvBFuvCcEorMn
kZN4ioJ7RhQwEuuhNRgQbRm3tyDyl5/v75M1lFCeSJcubVtIQn8ISw8GTwjw5natKGZnmmwabmGu
iQBbVPNIedJP+XBoqB402iN5F4b90pBCaXv/jwjb++PtFlC51NHEgc/FOQHS/K1KDeQEYyfymJ0i
gMrgmZLE8aHxWopL4eMjxGF1WoCpsdKmIYUu8oTPa6LPmnbf7u12BKE6VknDjBgOd/CfJjjXrdlV
AXtqTCEVxlQK5JAW1BWgF9kePF7Re2Z5BpNCCa2jHCyJJxhQeSu9t+IMdnJnshlpMpofCwREocUm
vrmpI15zAmaarAK5GK55IXeuwdgBYLmpUjZmewibrtlu91qE+++hnPYVYDPrMFFHjz5KYznoSybi
vGt8egyfQJYhiKsxGJraRg3zhXvbEHPibXGBDOBUaWF+VUX1T+kbrqg9+bfLCeBO2Ks5HlyAMrBI
az43lTRYQnoRXS61iKO975e7figPF5YLNNU4S5I5D4zz/YEaTgCNueWiwRVf9I8nG90feyYMEMJl
mTyVFfmHVFFDEugemaa01vzDimal/jrEIcyxQ2XpxSAcr+EjS16mIvT5l7blbX9/6LLikm3e/WSe
xIXupatZUZCqrJe7xNeiKSUFgWXT77x1W1gmdc4b5DixspLlj/WwJtAGCSAQitR/kAOBQwFoWNZ/
NGFxuepRGu1Gb2tnvRXnrSmtdYm9F2RQc+vHJpZQlZExBLfbw684iJ+ISKXipDYUqnNUvLjaJtB3
rFcaO6iB6hBa3F1giNToz02DhIphxQa8cFxVLX3nxeAOhDQL0S8gNXTDIy4jiFFbPl/Q1eTnm8Lq
tVt71V1i1eo0xh653CUGe19um3eAFBUcu9vevmHYe1sGp3GPQexGGPtqlfeIckBnttdIhOkv0FsF
JPlNyZwnHzqWLTYnK0OqB1pEDQqgfBDWdh4XX5zmFZXAxq8nKByt7SdhOir2sjpaUVyWDVVBg2EA
kWOEM68NdbtsrJz5COvyGyrZs8ymvVGi6+KO1KaLvp6TN784HvILOnboMZQwTqU7OoUrwlDaqdWx
SkT+PqX7jLZD59QegMx3XyUiqj+/wGBxrw2tCC70S13lJ+qAvaF5cz5V4TJYxYF/vH1tKHerZhnk
HQugP4CdiZCt9kzd7BLUr+5+Ys8Op+bS5hU+x+2xWpVaUI6ieijOtVCoXPVHm7lveCDy7sE/mDSu
7Lw0JsL03BW2wKpbHEOn8L6eWfnZtscWGNTadH0WO/+Pqf7flFkusJLqNyXbnOOrTb4rGvVbpPgI
4ZsWRHyappIc9FJI//U6ZaPTgSmI17+XJ3xmBhm1m/skJWmJz8MHEacCy0MRibC0ZgLG4V5+bdV6
jQEIqtEM1rUT1fBRs5zj/t9HkLX2TWRQbB+S1qScGP5Xy/1iDXLzSMSWDlFYJkjIO96ImAuxP/CN
q80h5ufXun8XAXowhD8DueXddAsl9QMP7aSKx0kJL/TODlinXq4H0IkWXtRFGSqhjW5CwEOo32dJ
/+SZT6+Bi4mBZY2MAWo0haHz8XG6LDLcb3xMWbZzrEGszfZ7x6ejTT3fkHRD8KUGU9/bScEBX9WY
QWupvuPSwTxvAzRB0yHj0eLkTrLDnt3mekBSJeZAEkcm75cHKzl3mhC7b06zB7Ekt38Hn7BBDiu2
3x91vyHcpNc/trgJWm/+t56uM1mmC57SkEKLpA7AkiJkU+5i8TmUt5mSLLpE3bXRrYnBRgcsvLCu
5JqHWXzi8n06s39syKZvSo0wBtYrbk3UZ9BaRwIPRkBqBi0QOL+QRDwoKEUTOs+NRUZz8tm4Uyuj
KX/+rTvIYLlwb4ECjVGd8DoPlaPFuNePZdrk7udVSP9p07NmSB4dohowfOGV5QoMQZTrvB0fggZ8
LSQ/uru7F49IbmzEQXoiRDk6yFUF16dn6VimsSuGB95RfIzvf5HWF1GfhqaGP6RvWteP3kyLlmNj
vMs2k1RdR4ZFfJOwsIYdt9J1advOgXsUzo4UL66YjulWF28K4p/uqgMxi79pd1GdC6+KhvmLDyqY
fUJ0qujBNW2JgUMSvYhvrua5umDm2LlbtbQK9zUNXp5qT8MvF2VT4p/MAuGM2O9XJsJV5SbVU1Pt
Ab7uV91vKQJNfwvsznMB4nSTZ2GicNoG+l5ksJ+kAeimAqppdBKHnHB5Cj+NNO1ckdI1a/UBi0mS
kT4cEMOsQkNt+QH1x2KK7WOmvqxFRiQvjAqbhVcgRfIyumhoHRhwtFPlSmUkFpuFOFze6EOhCQdx
9amkij/K5HpuiO5xE5PyGnQxjA2xn9e4dzbS6odoBwZLE0u2Isqop2DkC6FncgYqbJ0gI95A9VBH
UN2slYk3iwl4tw+36dPbxa/Z2E0uoSlD9MyNRBAPwwBy/pxcki8x0JZ4ADKfcI0dWmLU0gaqf7oL
XzUhZfoZwm3f8hT30Zu9swSuYqk5vMB+wVPgDV4M/ZWm5a26yPSKdofruLekAX0JuCJkrR4hb59U
t29X6AIvCPTo7QpPnGhBNxawkeD7by3J0yykSSmd37u+KK+Y9aCBOzEh2pfDfpjBLBjDoKbPXJJu
E7NdxSNgURCUI+SGVvAswFTybJ7fXo8YC/RqkO6RzTv9SJEaeAsx9ZA0NOMln0XM8cKi3yzucrMJ
pg+K3mAzSf0iH0t/YvTSXEdlmOc7hFDkvcaYtgy5T1tGIgNFfUJpTuZL0ARU8payiG8aMZvFqkBY
XO10USDBAd01h/vDSpz4p7zih5ltmZxavqlB0gRz2DTZRaC55MsiuN5gELSi+qnC1h1SnxbdZ9IX
RqM47kC4XlZpjCLHyIQwYpln8uo2UKJfNWndAid59F4hGiMbC9vAGmmtX1fORnQVvzIiBIYuquZH
IRfpX61GYuW/ngO1FLcc7xcw5QpTmx9tnNzx2lKyIBa3MqsZqV681VioE7D8oEmEsEAwB6Advbwo
cfyqUps1G3wLCupfdajtSzgCcKwc6lyo7Vlul/wSyatfWRTa2+lU+7YU5sYBDRkOv6VHs2T9Dcdm
n36giNm+7Ll6J+kCehuf1F5pdaGyripRId6y4GD8q83hLultENoNBy1O/8+8xA5ukRbzETdaCV1o
CFLjjHNLz3pDp3GqfF9TQwX4Zeii+5/i5kV4sE7/3tKT7QFyeyrRzyA1+hkz4NXYf7jOH2WPy7bs
baMjMDnAj2YGFEvqqjgeJDJrmw5nY2o1OgAO9z05Be4oMfdEigt0nGF0/82RJS+pzln0hyw0P03X
iKM/nylwjvxmmM/WUNucMNwQr/3drBKiIpCEcnCXG2Sn3kmmDkUNYsACPew7sdPxmAF/rCKwcCDQ
EbH2HQ0O5hgHjvESmpdujGOyp6bG8uqdy3MUlOi6ejCTyfOrKLWY+dOlXUtduS65j2LfaYVWrsL1
iZCA57LpsSylpouL/mL5gJvRU1VuBu5DzSjNNIrJrfY6XThxPsl6HHy1tnR5boR63IeTGgpx5BWv
ncy4tq53/D1fLKNvjRAWrvmLeQiokjobaUlxLy/iSE5S8G4vKOapaTSuPWe6qskks7RL3b8qZr/5
vb2Fp8FhFR1YCDrb25NIFMB32Vak+Wv5pfxmfG4FPqWGZ3BzUa4LsW82Wh8fmLSEKj2tKYeqY9Rl
arxDzeW2xVOgHQioO1WXcNaiRA5fGcLweKn+T4hb9g1stGUX93+Q/KuY9AXH9UVHQYkBswuQwmik
Rx5Vk7s+6Icj5NFoz4/H+5oLffe3kK90C1gIJUCrFLJOsWBZlcHiAYYDI1aDiNDQGDR8suDCkMnW
6JmQQf9EqLoMbdA7uttsCtIgEB4U2ocvPfRHCTEmToMDp0y/dWRzoUeGOFxgmFev2UCTrwSkLEaS
CCYHMlYg6TV5x6auNFyb0edrh9PDPmj5oMMMxAAhzKIngiSmsm3p7sXqdpY3iPUKuLarSZpA77Gr
7JuPEuhCP0BtpLJWmhj3FLIjO4D2lYysWL+ArMAnJfh4Hiv6t3rHX3p9mHCDH2d8SUZA5eKq5TwY
wyHDOUiTNNbDQAxQx7ZzVcV5/5jA8eaSAAsjuWZGreOmOH0+ZF/Kb0gPN0c/+EYIrDTcXCRCY5lI
z7pvgELO7f/AquNo+6IBqFUpFHywz89M0UfqQ4WW0XdXG18W0EL/v4/O1qdb6yYIH1Tt2P8DSbo1
FVkkMCS5dLUZDL/IA21LLb6q70BZ0awR3MRKQZXLYsQQrzBKiiAgN/6ZN5Y3y5RP4y7csqUxFjno
OpX4SGXhvhMhMeEdWYm7hQ+GcV8oLU5vW3WMf/8WJdGgbMNSjdWe4/mJl/r/PCOJncCENVz7jLn/
918q8cl/B3SukotmYBYlgQHc1ls/IXNEBksrxwcWSe32CcAV+nWo6ZvRVl/IpYT7U6aXnFSzU+GK
RLBhmkSrp5uZOBVos8Mkio5/UKEK20T48YQhWHsQsWKzuD29wF6mRWZ00dRmqZsCVQ1DaTYO8V4P
VHvpZIpTgvyaUwRbyXf393KWpEAH8HwYhfBEzyO5/bhsZyPB3fJWzjhs5qA9JmGKY5TTYNrvciQg
XTlwdaNChv215byGyn9lqMWZ0Sdi61Y024+VAn0DFGN62BNG/m0xI6TSaczwVXtIPo7QIDoQ4FnP
hW1Asz7O/qWC4PwodEo0mVX95CS/MCJqBZ+mBv2tMgizrv7f/wpvb2n+1j3lFiL3uOm+o4yiuADj
2aeVyllSzCjCy/PMdLmXKYQDEfakVmf+kqGlbXb0kRkQ3jLffnj1sOwBn5tVVr+FjIqV64U/expX
xNRcZuwdvqUTRW8eY7865jT5Ny/mPmRlGD0vx3z/fsyVFOubSlYuBfzP0tN7ORhsY1QqN7rL585k
jY7wKfoSrapPjD+IvoGw7ooQCTUM4mxe9bTSctULugAKCjD0bQIjvYHytwuX1OFmNhsVOpQ7S8bK
OsluV64XQggcbR7Q7glquanBxJsqs54lZ8nq/tjQ3ZqTJjpiHGYDmZOahIMb/56N/wriMHEFhfC2
duQi6RjRol/wjvan5iXLLEWfL7NGrItp8JXMigHmc/Ig/H9DtD07gNoktCjcfaBn7H1qb870T0Jd
LycxnQAA4KRuBRif5+KZjJtee0ZegumwMrDJl84nj7lSdxqDb8D8QIBUMcksTVrdR7k9RsM3ISyP
RE9tE9dupWd5tb8b5bAJX9MXlYP+Maw1jQXlzDDfkoD1Z6PWItkeUznTfipfapBBunMMKTg9SDwC
vKdhmEZnMFndlV5CMHygkz3hpHRfT/e7j9wZdjdmRqJyQewGwKTYbN4yY4SEdZKijBkxOsr6Mb/S
n7Xa24OwmcWP8NzFykmBXfAjy8AXB/kR3dj+gznWEnNieCG0JR+tZRl+Z9wgPi0SaI6jR17QpDez
f8CqU6v6lukVWAWDph83gO2+FO10KHYQl1qKxvvSekqCkSuWueaOC+AqRmORMkor+0+xftvPa62r
z82AALWTRzmyNKUd+4lRkZcUmmRQJ1nDNAj7SmUXwmMs52d0py0UriD5bDrUPvH0T5Y4O6eTrtfb
MI0zTBlDfP1G0phRqa1RveoCoArOS7pXEmPX874o+IldNsYpOGwl28Xcm3WdJwWqsHNwpMoLfGuV
TbPRgs5XkI0WJRt76A3b3CDgTb+9gWQ35Pp9WflVr7OWoSuEwiFtspuvo51xG7qOp/xuKd+KaM2h
g6trxl6FwZB3wznfIDwkowu84PfsKnMr8Xvv7nGnjw0DQOBdOdSBZy3rs2Hp7MS5HrIYvD0FJfsE
t6R0tGsPdFUFYdcVdlMVrbQLoAvucn+ltF8aRuajWnFVvdly+623HSC9XfYIRLqrv+FjAbgfkem8
v0qp111hFD3tFscmjnN5kR2TFRg8MNT7lAOcDkMOGtjKFv2viYbNUwlVPZnOzEe5vRXaHyLp0dK1
YIf8Wf43cKYDePXdNlqHUsy7h1/nbGQchI4G/gSH3Z5ZISypkHRU1KtdfnbMpT3PvuTvzqmD38Ml
KjUXVuwSebNKSN0tqaw/B5ij8e2K3dUuAJA5+j35dK8pDH6mjpYFU1L8+jCiizG49/tzen3TzFxv
E27ZSOFMaDyDFfpwajc2rxm0tj2QBx2TUxMQSWlSWP8cRsagfUBEjthXpuaK6gc1eRCb8SVpKpDn
j1TEt0D6hmTOyhESp17b1HNCRujdoRlLnzaYM+ZeDf8EqingQkQX/sm9OBV+57gPQqeiTL69elIi
iJXVSNr3hCyYj20RxLY9Lan9QiWIgc5K+i7SvZdHBp3/+buoO6j5149qeyGJluF6Ti+LxTnHve5A
UE25Y4dY3SE26ieTjPQDqEYbfK9cB4qxGINU9v34aPLCTEKysfOYetfRvrXBK+BwIyA+PiQ9VE/U
Rqobkqk5ePcO8qe9RtjHibf0qOb6pUaSx24zuDU/Fcx1D9wT+NJn3xUPPewoi59x////k1feXntn
nRjnvCWEBtbR9ZTopnFaS28AzpdfAamU7ScIxdIyE5ZkPfMWhu0puw/53eclVOJkKOXHH1AMwtXY
Nn1MwS+pv9Tp6SZii+u9Jo5OPlmzMOgccl2XWhIIiMsnnkBwU5bksTjQHZnZlH3YboSzgJp0lAPI
4RU3TZfx4jL1XVOmCZ6AxyZaDYamU1FsUMdtikonoiLnF8QvmOD9J02xuWntjxpdu/7q2lxSgWuY
piRlfoyO1DP9W7WvbC31uWDwNe+sdrst07s0h4EiByKq5goMgYQ1aPLjLqqgk1nNseDauGWm63M9
xgya+XbUNY+ub8k0S0xRXNcsGjqk6cePEhuLlzjVuChBPplMTkkUii4XORLT4iW5QuZW6yIkt65N
S81GwQn88Sg7cG5uygKXMeTmsn6RIHnmVIbmti77WlmqsjzhoJGhob2GywBgrN3VDqQs2z7hTvk/
HLoRmONZB5frakB1+3w3SBvYnUvlb1vW02iNpVBQWYjN//JapwJqkQV0D85xzc0LjMZJb/XicrAK
vYijC86YQt1qJzTefkOw5uXFQH1BJUqqCq4E2uXfZy61/kSuBLzsLINuTvThOfmzKt2hWqDAfgfD
ZNb3fxTwb7Cd7EAaUwhSzygmXIXxzGVBeMjTkLAqkqf/I3fKWhSj8VVhHLcQH/9dY0IDaEjgnqlv
BVeMzjOKCdf1LA89ijPhv2K0e52XUbpKDOi0PNGYTWSnM5F7hmxA3lPM5JM8u59QA60fVLJCTEVo
/BmqsNiMD5JXWaLBZUxsBfV18HdTv2CBTFzstN2aEfyyl7M7HfniiFsH7V2tuYp38ZpZVWrTWT1l
fB2CO5u/GNXwpsy98wD/021FfcrTH/OXFvr0YgMv3+yJCh3tEZyglEoCuj63/bzvrF9t64LTOmKm
f0uuk1WeQjkkI3IRmismnVun6whuuiPahi3bvgWkBnt/2p0dn17eT7NwYTWXUqouisNo0nPRjpXU
aTLcmWoK5J+Cb/yW1znR8+Yra3iNxq7h34Ta6+hHP4ZfLYtZLAi7fKAYyxNQiyrT/PGUvYxkcgtG
KqkW2NOrZuU3+KhNF2E+pGDdcb/rUzPSrIhMRDVl70tvJ1tv5ntDQN5yqicSk0fZagLL3wgoMiOJ
1LE2YBn8WhEFW3VXFc0F1TuzjEVTAdMUacKHDx4MdOLJMEkRydkuj642z9N8ih4rSG3kuhYDCpeN
8oaRRod/tZ/6LGqxV5Xc3md7WjWPJWxp7d8T0g+NTD0EUj0KLZVoL3/WH62rd9TFMNqQtzEaV1xq
RX53rsCmCmWIjNLU+jTgo7OMakpNCki+5I4iItlB+ddyfQEup87awsURF9V7youRkPQwWhjhd/uq
t3LtDlvpros7dkwDAxYja9JISFeYCovMXKOAG1QsIv9TXRS7hwbuAVMILF5aZCjLOchLbsQ3GZlE
fh9zIoEJY8UKMYUh7CDlczf02dhfsX2/rKq298RI9BeoF8iiJzIYt86dqMlLI7D3XcS+ba208KH3
qb3igEVf03g5rIsa5+p9vth37ffM2NMCAQxbP/9EeaXcy8Ui6CZ3cIqn5bMesZJV903O+2XnOSJo
Q7csUdNf1XuTEJZFRxfnx94nlVoy/nTTD2sl6WeOvSYxCShM0sT0SD6M4+7cpge1dUbrXaqmc/Cl
PyO4XZeUtMumvapbE+XTohcGjtxKOY/rK9j5nmaYbuXITF1sN1csr0/sMPJh2jq3F5XkFMnfNHTu
yzPyBQFtBkGnmWITUZuS/olcWYmWpuNI8g67luKgMsNlwWeqR1WtQfyTp9fECEl0eVVGcGasCf/k
T7qhkc9DnGYi9pXgsqpvvoh0hz3ixd1qBDvzPv6cyRL/i3UEeet/2YgjeHzCM80N2Rv5Ca69VR74
LjGuCyJTTp8FYnIfKfukpMJwA/y78Fz53dwXSaEGfKI4yTtYsyxM5wXFpf2nuQ+u+h6SvaOJLPz3
GTDQ68+n/F1/+njlqL22YUXpAS/oysj4Ixul5NWJtPVnU6VuwhaUaxDGlWVPFLUbc0UeSDU/ibMK
O9ZcFH8hQCmoDmI0xNjLOcEyix58uv9pm/FJay80eNQuSi3pka3AFsJFQP1DP2PCBkWWbXWIdWYk
r4N/RYdH06qXS7N0l+onI2S4XmJbc2IXdvS43HZFjMJrmjCM6NKLwCQagmynuS2PoEq8WloUwQ5M
5Ip+4r4kWYKNkRvILQ/wCrfo1Ipy7BUN6v6KP7NciCey1z8WPc1ALeGeeJxhy+2pT7Ub+01w2o8I
oaVvj9BF/UGZY+5XAxjmXGviAia4pxAG69QVxB4yJMkImEe7RY+W+4n419M8l6b2c6v7FmNZV9OW
E7rCt7s6ht+8Mn2v5gvQvlaqgq1nrhC5wIyDZRbKt2The7uVzqnmGkHzVYN2Leq+VWa3Lx3LoFWM
taAyQIeD6Al2rl6bAaX92kHeAmUjBqMxyZrpFwulOS7waYVy1BxgCV2/SqvjS7WlJfANGLRdMuUw
nCS0OLUn98QhoQZvzPtaxvYYkDfjyv3tzDU2K+h/vjiTEBDrTFH40dEqcQ5+qOrgNJfU2WJBFzVc
IV4XczCFKvEHMH2WZQsyhUE0jVRQ/5MnhFrXWPetf1Fbt7GoWgXrtGYsq4N/A+tZ1AK+IQGGFSAM
k9ZzUmD+lldrjNzBbzFxeV6vCKxw+MqlhCaQFcFdX/Pmspp2BU/EMklvbkR5E0tMdpCygz5rv4K4
MBgxun4IXB17A05FSy3E5b7lox8Xiza/k1EUuDXWtdavuEz9Mwa43P9lQS+Yf4ptX6ClUlWYGTUD
LIAb99d834t8y55LPnrTaYxdhoyedBrplOdpZ91Ot8rTgAHb2f0kygM5Qfq2LrsRStnLEfgzKReJ
5hGxFwRNYqCXI9aaWrJmzbWIGP3MqE56+ki33d1aulk53CM1Vn5ce6+/f0xcyotCiTvr0/0NJxpm
myNT+pE64CE5mHZ83unzxsJ/4J4z8j7KGVBbKFEa49/uSpJebtsnEx/7LK29AojMN42boz6BRVjl
OmpMPpN48pbC9MT5p2Wu+h/6WN0hIn9eDPn02LfZ/z9JLf6AJXC9W8h2rvSfX5/6vNNUrXDVgm9o
e9n5eSVVLi6NvwpuJWOsa4WlTV8Ua72quHNfgyJOaFgatwNcPnDVlRgB5ISeJmH0Ibx/GbWGKOtu
1taCvbqzXO6Dz3t3hT9vH+khW6/edFLU0ViI1D1tonbE6FgME9VvxqNJgukJN+0yNCs5eP971orQ
Nb44gLPlnLgDxB9FTkurA7rM2loF5w35nQCzETd3kJ5nZPgOBkc7Lwuov+vFYkFGI9w9HhbvRC8L
50zwBE2BdQ2VBo2vMzwWUuRZs9Uf3oinvbpEoTE07DvnvIo6xflnQ2+0ekA3eah7einQsII7vUVw
n2IxW0pPQ58waZp/ONBgWg+n4bpRlehUWSw0NEWT/OnYpr+S8mVD60JyEpkrkBQpJknTQgP4iL3N
7Q8bfxLIJAFO1rVoEs6rL0IcrtjtHf4pp6yB89kMUfpMIYpT++hr5DlvsdmZGqO+BhNRybsmvIgl
sVtacbkVQi7E+7INSjccZNS+zc2XamCXYmTk6OCl7VzRgoW1oBawpW5FxQ0b2qVXoz39x2Fit4w5
lPVHfwxaxAhuCatnM9twDXWntMaOlF4e4ucrBqFyJiuqfXVCSkHINLIOdwfUG+xEmRZIF8COdVu8
yio32TK6tCQUi13jv+csiJrg9PA6yL2/rvTr0ucpcAF7pLk+IXlYgJSAu2I7rnJFQm+cE+lbptWr
M67kYKcyqQlXd1IYN+3EPs9CJSGsShJhjKJ4rmZq6bUb4X+rvi3HXCMfF0Qky62ydSYcfhuSQP8i
m9813iaShkP1mBy5SvCcTMrmxfTPy7yOqMICjw046dviXOH7BE961FCGHRfd9BrQ5pdnfM831tQZ
/SD9/PXxTVdYyEsB1lzjQoPhtiniKV0ib6gGAS7c4EPxCFYEqSMM2oUxxSeyPbI+7x5vB9pOCcXR
meWIz6czqd0fFGyF/mNsGLW6lZo4We3OfuBMQGFm9elQGEFKn73qHRKqn7xMgtFr7QnJ3SLduXNN
b3cYcAgNxp9XN3bD3SL7ybz0sAC77ssQYyxXwwa02Li5EyJesQp6Kspqd/DfeZglJdhzJ3AFbLPT
kQBDda1PLoSmtFmzfIEyExvAm7cYf+XfsGAjB2D8s752AwWuGVYBcJcXToyh3T4+fpvAVkxqLLMf
dU1E//9KAIn+gpGJKTdKzvtkMjzQx49NPkiSI8B9TIT/sXRuz2gEE6rFE5i6kCEFwFj90uKONCOk
Y/J9jua2d1ckJUmR77Gy8bIfdYAJBccsqHlrU+CTHFNVVhGNy9B0jyhESiKphkgHbnfMlaDWjqxD
r8Cb4/vUtTi9itU5E+ooYNOoiBN5Ub9zPUHsqEYjxZr8x2Aj5DDgx/ofDP0HrIyKBXWBTKQHVgqq
Tnn6Gj/C1AzBXRKx6B+hHA7dCSQ0xBw/licRVuka62RFboedPCrj3+FROicrAIl0b6vbdCQzPhV6
Yx3H0wdPLK9dnnOTkJ3Db26HinQyb/Z6n3PLuhS55tsVvtYT/Cpnoihl5zfe7ebkZoPVIhnFFXfk
gqcffMbQXNZdumZ2QxNg/d6P749Xo2sO7Rf5yn+zxWowYzvh3YVEZgEXlPBmJF51fze+BTqvyXKQ
oZZifso4yP6dhYeZEmjmyIfB6u7Lt4LG3PdJyksR4nNJmmLGrdd+pZKjd2Sjgoh0A9i/OxwoaY4c
mWLAItEyh1F0g899t/mP9Rt1+W43sfxJ9trlh+2/Pr4lhScUxkF/cQ8mq7BjIk/+u2kzC2Z+9G3v
MRHOpmLLgqi+JL3BmiQY/s2p0mtG8pAa+1wH36jQ8aY4p8hqlkNTzVoTfAGNzbCEyzl6NXzN1POp
zahzd+rjgbjwnjJRqNw9WN1Fu2zJGKUK4UviEwObtJyhSjVO7hGSMccPa1QjbU762l3a7pGH0x8Q
w0O5zOzHQE0qzN5O0EMYCUOqDYyLKOIH4mOrYDhFsSZUp2ilr2WDYLRE/hS9cgpxkbwzghWMU4/F
WoTuMN1vpkXNkf/QZpRjYW0705Uw2+UglekcGGat/vnfYTXCxOwZy8FgL52ZVQjqgh89x5evyhHQ
fgqgCZGppuVjJL5q3Y6vKvR08TkPrQisaxNfjhi6hO2+YIJTxqa08aOce+w6qe1lVivBogpDdvfV
QMFIbjqSf/vrIkIwrlD2kt5x1LoWCpeQ5r3gKRW2iM8eLwEW8kdjBTdUwScKH1GNLtAXV8Dybq9W
eenA1GyUvirbGD/8IS3ZBb208Dd7Jb3egqdS87LwN3ZW1V2tZ7nHBZJT1WgWf+mg8ynTWdiFG6Mx
d1+0PIdbmi+8HeEPmqdLtgUw1MWfa98tpwhLiwAZzGKW7eX/bB67Hix3zGJDgm9aAZJ4sY+5sn/e
pebcIhfz9Uen4wLM50FpnB5qh4CLOvF8TVFoLfl95RZ0iZi6E4AcSdTaFRN4nRZynStZCfFW3pGn
uQCCeH4ULId7tB9SErn5NK+nEftBWsvWaKOXIqWf5Zjqn1Fbjdhg22hMALZfBNPd+HZeWx2/2VJ6
W72ERI3zQWUYlasWSqA6+wofc52LdtPTFLJM9ZKOz09jTR1wkd/VJaIPcCZVh7kFO68nTNTHLzVa
btGgZdPvOaLulSDzX0RK+zs2zTxCrKQZI50/De037c++YirN6T/jyUobw1Rb1W6/0TELwZxOF1l4
VrO0vOEvK9Ep2B6T1gncfPZVF4vca2EW80kFfc4FLxqfBW5RMYu9NNq72MnZYsb3u5dvsQ0SjwNl
g+x4/k40GP7LirYfpsL/K9GOPOJBuiSYhmQN8cEEGMDcN3U9Neat2kjejPTDXbObwZ5UEc/YTgx1
GBfJbexfnJ2p93FpVP0qT9/7rxHUYVHRjmC1y5QYWoHai+bPhNS5g97ISWB7JDMTPHnD/6Yzcpz3
bI8Wkt+8EYEhOShDTkr9TUEDWhgVxoZ/VPq9x2xn6p0D1OsnXVGgLW47PdDFDNRjWtLhAkomvI7/
nQ/djbZwu0Z0q4lc58nkJeyTr/O3gNcX0XtI5Du9uB+M+7t7gVglfxuu76MYoBtVNam2TPtoLZmM
y0o1ruPulI7n9LFEiDX+LcchtNK2ePw19BTh6bQMMUPHlKqzC1QXeozkZi8M7BoSL9jblR6dtTSH
GcgUg6VqK5qR5/ChvYhmRK2vXe1IkommoVUTzCB2LS6YDOnwCrLqz7cEPTRWvlCYkfSMWgRhu3qT
DJc238xGI6F2QOEYC4ba6h3FBlSyIIkq3iKsmIFuWJMQuF9qriWT1IGyX3i+/DA3/AGRzmHN20UP
dbV6gbVLQdEmoNQbYmC9fJKJlxVsm7RnjGSyguH8DrAEQ7AXRVCJUVqy6k64sD599/aYQNSemClK
Wm4lPhsFusBKxm7ghs6ySZJjIprLSJKw9idPYHopsKMG/CPqXxLcH9X3jzbzzo1hqKvh2hRDjv1L
sbsKsz77wRRZIoilU2U/1mSgtDXz/0CJExUN1vUzTKY++BcctyV1xfVEyDAFiMH3hm/lliegKiCN
5by8gaH2hIebHV1bSc5r28YcGtkJOaciDCZMvE02dflgC2WqcUdrWJ3emZFIZ3uz7us22T1ZnCI4
2EHic/2jXx42R3TOesqatYhnMnakHIroPWRmdwReI2PEa967ftfy/18HVn1/VeM3+l952Yv5VfBE
hgI0tApCAVMvojkqpoKbGCxAYtwd1PEuFC2AFNQwYTPzZJtIf5HoPwvNMidMX5UblQyQVNSRAeWz
8lQc/Iv0SVAOMPo+jMipT0hyD7lEbeszQAiiJ9u79Bn5A35aBa0fwQ6QyaP/zqO7OXfWav1S17nN
txJcDG/KpLPfLwriEmPK0K25WNRdUXeGSzJFgUS05hiqEwWO4B/81XmdXJUFM9INhSdyElmwsOoC
dz4JnheWA4UDUJNX3uwFDFsfma3V/YGGCaJEt06wBIWXk9kJKXoDJq7XvNNLhhp+bRhP49wAHXTr
t1myV0ECLNTwsv/Isq/gwdKxRPauM7Dcgsp4Z/w1siMuzpeYWSIVnIw9L42L4mFd7me9GB+lz+75
2m2T3PxGYJ43bNHiOdUogVtBFk69zuelPJpP6ZS7UPi0iAfdL1lL99eCsrO/THKBx4zakNMiZExq
f/k29OoFH7BDO7ipVyV5tGT4T50tPvXORHm5ONkb5oAR6SLL1w5M6anHPafh2CGbFGqX1fOyOZg0
JTLGDWbEO3g3RFAbt8TtLLXZnAP+FKyKalErkbTHzrIswNyVwOxbDgg43XEYO2KDqxNJvmuvKsPM
i+aIQbMo0YajSmWumfN1ygZ0IIq3NEVQhI5Mbfc4lSgaJp9h9a8d1OEvicTsko0eb7vDqsVW1p1a
men9c10/HSZlQaa9mTi5Yyhni/coVtB11JKbQ4eeKwzxgvZ1G1cc2F/8BK3PkDlumWzN3F1gK89B
13aR2e6odZwHVKuT1AgnKJXnxfv1kjVil70mjYY3hVQnDlO0gsUGsndI20zL+IC1UcfJUbJuouhF
CdZgGugY7GpTWEkKIVgvoUHWu37IglCUKl/E4AcztPTB4c799CXrYME7ruYOe/ahsyoT1/SpMNmb
Fw++fS5SKDMrYgFdD/OxeQ9O1Rf3XLy44fPkteWgMvFHvGQ+spi2vbm8VK27NVAnmlv1Ue4REri6
MSwqq+nlSZThysmOKajl0Ykq9Qg1NRt5eJq/e4Ty0ZoygioMoj0rFbpplmd7KNLuekYgWgfcRGms
bkvyNbQ760rrux+MT9YNnPLKN0SeSqXHh6suMEnXW+BC2e5Ybcq/oJED8gkNsFFXoynEkNObQ0hR
fNhfYuNQO42Avcyk3V9zSqdrhI5V9FGHjj6TE7Q5x9be+K9Mtp8juzXg9QFVbnD3FBfIiyJwj9Ee
ih6Ces4eJZX6LgGrTde3UILrG1lmtFOLE4+QMcw4PHbFHCcXOass06w/Sb4vmVRLOVHB80+bR1nV
CxXTckngnOE5CmN6SpXRkT7Gnw3kv9o2pGM5qp8Yq6b0znD6vgi8iomHH6TUda7Apq8xSZ66F226
Sx1wj7rfQ927Rragry0hq9fv/dYAwfzmPikNhsB3Il4cA8GQ8w4zpsWpWF2PgI3GTpAH5wPjadzS
uPtwI5Gug2MdB+r12CgxaXZBh+TrBAtN3dav2UETRYcxJVfwSoNBkUeF2QH/tw5OtVBtqWjoL+1T
bkZn6vs7t6IwYyi+InnNMsizF8Papth5/KFHASiyW9yMoePmQVl11O5YGDFJjo5dSckrmOBAGC+k
bgshC85E8FhK2Njnu6hs15PR6W6twF/T9wnM7qL1D5/aOS5H3LOskbJi0djZ7N/MCee2+sk961Fl
et2bccxhUL4FHNBlA3K9ItgJ0G/ASB3S/+1vMVfH6XntGg1hGuUV7Z/IzVvPq1/VZ9K3J3ajZFne
l5fSREDwLMot9Zh2VwDuAybSm3Jd5nEJ+uQKJuzlkQr8bPoyj3ZWZBooYqjxk1l3vB3DkFA7EnTg
Nqp02bj+IUfWuJSOa4hYPC7eR9YFdx85eCPiK0/6b6P+LpBXSUygkLp2Nyv8PtrNXABMNGlMLh7j
Lw8f2Y8N3dgBnfbtVquLozAKuy11heURVizhKDD2pRox0fwewRC17Frm4jBChkf3SucgLcPHZZ/E
6WKgy/1DyRBESmQgRNhd7PZBF3WKWrdQxJg4JI3n26dOSJcuc5U+wjfuas4NJXCeTkF/UlvE6QkX
jZDuajxUVSHbgz1+C406sGLjXYQdRCz6S4mLjcDp4dFg52feVglDXUkwNPivF3VDnIG0QJDp8oM0
BLe6VJ1Q9fb+DZArxuvFeqXUqjh8TFTSXafH5llAhPiASndYsgsp7g4qUwUbRrqcm8DNiTFZM3OS
vD8zGxNA5wWB1I/h7TbWXIM6jg03zH6XvX/1egVFtT1Z5mkp1ij6SiX2civsTDwXYArkiZjrhu2R
o1TsiFaP60MtOWi/Ozvg4R1EjWiJtnC/l8pt1tc6i25CkwrmYSkwrIVSz9IyR/31GfyFWsNJT88C
xPind5aNRHA23fx9ORRtyC+QQexmuusChXBPr9uZo8TxuzHPySJQEgiu74kdGauxhbj6lGyU9uWc
2ffFamzQjZ7SYOlVRQYL7/huaspvWtgyvLNIrQh9aTRYUi3LkPyNeW1R1K/cXc7nndxRSao1LQ+3
yjAVUsmTxYicf63ATPW1DAsEJ0FWYBVplUF729LeA+tIt0nxBZh3aVQ3GfPllGLBK3G8ge3DwW9n
ZYJxPiXqd61HDnRjYhzS85Le3ViBwF04W11essmb5pEq0RFBlOGffvAsU3YXPVhSOVsMej+l/J3y
ew+k3CvhADo8Fj58+CnqsbD5mrSMvU4KrcZPgjtDc7idU0FhwfPX65PYsBBrC8WkM2A8JBFoh3ni
NhhX1fhSGj1lGiNj0Y2kY1DpPsuzkLBw9lEdhyYyNikEttIOnGY+HROkIlwqQuhNTehxEokn1F+7
vlVmsdF3Y7sjK/5elOuawkVC+gnKpKLPXX4mjtRrwzPiM4G2K+bZ453T4M2TMg9Fh75935XF1/Hv
RDfgXC8xm4vsg0/8kP5oRxuMVYvndg1cz9JdApMgrwAJYrgzqw47BIPOltk8KymoBIfymB7vPTqM
0IdoO3eb6/E4JDb6Fn55NsTJQhHRPBjIFETo1OksAW5HwYYQiuyISjX+uQz2nm2lxv0jp7rbIiD0
AcISf7No0POn4Zi8NGXJoxMs02oeLuzCxhY2DyDCiqa8BpJdU5KkzGk27d4l3cCxJYXA9lg+MLfh
L2DV1HxhtDNQapB2tv4rX2ja6Zsu8wNbFw2Oh/l1ZiIecWzhVeQCEA1muTzyE+rPjWAGhU7YZzGJ
7fD8gRJigeqKeAW0PJIPvHNjMZAaSnDXH5r+gg50v8H0b7Qy94ofqTzbPGCCyqKsHkGLw1A5/iK8
o4RKjZyQt9ejNpRdVn9REDZZxI7vp7V9pMEwvkEOm1jPSKCxWeJmfqHJ3lEwKJMgjKdVNoOyDxNF
i920ieCAAhQ7mkZ/Yy4S4F+L7Q0FpZI38PYP8TTwf+PFtiN+Gzw5r4nPhs4HVKXIu9y2kY2wknZQ
ehmx/L8Rr5Y35hYGG4nksOCmVJ0HBhq3l8p7X6TMkG6vbXbXM+FufTvxecFEA1N2WJJpOcfeIB0t
0xjQLON+sWvWylexJZ79ETejHzciVHuIl20M4FBRsZnfM1d42OKgsydBzP3udeJocjtXhoejj3wi
OCVKmPHIEciwPSWT/INebc4jKz1gkRy3kbh0RD5rGHtLpPsn0ZHoOMInASpZC9xiEYRIKX6QBSNR
exrbBgJ5QJIsHanMwUi4jNhxTxqCy/CIZsy5KI1YIWyT1+yyv8W7XtbI1qq7QfvnUOy9nSuCBJ5w
XpUXpuhX8biGdwFffUwyVWMnk3B9dOtKYICVudpcLrfFx24kFqIgxoDJrq4tqFmOMy8kQKttpvkz
3wtNKnKA1QJVKGut3HI7KOMcsQGgjYf3uuEdh861BFSmd2aX0Oucm3xg6p40jBG8SoScbRZjYJkB
eV+ypUSZALe9JdKbGCXgwkCJD3r5KTaXtOv2A+82wdsvhonwQQBIgx60XwvNQGE220crhpp8v7Hn
uzVbDsUKYnGS+I3BdQFe+S+4yGE51B1gZ6CasJYhC9kXeVIBi31Z0rBRsgRqfjDSALa0M4+lllJx
YCw2sWGhq+jk5GcofgtxrtJ2Go6pI5phYWpI8W1/3pBidVm7XSbt0f0vo50xav6xLEKagLWqb036
dkK+k8uNfNQx/cieaHK9Z3NmNrw5NC0fFvsf0Rj6vubYw3plflWizP543xqb8KxWm5BREtsxbNNo
ZbMB4+0lbu/eKD6XskqC41QwKugEMBc1Ep3EgN0zewrkkJ8/aOlUAVl9lTCRE9bFw/tuyCBpIk+m
z4hrI/vnAoXE+K3LZh4fhEPGDzThqt75xNBRhgovJNDVO06fB7X1jIl1ffwMERZBknTu0PBr5N5u
ZZyOVrG5jjicvdiDZ02/a8rdKrqDZocgM87TUhXh0WdS929pMZFq9G3MsUEtY7TQjzp97Jqbzq9Y
aw1x07Hyf/eHc3xtyOEt30689yBbC7oQ7/R/EUGH6SpLSJOLNq8FfMj1ftSVAG4XBkQhJewz1vFD
0RgQAufSp3nNyYywWeOQ0/u7EPD0f9U3b3b6BCq+10yT5wqYbgLPjRmTnqmgslN/8M7eNp5eJRSc
RRQgf3v4c/y/4Rx7UW0nXtw1xfZWyUtBZFLiEVLjHxA+lIGSXy6ZpKD4zDMF5b+nP6TRBJwZeeym
M5ivDZZXK5uf3UIwo3Dm5AExmXVejTdK1T/aLt+61xqllMkUqxjbV73qbrs+CITMpDBN69kqWUEy
GZBE87B7nk1Gca0EkRug9OaMxa4K7cnJSGBzIuRKXpm7xMKjx6D2J/L3GtW7TIseyIr6O+Edi0ed
7XNqWaoq14zbOrG89ntkECLW7dZGbB+XxWk5UQdhoIvAH3SCljWHoehiyWVI3puU/iVXvgthTvZq
X1VcgIlmtDbhUHhZhuWXGwSxug+YhoCZfnXWL59QlBRgepbmuBWz79Rh6pVU9o4YYppTtMR5zKDS
dGGG4s0IejkPzKf0wnCyRQCoUMNJNTzen0dGTyQV/jUM/x4YwsnT4IvVxy9gWqsebBQ1w/Ol7rlJ
99GCNA4VchyUzcUWnzVAnO1NJVLLKoGSPNBToNsds+dB6Jkvqa8tlGstjPzngrDHOVTWGV91NsVk
Ah7wB8tzqfBYsR8XS5kqVMQVtTmEPep6tyTi5+dAO9vhncSr2f5d9mDLKnlA6UtwHw1fAsRkpz4P
/DKCt0GkjK6w5nqn7gtzbmSCPfqw8zgGZB7BBkJ4XR8iXTKolsrnwvS6Vm8vIH/Z57M5x+sKsQf+
J7jzNE2NdAPCKXyFYxtR1iLutleFAmEFwfi0zIZ+z5V9Div3kWdI/B+nRqbExyT7yi8Hoq4vP8xP
vh6MLowgZPirmgwmYYNcDXa35LxG45RKVsuLxcVnSXZTAbOaBv2STYC54oGGB48aubsHIJyzTepD
Mj7ew5KpYj5DfED9vtzT8f9pcveV8OoDxTfrz/bp0KlJClRMPHXI4PmNNyGKXaN8MTh1Ibt/C8ua
KhWBvOU+Tx/7KVUPT73PBjSoLo04hYdojaNnPlwOYfe6x4CdEk8ypan927TRYWSpEtxRrGZqD0ws
RdFuQcs7mWbZihLb8f8Wgx9gWS0EHsEJpU4Ff/g6JHl4GouemK4RcjPyIGEZoIHa5HbXx0Gadgg7
22FjbdKLqPkFy4NRBhzFPidbpPeGoG2pzugk3XfX836MbueX3egNEoudxjWebWY1G0smX1uQx7Yi
3AApaXkww3OsdGUiFigcWi6oJlMrO+Pk7gpXa0oENUw5nNiZ+HGBAfgEke1JSG50YuOmSOrKNHvL
+hIkzOVYcv1hfud/od3rsmQbZ8HIx7vFInln1/o328k5G34d7IddZt5t90yi2MSX2LwV6yrjRSh2
BCUmV6ym9JH5pzO5J5YaNAfVf9gvh/omYO2gtrIcrK/xFFoqV448xkTdyr06ubHa39DAARFgiptN
l0XotWiJGIJ9Aaa5Devjecce7v+u1+zj1BB4YsEiACUaQiJFWlxyCCNM+Ai3UVgrpLkWeH0bSuZN
NK95Fg1zrcD3oa5Hnn3S+YnXwYcGQh9HSX9IsSWuFtC+ggVbSam4SGvygAFU2oPrXUZESx20I/nc
uplTiL+rrQcnYBSHAFtyHCnht1loybCP5yNgk9afIco2NFuSPP1HUxI+XWGeiqjHU3qMA9lEEL7R
iSRkVhi+R8je0VRobZz3Y4BuGjv9u/5bW1lJrBwxh17NhXdQu1ZNK8FC0VwYh9JgNfzL89Hsj4MZ
SxkBSl2RCq07fKbk38s/C7/luUGLmXVNS9xO/KO/XruPDAe28cPEsG6jbMWPGzzkm1KpaVtLXHxZ
PAKFVvwM8mBC4m3Ywu1As6bOJVHSQ5VJ94LpI4UhDKzOHdI2lpDtRAQAUtwlZKkc038M16DKCjbA
ea3fJD/mH9trjDE1Ht0fZM69cVAL93Ulu/QDM/4a7CzMjQAFRLcD9qx6+P1aXE0o9kNxQ+dAFbag
gEPtbEpMp9uy8yLQreFitvQoZbR5q8MFn4ioUZer+b9l16SiW/YGsMvdJAz0ByLS+QWd1fCApGtT
OhAMzCQkCIodWecBFcaO5Y66pbfojgxLHWKHCysxZkVTzxCDlyYcIfSCKDfCMLVEIN2w27Rxi6S9
kv1QZe9fzvazwW46N9yOMs/VSQaezzlVQ1PIAOKoL13+4NiIkbNj7PRiHujhaf1Mik1FgOc/EbHJ
BEFeUHR7NvpOgsJcotn0YwCEPm7xVUxMtUjI5KJXzqu28K+x9NKTMZIFFjVuJcX0w7w9n5fXnFrB
17SwFNz3Ip2xaM05EuVZC/vuIjSeB7gux1mm1MmxQsV28rF60+91xOmpjpm4LX9Ve1+5wBCf2lnB
aCI3MVo4Nf8ArZDuBiwaadlxFv7FrQg4Y+9Mk17+y79CoOnPzEjhj3MnJ52flsJ4xZ0zFuCMvklh
i1MERWYIOxOHHzXYQpLx07GQaOB9DVvbUPsHTt0ommeqUYKS7qU4tZfhS0hNRgAm8o8u2StHXJOO
u5U6MjdnwmfJvsFrPr40KM8vPbsrMu3p3wgJUTUCvteG/cPGVxNot404ehLl2kGyjyAO+IWvjsjQ
qnUFP4zwsu9r05gW+YX5A4yJCv2I+ENcpbgj6EITh2QsYhFUWSHP2kM9xPReMRJXmDtPcsJEamIo
kx1/4PFXHy0VNX3mCiT/WKreSZYu178C+jjNUGcVz/tkDJnvHGDD7HgKBK5+mIM3BpkY7m+zrIK2
3z82jJT+pLzbzNOmTbTdDKlXOX9ndBn52/pnOVvQ+db9DaBlH+XxNi3LZ7Jw84GVkeyORl5atRWE
AWk9nmXkKrYjP1PsJn29w0dMoqYOUCaD2rFO073T5WvFF4o0Pv7hBX5uYDI4Bx4X+dygBV7jYA58
I+8kXDLJJC0lfNhFVjifh2jb+Plw769j2WW3T1IrqYH7nj6XsWpLcPAXbu1e6QLObRwpDm6Z10mE
h38OF8yjF0pEw6KAIwEG99paIWdm4JwYd2EcCf4eCyKzMKvq3lNEeNcS6kbRmius1lMMbWIx2APB
xrDcxTP4BOukdYx2QJuSqiaMrgRdJYHdYfKLMCZn+ArZa1j/gGCamnCiAjHs8tpO6zNyA11y7nJN
VRlILbOy5/sU/H0MpuPtT4CjPZjTz9dRWpGLBLmsx4EQXsCYo+Dq4ROPJKG+CMETaGfs/HM2eL2m
5VjHmkqOWQC1rsRyighALSQDk0Oo8y9n5nLS3bmjarFyUqrGMuIjq6+g/72jTSiA/JLKgOvnNKME
WwNOrMpc4i+0ns3sIWUAbXP8V7Y+6EsTuFrdf1p52p/aVvWlPl0Pms+Z0yLaW7xGhzFEMdBPhW/Z
vhVY6JCXNPUOwe/Dv7loVDJnnR0KRnD0P/5nHMfQSi5anRO4CCSKR42UEh7Ld5au2c4ZLgPFE88t
WH3I/ArisOGV8ruI7bQtgowZ4CAVSTHy6M9KcxPvNIzlFYB81stEZHI9ies8UIY9LbN8dBx/EljA
svsNy8XZ1SZh0XWAkxkwI4Aj/P5jzqnfCprzUtAoopvr5eqQtHDYpQooKTNNGXjKkz06IUPAtrph
FyTZ6IksM+DYQEsE/8BQRug/us7mfGgGB8LIbXmCFMhb1yr4Zr+K8greUI1Hsl/6DZAyG3AOSiH4
dibsZjjP2qGz5BYIHiBK42P+eJr24fnNtphRcw5j6nWG0R7n8WNIMxejCofEhoY7KHyuBOrZ7hgu
ztAWzzKXANeSaz4GBVo6Ah3+FkcZnxta5052Vz7zY6bpeg68x9JbrH7BtoFxAca+AUv+LUYSze7k
KjQgjWFjWURaUbrxT8TStMKFogzbsC8luFCxOuzyIR6KJgm5pqOLXTj0Ygeme4Y6jxFykwIavwct
DyVgGOC6UUagabkL37Is8UYvjqAGPAX+N3UUN3yopzfGfC1cTymMUELiFYd8gBTwpi6adwfV1gxe
kU95QVh3Jtlw1TdS55OZizJ9w7yk+kNsVFHlwZi5cAcsMaXadp5Mswt5FkDdilhqRvK8m2w3CEeP
e0YQJUz8pe+uMAklFJtk+ZbWUr9KgUJPzOconjN04K0tt6E4P7ZwHhylXNDNp4gjKbOe59xlDIY0
hzNg1YL+OwDcofDT2S1thhNeq3G1eke/j81eEg6nRj0rnQU6ObJo3wnHAA28S3lrTc3ASy+zzYzp
awB2TCWSFuTVrTby1Jc4cgVgAAQe6CBouYFeuv0WvBeD7pU/P8QtEO7IIc622UUyVZWXVLUmOjyT
h4eRd8tMObL5PuvNvrTjYovk9RziX+BA0umXISWGrqrtaji9RDwbpQ0HN9BJ6tCXtAPUbb0xU03Q
ynxos2UEruqbAISr+EmuQTobMv1HD7ve29enm4TByBr0thimkDCGxkPcYpuhw8KCZR9HKXxUKAar
lsfYneT9L5orOpVotoncXK9062mciDGYDSgRlgtTtv4vBNYvJeLMgS3pF5RvdT3+3hERNg+Xcrcy
F2fzbrQAPoyBwtBOzBfMxVtSb+vBRRr+5BfOdZg3Png1SUA2DL5rQpRYVTL35KmLOeHnmMzbA8p+
ZADGxbS9JOqHh3AMLCDCCin3fX2fUabhbErt0rVAGpBmvf8NgBuOsetyZMqLtnLfi3plnqSPEium
fFjOe9nDwtbX9lTTOjXK5Ciij6bCe2iQsIxeExr+PMhi2sGIwWjkJ83Obq8ZKA3IZA+gb1+Mar3L
yU86uXBPyVnXF695l1b/wIZA+kQqtfIbjq9d2nqTnwyMYSO2rEyaRJvvvt0e0OVYf7XklRvrIOAn
py/M3ytNquFAwVaUZEni9zcVu0QD4Dd81N6CBHhQCXxYLssyVuaN36IhJql73RL3LRa+Byk58Ux5
iR8dx3iEOFKcS0Dn7wU2/LDeaBilpZksXeCTSVD/Vdwh07o1IQ1KZMEN6y7rnYBaIVNUHs5nbAZz
21Cb0p/vCOy0DPjXc8KSymjzeqJuJwk5BI8aN+KHdFNmsCSPr8S1rXGA8JoWVqCCIMhIbhzlV0MX
1oXUcAMB5UOgJKtndAVAct+hxeH7B7l0zqEtlpqrutodD/yvBBvd5OSvk5PLpQtG6nR5nSGRWw++
bYdVYO6bRvg/CRF65h6IBu33JBIRqednhfgOlHcaa3gLvG2Z749Lzc1E8oLgSChLdzlBoakBktmB
YXu0ut5lfS4sTgQyWVa2kkGNgehmU6ytfYqtsCXg88RYor7So7sgdsGhvtkGFg4rwhdH+oqKdu2y
K/2Fp7aajEN8cytEioFNRCURUoIwHdPGZ3Y3a1TTaBST8Q1W4ZRVNzPoa88g0wvGuGl/aFVB6nyA
v3RqJrfbwkZVytWJdFLTk5qvoRXYy0mgDJK4rAj90kB71ctBT0fHLeJNVxaCkm7lRAz/zxHXkAtD
muCgjILpAPccUCgD1iwvBCGTrggUkHCCLS+1p1hVzWqvwg1fBi+ZBbGO06fz2w7XFvXBcXcUPSoI
+cHpb7wDPnjgL9XbtCxSsKKWCnaNYyXVb4Ig5izzH1bVV4RYhJ6AEKwLyGQUuTwHvGhxtgzGg4kA
swdoG4SK0YTPTlTwB/LPTb8xDQOBoAlla/vymMgVaPxSZn5jtUFn6IF2kMaG1PQnRYO/9embLl3C
LF5Yf2PDewNGKBO+HmMa19hz1maPQahThPbnF6LHAbKEzvN7EoN1rI+dO11cZSBWRXCG9c/yiQPI
M3sENdcIkdYTDKEpGUZc3tB6ThAtZLfVuKtVQEWRfVMAnq8ipLQlVahg6HtsvAAARrxytkwpAoQ1
oJ8T1yX64msU21r1aNQ253Pj37ohc/h94483L6/YingV2e4xrVu04Zj9c9zP1Eu0MjUyYX1BCtxf
Ck2YaZCr0NJmxMUF66mcARqGG0y4qpAjzilRo5svGUwsRj9sgYSv6Aohx9qV/yLBB45T+KK8lABn
dgqc8wAjgwBj9grxX2DRrz9xptX82NE07YUO7/gtFu5Wcx/K7nFIxOht32AhWkoF7vjyXz+UnGTM
MYKhS6Bp99k5fsTSJh9ga4LMmPk1leShXNlOrLRJpgdNyWTqfmJEpWidDS2QXafQiNLr7jUcKuDh
mKcwUYvkOsN0FPq+I3SS8+AtOOX6FEqzjQWR0NtfdBoH8d1nO39jSuFRz13fWREKo1oJ6KALAl8q
G0AYOh1njR0VM6xswHGZwixWPWpLpkNfm4U6A1cCapX9srhAu8QHwKPTUfClW52m83jF39DMs9e6
e8qPTm6z3y90VjEiBq+hyMK6h09ktF3f5NKR8z3Jn+aY9etUQAkt696ePOvzCnHGGep7zVkuc8LD
YGpxWnL/lrTxkcc6uAj8VkoqrJsqw+3CO3vkyKmIZa+4UVOV/RdErMWYzrzvCnhcj0x7or9foBE/
zBuQWlAnrhTlU+Gq/bXdqW2VRnHK6IkaBDNndMXCB3ENHL14owLONFX2HuZ3XVVk0TUlVz/TXV9u
vb+Xoa1CNcNYZDY0YHaX+bUM6MJ4DlRYS2FenvfUdF6IVUr4lOIJRmgcsR2EZigGlaac0scBBf86
O+XSVuIBl2GPxzMHT4Oa++EjfrmbYtv8/X9vES7Cc4isLnzjFy/YUXq4GcaLrXy+3bAZ3QKGoIO6
gatEIqYODRMnYQbVjAaG2xTlEMDo6zmIoe8dJdUY4qX6pdH+kmm6jMrsOZjyoYpT4JJ6HGpsoyJa
t3u5UaI+iUe/gPsK9+f/6TzOpVwLpesvu9bYTIbPPkr85l+/skV2yruX7z2HUHPYefODNgUaCaJP
/fNbKQZ/hRuogBpvyS38UPvw7JPf5rzz5emlvwQ++FJhHQlQPYZ3PYS7PyrDyNntnpe8gIqtVvYl
10TY747FluPo9Xdr1icmTTJFSdmTASOD86X8xo8Uod33+SPpSrgzy0lfV5U8LPZSylTfkMNC8/KT
EaPf2TD4nb79TNYjWCCc34iFYyFmQW85GcvD5D9bk78WfAnRV4suD9exMYS5hiNn/EPfZLzNBRnZ
UEyo+7CIEd87YgTFs4Wu8Ug5MW98GMt9b3YcsZxT1lJA/xQzcjj9/ssZ6QE1BucQftTRFzODpsuq
1EsjXFctoSs8fQyMxt3GGDyNShQDwEQFwzA/j5da7w6c611SvSbi7dIVBK+2dEWRQGcsFnxBf4Sd
2WXq1AdnTpz2aW9J3eN5YULtHsZ1bHdbqsaL8lF8xGJTobFs6R8+87TDo1nuIWY/Oe1Tr9OCUS0T
DowlDTK8fJrKpvm0neFhM1vLselO1UQp3tP0EQN88zXAxM6A6NKfsRZsqrZLnRpyFLQ+6MYsF+/R
jY4DqO/ZNqef7R8FkNtgz4SHZIdGRUQq2cL58BMj2dACpbNxgh73CMz23e5Q9S1M3+45w7Q3F8So
Yo03F0Ev5StIP129tr/1Jn4n1Li6BOs/qYa7ZdXwQEY42yUFsxYb9fzUJEVCdoCGEz5wCeq/KD9W
qOHAbZo5qL/hin6EBUY3NFXSDrBMYEvHreLLbSCZEvYw6x5bAkOZJ/wpE2Jy7hwZpgEbzPGvUn+x
/fihp6SiXXf7DXx2H9EuloSFkgWJACX1VGNUbaiiu+Z9O5KfsIlNZPVve1RQyr68INmm6zeP5OfW
mbq+ZFYCe5FIXYjcB+91WZ5Uiqs2dUj7UmQlnPxZPKcAmASJxB3IkocoF38hfsIga033m1Gvb7Ij
0lbdeL+6yPPNSbfk13mr2KNJDTQ78VanKltXqvuQTyHtW6E7xziiap5+gi42s/t/VGnLCBgRo1h7
m5ouJSA90r39EA4tCdhhUSho78WWJPlCiqJs5Dvx5PAuop7cV3x7B0wo9PWcOdWxeWt3HJD3Ia5f
qdrqiR7YBTq4wbhJ8s2qzm0vMvStszIKR0TSFre/u/+VjBX4TqxpRI1kTUIRXkjaoW0SssxBqPSi
P5SuDgpE3NyL5fTz841R5q7HHts1dG4j1p5zET2tBfdahLh7Kt0TjVwZP9ycjZ2aRums6AQ6zJDJ
AvZ7lqGiq3w73kg1Y+6lA9ERTAu+rzjvxqroR7FHRGH7KZFeq8yAwUfhmCR3sEueYy//Y3vtHAEh
2yUqEAZsrrZjJQGSecVehQJaHH8KNL2B4xI/S/tBo3MuDWgZu+UxZ8A8kDUqsW0k/PxojxXsDp5h
TPadjrMNOCR/VXK+6el33jbU4chZiAXQmYcNK6qZqNAXnCtSa79zFos35ApIuyejd6UEfjmK4Zg4
LkF4TODyIEOe4eW4YmDGXDtdWAMCqlJAzIfP4es7cHsp3vnhiPLc2U73ZYWGoT37pWOFwguCJDLW
C5mcCDJmVEXQsJe37CxQ8VfsHvZt3gSRjpMl8AoBNPlFQDj+eBN5T9KHohsNrwXV/RVaVdjm0//f
WdZqqfWv0RchSyHkdvPEPpKy1IQT6MkjnbS45zEmrKh91Uwf6ai7b6K6hpXck9bbcIXxYBH3IiNc
3IxDkPYr0699+wfsZA1afxBFoxTLpk+etMdg4A89+ma6/w1oaVWcR8Wo1yefqC6zHEk4x0t/VYr2
SnZu0HRRYfKCgYeb0neEe6sTJoYZdsNFKnxszcgI/I5TOxUOBk2aveq0ld4fHq0LZT2kBoNqixIN
HUxpaQPWNzcthEtniMgxcxyrW4pFIIPGe1260gEqdbxtrC8Z0IL6oWsman1LtiZAosaKKM3IGJ+J
IAils1wyW8Adt2K3xl3GO2nEqhVI11ly1hdQTjyHTH8iIt7HVz5EE+iP0/6FAdE/hGlRu1ECM31v
jza+sTKndYXJ1wmKsm5cZe88ieEEFiBy5m9+kYJ1wU1P1aU4mPuDqC8h17YVxmmMTdgTzreFRC3A
4yQoehr/NaPy3duQAXniO2vUtiJUY/I37K/NSAcDr4BTYIJag2qSDexCyPFJmTB7OArWa6RlvFCi
EeJHiuI1xeqyRnBeGP88A/5VnyuDD3okMCFS2JT8CJC+BaixPQgTxmPIECYJClt31ojMCPSlApG7
oP1fTGyIcyfhUE1JxT0vpMcSY3W1E0vl3hRiasBOBwRaBB+pGAsEEB5otTLpV64nD0n+LHbSuzG0
L+hENgoMuGcZIdeIeriOtCXyxb6DtK+vKHKGxteN6F8FyYMeUEWu8NbaZXoR9RGJs+na4Rmvx1EE
pJVvJhf2ibKkiyUwUUokQFjVGXZ04HnzTDO2rx26DIInEPG/8gYOF5Pvgnp2125DEe8yy3tW8xGR
tgd3yb33YrSYmUG6gv059UU+Amv4eML/bZgm6CbmS4F6GFFSsFhiikUF1G4MLAfRlStn+hFQHF/I
Xy0W4zHRzP462ZquidJzpAPIxSduuCvBblRv3OYq8LuSgbA0RsB/JGrC4iJLo1Fx4LfI0g32hzXC
INIu4Zvx0PzJlcnWev3t4p01RhqFjiIE7lN7pc1/2jp3WIDBFc4hHt1KAWyASZu4WqhLshOoOF+L
h8Anf+wGrnhfDZZGHyENcsfsBCBpbVhE8LL1Ts7pcxBsPDmrBw7GtaVCS3KXX9iJnRFj0xD6ui2z
/djAReoiWg/xSEPKRqdP/mHjDdut5ag/hLBjOMJ/1XbuzCR4WF6yvi8sdAojg5HVpPxdZaaeZVBX
HCh1Ze1slrTiL+0mebwbRfyKSPA++c/eY8IGjSjCXa7iWdxiNH+GIAinkFYGkoVprLxFBGZQ0YVb
GaJy//YfxJN+pxjF0aWB20Tyl35HGpDymQTEJqaV9PQaOfTdSJqGr9Bu4X0ImoONiFhkfyO7z7yR
b4y/Y3mkiWsOh2ILhKuntEdeSka+n3N08OEZVRVdhVw9Jlz9+OsJF8xQOOEG1AvQusfJ6JXzZQ6d
hYgae/gDHQe2jByYIj+1oEnuAvIHyfzHdQCFEvfioOtIZJW1vOe/32qUCYLzvbr77nukENoKXSuF
DWExAUm7Y+qw0+nFQsaWO9a9fIYCbi3BoQsSbnnmNHOeo0UO25o97Op2Qsq5+sbXS202DBn2mIM4
q8TSnTQ56JnyQduOMe/b0ZnPgnGZJhhQZQ1jCBp9b1FgqUmJvsWUBEs634zwfFWShqs8lXbCF3YT
6rTmZ95TS9rWZghLVx2ERExoO01aqsovV/b/qhejpMaVG8vZ0+B5x9UWVuppwzXvNRrlrrxX+/N/
VISEmB3Ql8PBxRkz7kpkXiRhymlCanJ55vX04/sAMYun2ehCJov5AFAqP4dIenyyjgo01a/Mfa9F
WfBA1sJ/tRnhC5hKmlhMzuMUiRtx+96AU87Rb33es0wZ0CYuzdHdeZSghjl/JWQswtxOFu6L8gxZ
ZdB19Ps2wuUnwAahDbzuSqEGrbWnK/VlG6yKjt9dZ1+YQg0DipYNHH6Z2kGk17xMiC5qay1opnf8
SAxXpbSj51KCkyHJL7irAqfa+na4koiWsl/oxbvXPDpDqqy6Z7o5wxDCppk1VAEkGPESLrCoiXIB
WG/2MipaVfWIP9CTHNvONXJjcfgwz7Amp7RweeLGr8V06yF/IZS8XavdVCHzqxXSaXUikBr9x9Hj
9nGgKu71C8W7ozoV5+ZdBACD71pJGunR+JZI+F84eKE1azQjV/CcLePKclGMaabv4ZDqwvsQ/dwO
cKDnOsihY2A/BOpPL76r88zdGjDAySkLZwaORfWPQLSO33c/mG7wKUMTVvbb85Hkuq1poM1ClUFA
jZeIP8xixingvXst7q9sx3de0xk4MP/MIrx71ptHaLYf71KQeygdPpw0abIk/e/trd4DdkuUZW4u
ieGy1iaMA7XHxZe/VSRlpp4KZNU+cqu1h3cQu9UvOMWo7j1nem5Tz1MY3lyiMRoYIJFAj2NclwfM
HOS7ObhdBwO6XR7taVPnsZqSyu/w7ogTOhumY6UR9865xhJMqdTWJtbcyOQdh8l7KU4y2m+x3Pzm
8MrDLJiVLYBUSideHVrOVb6UzpdGhIoBBr7WbytecoZjepP8UTaj6dfgu/gX0Uksq7OGkl/lG0Y/
jF7I0S0mFteX3UFX1UwbzZ44Q4Yl55tiwSadPaCk03ESQ4LbQDHwglOsaNUPwJcSK8Y8xA92ih1M
OMMmrtsDr1f8UF0FeGbz/VHxtZWLW1upAj4nwIstRBYfJCFLMyvAnFvE3R76DTlqauE6VX9O1SmF
BIvcsHevJPrucFwTrtWhv39whDyMwFayKiJZ6/OLggv7joi9z81plCirJTm5rnVmas8h9eV4rJq+
2KHYADuii8rARvfGznxhce9E5WrEKH+diSI6JqiJlJtB1rB2+Pt8Z0oGxyDM6XKgh7eQUGpCq3Gv
xn0l1jMpNsH6Ua6Tslj0ZCa05e/XA6cqQZ9U++3G5VJA6JvVScNQs+jAawNlRfEx3ZaEfjnsdvuN
ITNrZcEJppNOMmYJwrSDL6gdQBvGi57sxBLSiPVAhE/YhrVAqBZXWXr1GcUCprDcarLVXy9f38Cf
H94DOtUrbX1b0QxltAU//Ytt4qgxgyO3fFxEb2GFI9CmPGq6rYPQQJUgm7ZUuJB7nC9qGZNHr+ds
a3zbqVkDlnBmk/CB38Gthl/QThiGPx0WcSS91TBG5AU+3UnLTWjYKSI1ovVqqSvUyKeM6/sXrCBJ
xv3+VeBP6w10+0V1fTnHVm+c7bhAcIkjw4ouHNIlToSl1VRqNojuIiqDsN8I9JUuTdb+udh8Plqw
QYyzU8TIs6bZJHK+L2IIrU1pnsCswFLtz0zX0cnoNHTmKq1lm741dM3OZwuKityLMEyfrdumHk6j
yEnoxzqJ4gYVX+uz0MEOOvoXqC8ybjwee0hhUm2gzUmI2QXPV7vaNiH14uHxpFdak5vxje/RhLSd
dogTnlDtzz8TMuSHzmdOt0PqvIyp+JrccXFd31eIK5jAVeWSV1jgFQYA8PAt+mQdLFCiq2HMebMX
n2/tb97e9OlQVsSVso3j10omHm9B04ruWWWvcu9bVKyEW7vBeEdwJemNIz0F6jelRNkpotJGM2A3
rA+P0IyX1v9OF2/gJhd/PD2o7Pxx+rknpzFP/Zc3lF5NLqB0/vVPNhmeMo/YIu06XqATVDehpfkB
pQJLFpWRe5vTW2cYxVsAbYOiaGC4OZCfiw/syXQaaGJw1THbvaukrubEQuz74p7tiC0hUfVv5mRs
RWp6J6LHYU9bywNdxC8SI71C/bI/RcBm5uFMwZyVyjNQCukZYHXnrUvbhKmYYq2S+5aERKxwYDgy
727gK3MQ96q8bJIZZdDPQd3MAE9a/MW6IHoorY5y/lWCOqhChkGdCEEoVw77SqkqR9S2i/ZvIYoN
hweIFpDCcPRFtkJF85bqtem+HWH/2h0M+J+TVGOu5LGbmIlD7mYWRgQHqdV13Xmh3WK/0UClPkFy
Zax0MV3ous3fZQq1p0xsCLhlzGIqK9mNPIi6nNElzuzAIbxhabKlk4MH1tYAgF2T+QrjpIsaMvML
wSbJ1wbt/iCjIGcRZemYrAQBQ+bv+CvyR/VFHoWSgpeojjZRdosp0W+eKRDxHGOv9+w5SUyHjdUX
pzXggAWhxMHbq7wI2YR7he5rmDsVl14atiK+aSMJ7UiNCpMkdej1Rb9aIAtMuthuDtp8sHsWmkij
QyzBZUBUUENeIdB8NgT1XhhRcrOF4eVFnEA3yiUI7PEtPmzx7zS5fPnbv7f3qghkDaJC38OVyjPu
6IbH5yMG86huXXuggBYZ6t01jmVUXarGame/fRvd1+CQznlbYFS44Q936pmCykxxXdFLafy722qq
NouvH/Dp9GbBsIdqZ+9ncf7jOEu7TmO+k24DqDFWwAoj/DD24IZoCml+EhgTvXtNhRcaPiVzjLGg
BPPQdz/nRBRB3H/pokLIYbVmUjqyT57KOBDdNsA1HBzbeJEwSHN2LfeJ6gVYQRPQtb8X25PooJv8
S0Fnh9QnhJdIzfciq6RSr2z45jD7hxJAO1gkrcfCKTRvfrdwIWPePZcDP4/REQtMvviq9o20wu7y
6KkKq1zqlQLyi1bR7DH9ulV4Bw/2VzYH2ZVRdD6QlqQ0dD/hv2e0oRz46JRTsKPTMckLvUIngU8k
/iSTB9XrSCgrcVuVCb/iC7pv6s8LxXaryy8JxiQ6uLraKoyTfJgsxANTmrgqIS0fM6p8eEDFabC/
GG4YvrgOrJ6XbjNBr9ln+/bU0SB2pDb9hk+XF20MyPzcUxb/AE+maHNynrpveshApLwXXFeTXtm/
FqXLNGVRyyrcuWjpKUFTPbh+KLrM4GcS3JYOhATx4JDo3cQFINld4XBn8BbW601o+Di3vte/+Hpi
3FBYV2eCouzKO2BiY8KQCr0hNHNLT7pcMD03kO8+SSwaD0e83IteKf4xZ1Jtpr/ge68mi2SfdRqv
3w0pnnBgRaDaUiwZ2YtEsOnfNU8y1UUheXQOuNop155iX/xbgFl25JpmBVyYoeS+hFlSbDQmHCd+
utq7qTI8bGMjxnj3mkKK3YDuFLXhVkoKqFyEVYnZsesN1td00gyMxJpewNV3U9idaz5ELwR0fX3G
5h1U8RwU6aqQYUxrocD6gXG1M6UBNn4GIhAaDweo91pnYrdW8osPJOtON2Ou3nzDvE7RcXngz+Hf
ra4wNflP8ZL4cc0KH0awICVzLWL+bIEuo40oPnX/OXM244+H4S0iMw2ueZvtZVazPF7gU1hLHBtf
Lnm3guMzLAPt6VQIGHYfAsQHOeyTWTRJMLPQhL5Qv73ikUaRywcbzV/jc/NTBaj/dPuABoTjINKC
XQUYux2dJSbUFQuDfIc214sk1GusJsvNqb7KroiHifoqbmB2biLVkvtC1g2Vxm8WPwtKrI5O5D+o
raLIVoCxtbuf8HpNUOfUhizmaw43A5hSkB1l2po6D/gmVggRQKTbZADtIrfPYAM8EPasasg82BfT
k9jPy1FN1s9xkc5uwFOkUDbY27tGYsaYvLG7Rk5H7G8ouNCkBI126rYE0zvENHXwPJXlfEVCQwOk
eLGgeNn58EcgVGdmwAAF7M1WP0sCG1C0O89VAC8IgI4WePp2ibV3NKHul03i733fppXhdIrSHMhF
WieSqq1YCa9y2OAVmqDylPmNlRWEcRxK7du6I8//Z10qwR9JBewBLj0vvVRqjfbTyRVGUxuV0rKI
Az/81lfTU5/NvzTUKHr8dGakcTDUBrVy+xIfWSidALPQr0MEXAi/8fWpK14cDQjgYbGS+MJAcFV9
CgO87BPrqA0ASV7Qzg2/SuL8x1/fWThJAW+D4Xpba2PK2PbiPpldAJ1trvYH0hDmmjH96dzPnqMS
9NTMgta9kl36ruXa8GIdvJ4JSXjbdh1zId8KsjCPD6N6tzvmyr69GkqKBIUHpsfCg2Otj3F2blQL
fHuWOvzhZBMbfXhGLHKfiBKtTqztndDACj/zE1ZPDMsjV6LIt84xcfUkNqL5cazo78hUiMDf7vVb
e0iCM+S9tx+p0dAYHkxgnhzuI1PiwJzvSUXETWtlgo2rzE4uMvsk29BW7tOIXvPZG9d2fHR6owCi
9vc+0e2CNwMcSwams8HoaJfY7O6R0sp8dojXpZH/Oid+30VsF2BJprbLkLxSuo3Q3Lmz9OUZK8Ll
VUMsKO/lwC9GPEaz11anWOi549lQVQYa1RQ9kosrTesu/vNLUxpjvVp5qDnUR7S/7dAaVvucvEzq
ORhw6M3cE16RCnxd0iJclVdWLl7E2BTS0DUwOAizbzUZAEwe6LCI/jsZJmEkNJNztIalxMqZvHIy
YaDXw02fdcvau/eXj3Ad5ZBU7n3MYP8uNiTYFH0MDommuC4haHt/fMD3ZHaobYBWiD0V8/q76WRx
gS9abHiXXhKU1AeFuaK8BUt8dyRVdGOWPXbdijlej5bMYkFbx4yzVSxgw5uPUoc9bx0PZFpE8Mau
XvnX3ju6kfk6GPv72zjlS/c0ihysUJiN6r4gEvG+Ba92Qfg8stHmHdwvLqbJI3thgbZlMU5QILrV
mo9WfPc1IJn1N+lB9vHVjINJkpFxFLDZ8gPST1umBemnbM3Jjep+i/pTMq1Ae1yYnLW6V16m9O9g
AQydKeF/5feVJaNtVeSGgMd4XEaHfby1/ZGzxrxJNbKDyE4UizgMhOrgLDvdCY4DpRkApYVYrv8K
SIIrVzTWvFBADHwkYx6s1HJBZ5tgObSLTMYei5KJXoyhUERqtueNsP81wGb2GrheA5Z62MAncvnK
FeszrQs/KcFqCzkliJDMumQAD6/HG03FNDnNSXzdtQJFtuOBq+Q4E2GkOauUgSnxZX265jQG8BEf
DtoDFmM6o3LLNHhLG2PLxvjo9p6wyZhw6zqJ013iYHGfsPX7T1XOlJRwnARIfVbNGKjRO3ERt+ud
CzIN38xX6Tr82we/YrDBcOJ9x2CPm/KNNA49ocRawTly6SUvZXwV2XDc4YaTUf6LdBkmnplx1NE4
inIoYJThadm8ERHsmFILx8Jy3SGlU7WldoqsM+zwFXRttiydKK7+gOd9ziK/ETY6D81IAdsCL6iD
SjwtfAsLl6y9/cf9bJ5Is6oXsVXCbiLuvahiArUVdX+8s4PxDbkQ4C9K97JH7b4nTGRCxcsVOrkg
DhGD3EoPNdCiOtXUKwDg+gwxyp93mi/JAmGn2WfwKfIIlRJlmEXTCz/z5oGarwi/p2T4pz9K9fJi
x5kBWr6/FdfFWQvtw6gyNK0VTfBF4HB9qSDOs/GTZ+3keaH1tJJl5fjTy33+I0AFBWCeX0t3q4Gp
pTSiMd1oUm3Tpw6i67e6och7mtfFkZVtOuR4H+p+oppYEPT8zAvI+55wDedXLKfmAZOXdQ/ry1FQ
/YeNE6o9kxFuzpvMKt26daqayA1PrhHJ29crnbdtT6neg2RRLON55eYLXuYURjOv6px+tBf082PK
nNvsxvXaJ8T64hDoC8pVbOnqSD8zQeWN/+n1EgoAW8ErHdV+uiOWlyU354dTZfvLViCiiXdC8KmG
TGK5J3TY0f45XnJRlnz1AnKZKtBwi2sDSYMW0rK+07pHpEF7MZOh5eThWFhLKkwtcWEsa2CpjSx4
dqNHGgeBjPWjFeSQk3pLdwu8G2rfjqzEolQtSBvkWOxP8pzCAys85/rVYAc2Any+pj1NNeMiJx5I
lNZNjlytvdeTDBi9q73xsc6q8aKgSnQvT9+rK7lpX52BMTv/hJkid8a+t++ZJSfvyIUGsL8rX/o6
r0BXOUQROqWhEyucIqsdzVm0SlF65rc6ZA1EClewk84moiaY+IvrEGfXwybSotfTI0VBc2umaU3e
jy9g5xUqbFHexqTfhLoXmpGzAt/8Xo1u5/VwQ9NJ42KP1f0NJKYGgBIn+V5VoCLHFYrVsvgS3uHb
cJp/tCcllaE+vC2mF4wfgfyjNxWxwtkM4SLJAIvR8E3luhG6tJari/uAiBWV/IosGxqW5/5VA7iD
YDbSj4PB0bBYk32udA1vdap7I3nFjcGfQtVrT+4BVD99OoekK2gDnCUfmxtyJN1cEuQzrcIemV4P
vpNUUNyv1Ywchf4EzTmA6C2ikB38IMyEjtS03s7PsmQDx2w7AlmHCasC59YLEgDhc0sjxFI4BOFr
mIhtqkt6g3+WImE9ilJJh+E7xCb4zagogRWWOlCbCor1ACKy36dSUms06VwBfiDGtFn+kyKaVBBO
8ekw5kGeCmvN+2ZbUmr26pQEfHxrfg9GkTbj5sGNz3qgmHInfQ/i/K80AzWOC2Jq0jBWxsM4WqlK
Fg9v2aDh5OhlJ/8CP19ZlCiQ3aNn4Fnp2SJNOpIfHj6bqctoD4sFeSi6wzaC5dc5Ujwj13Od/I95
NrKs039+2B7ZcWVog0QrNWuCF1ia0OfpkpXwz4e2En1ne2aEmMOsADgh63kv7bfmi1m3XO9Jm+Vf
6lDdjALW6euKvNGJm779t0TcJU2w9C2Qfdma9ryhhaWG78+obwee1++8GjrhvWRZoScIl6kt3cxb
YoNmW1qZ+BRP17eB+1aXd2UCW/T1164qg6Q8BwZyJeU5aVDt5VjPfLZDESbfWegeXkckpEk4gJQD
LLtiXUkCH8Z5X6tzKTFtDc7AfsecUhGb6FnjDsHlaXQ0es4pwhN9OhZ+a+/VQgmxaW1zCuyCkihG
6mIHMOmccWp6TUds7rTm4PVqTLHDAYT/965qtiDgQV6stTp123pYDZ0KVazPRKZw9BWeA2g6+xTU
upcwNQvecUfLabHaQJg+2Dp671J5ac2g8k0Q/YKKfkiTxML6XOFsS1slKi5syptUaYz/PbY4wPf/
iTBfdgM4GomZe2SJIxEYvr/CEBu5kVXY5ntwmNBtN6/1M3rnR0xSdzAC4tYHlIPoZNmFSXZpJ2kD
4NyNr6PF5WN7AYI/Gm2JB8yl4I+7VuX0EO5NNX2TTKTs0Bpsrx+bW8ms3eyGwpPl628LqUkfAL2s
2ay7kJqwAiztg79gsdzyOj1VdnXYhS0t2zrrOoQfWOD+NBpug/RoqFgX1mrJdL8Z1WnqaN7V6LED
qMThYla/gHfoAOPd/3zp3L9hcMtnZpMXRH+SO34ZoKagLoXlmH2DooGtVZo+rq8kUc0+rubd73vZ
A10YsOLkKmMZ1vtsf+K/0ySF/oYF9Q8sjyV+TENeIGKp3WXvJ55qvY22ZZ6nkxfyUWemZdAJxWdH
FHNJzEo7/7eAM9H9qS1OkPKk5Ol9XnrKc0zvhS2CdZdyL3QVP6LOZnS9uL7IzlRTudC9Z/iBgi76
SFsyY6Xfdb3AIlnbxtY2CXPlgQ4ZTeFhgxoBgJCiBfmI0XhihGA+lYIFZKgEIi0i66dEWHfTyTvh
9s7lFoc0vJx+9SpkiPsQZciQVuLzK7IjmsyWcPOR88wKDQl3W3+H5RlDkDTkyOgYbAXGP0AQuIFL
Blqi4CznOBqZArERrj3lzy5Z1qaIzpQill3GPvCp3eFXwv7Lc/apKlbtZhx5oA4J/akNiRvAtpA2
HT37AJcMghIeQI5yrzk99E4AKHIjVpjVNY3GM+ka3EdDmXgg9Gbnv87/8MEeRFaxa9yK0FTDLAo8
5M8+DAkMGmJnbx9+gEBaTVrevOXnOaMGoA6vfUjwI2U9ax2hkiu+almatGYsj51fOliiHo2uiBzR
1u2jGwB10ya2jbvB0+IteG1dk09gcx17fsXI7fJrMQTR4f3uizxvOs75CVp2dd55El2m8OqpzAFC
ivYlydWbghY1EXPJG13r8beWWEcuterAv/aLM//3Ckzv0aNcicB82jOVNhID4bv1fclKoCjQUtDt
dIijYhrYfxu6lO2/FAfY0XXtiZqvkiY3eSrqkGi96JcQaLqRaYw9Q0t0Uu9tBRjnfkAS/FTEFEkk
9JW5fV69+Y2EtcqX7LhrjiJyI+moTjDRe0ewPfRGOl8KuxWHgH59r8hWa5cYvRzkCWW0KEzmbari
rWf/a6KaXlCGaLTG8dFzGJEIDutQ2pSIVCU9hkich5+0nQ2OewDmJKH8vqfX45xhfXfTlUP8Kqyi
r7pPdYzhV4b/3feXWetuM6jdkvfL3goiREABNKOEjlMWOcKPSo0nRE6+vvUPcnKqmTEUDSQsRIeu
kfAbrSlHOTLOiugm4mp8PyQlMk7gXfq0dFSyALJ6FnEJjY1SGiD1f9OsO5oLC2b55pvmysPkNNCq
gRxhRgkQp/cSxUs/6XD0VwNkH+ZUKnBwDDXsXePO8Tf08yvyJSgvCOgPbDNNXkhlPzY3CuLuw3F8
yPYijyVW/T3RKBynHbfBtJrE6sdRCdMuUGCRlEZRxNc/wRHTJuLeFs/98tYC6MbyLWsS9TpNDtqx
DcQlnRGiXNdeXmvkM82VcJ25fcCVWQ6anGehk+XCj6yXXsoFEWQOlTItXCeFSpa/7FL51MOnp7O7
NruVVpY6APZf6ZBGuzHkBhYXtYQoPz67tS6f0fjWNbknAp9cWMJXLAyCMrG8qmOzDrVNGEWVgxce
T0/g/uoUHgPW6OSkp6/BLfPMC1o0dSGeNGgGMZSQHdUestiW2aFAT93oLaSdVzzpIc8rCY+Twf38
vybjj0LhkOOT2kWI5w2pK2MoxYwDMGT5ThHxiRlDMybO9WpGEGDtRhrmPsCzNFUV9OG4NyzCzi5K
fEEGff+o91n48ruTMQiyTfEL7CRFllKD1NanyDbKW406kK/4p8eFJ2gTQmYEknyjmdnPQCnfZNNC
fEIvUePcQ2Z+a7S6AW4Ax5lLB9jKdlMI3eHkRZ/+SWcgVUnyuw4ur7OrM1TupfHe5szAzifM8HlU
3oD0zGIySL2eVdEWYAnFyEtAGXGCUa1eiMqu7/HIuI610q2Fit87l0Euh0Jfpru+uGW9hQGgzSJ2
SS0swUBWZKqdGO0OULRwfpyokxcf4BGmEfWpOma8MMYIpmix90A8Nq5BC0YQBNUyIrYeIbs71CvT
33wViLeG/tCyCWZoNl9VIP8hvxH8ZHcK5w1Z1Pcv9H0zn3KDq4+UMOwBaSMVjBsbz6QWJzUvyEFT
jvYsLHHez0Y2rKiTGfASFVN4JWgOaIvtaq3WqySq1MaLldl4T9QhCJCyRAqHkCD0g8LLj8C4C0Zm
nmiAkHAxcWuTtkYyhvmvzpOI6AKl5YdRM0iai52RBHckmEMm8oxpAta3N/PR/2qIRnDB0TvCwy5H
c7t8xd/MQhXK8x88nzePN9NrBHh/4s5R6umE9oz8w/fkfiJVNdDtByJBasCvVdHzCsp3SjFjoyus
mk6Hw9LKIKeoHjmQ/TdwYrQyyIlaBYjdeWteQecYiKSscANQ8ZUDTqgBy3Z3qYf3bCrl8VupWSoD
uuPUM4jkcXDWB0184zWjzgIBns7rlhLf9eRgbaciB2jAGBB5MTQYg8vp3Tlo/ar8TqwQeT3G+HKw
k9r9OB4/C4paN/UGvLyPNIx+WZ/5qYoLLD76KTma+Ky2hhmKEBGO3N+mgDbptaKjcc3ReiZXGzZ3
EdaepKiTesaKWwhUnkFijk7VN3NstKYyUHkXTke7BOCraMqArKuCqbZ4Op3YHW/AafKSbZFXgC3q
MzbtdoMwzjNDpG3ikYiSkzHROwK3EMTX+c6ZGKL8hdE82P6wmzzg8OhmsyWg+fK5rOfLYK/Ldnkg
QE+freCWlcM6wdt4RRTHWd+BrHcxe8DTyWsyUcri7iUS4bcbIINV367MUssHx9Y2fgY7z725Qwg5
kznAooJr+SXdHK2pj0dXzPn0aKQvqi0SLQcrGi7bS6YTFd4XV3l9n3GtE+uurluImbjQ9YdzLSxQ
LCD/8pmwHDc3zSqToSJsiDR6u7S65gC/bG3kWR3FtwMVcheOzaGQlZAvWcWYIYKLyb0MF5XrdnAj
7aqtx3eR9XtO79e9nW5UZMveaNPvNPG1yDtF1A3CDeT2dn/3CB9ORx2gCAHeVYC8MDnSvyn4RfmC
6uqQvnsuSQYC7ap86dD1/lUOZ83gErALvxtyck7LZIhC5eNa6qV04N9yok6EogmKqZr5z9WXWIMO
1TrG65qdevXEnazN01iLU/qENsksEywIw7kb65ybTzgtJ23CTxmoAflzd3DsNpC7fJWXC790rMz2
on2Dgb5FIZzAYw6Jn8c7s0X0uQwoT4h8pzgnJR95FXMm6x9HeZPwDIfsGzd0W1bq+xBildJKNUnL
fVO8X5jeZ65OXXLKSl9Qj4cqMYdexRaRqdY4kT6szsO8N2bLuCCO46zrtglg5tW4XgNxxqTOuzIU
mGe3MUc+6IORg7zMcis+JbtezWhN9HwGqHXMDgAVSAfqNmZSmqiI83hmeryGGVULWi3mbhHHYlsk
EIljk0sxgKkejg5iKkVnCPrhCGFjl0hPz6ZiVGKfwtztzxSFDzz8m3AMIS3EJmYIEglCrxybExlq
7zvXL08Ww1s9PFEejbbJ5LTDmA38fHuGTPoltS3v/a1im6CDsaLfhssPUB9OU/1jve9wrHUflKHe
gIsQ2Qkjs2IhPU7Yqyru0tGUH6jp0azFcCdR7JtHbqCSH5YoNPF239D0rXcWrWOjpe7aAPUMU1Wc
qId4adkeiMA1y22R441q7IcMX0KKxMv238jZTEtQQS56dwsqDwQmYkBSSwlbRR3Ve0klEhjKzFEW
yWk0RAATxuhcjlMbVFM5ajIf9uzLeWr+C78VjYkVbGLY+1b91VOs6bsyjSHLvOT6tXTAYDQ+X4BZ
ch7ZYVmMnF3fYlr17OPcmjXjmOgdEYAu9lr04TGwSqjty3xH36aSj3M56aH4CW/b9bb0TIP9U8vn
OLe8wLAW7JxXWHfKMLa+pb2X7UoAOJhYrwQ7AIjm8aCXLH+Zy0t9ue9BZ7ypSrdCc6x/viIrugCD
cLQuvr+dJ9d3JEREvCkvOHMjL5VetE4AUW01bJBuL/vEgHjPIAMJ81czAuwzhdqm9KQb5YKScFEW
qKc+ceWXGuLwVrkvgI/uPdh7C45JuGpLW5aWuKPq3XhS0TvR3m1L3x93VnM3MVRZyFSFjquZvlX/
EwE3SBfXSq+zFhMV7OZKuvMMK54Uovr3ePLJECDl5aG39grUSQvseJMtITCmpRYFshcaJOzo+nYK
+q2tonRu1O2ZG9s8y0OLczYIJFqatSHshiTAuKs1reDWP4oIyLi91mQ1jBrw/gaqZV7IDtDW3n99
r/NjrbuuAFRq9KN0slW4ZldDpQJsa+102x9iiHjqdrF/GjX4f6Ar049bfHsEw3IUrPXqdfK6DcXJ
UO37xBClomaIczT1k5gL6MaJPUtA5u8cOP6eabt8Z+mXMWSAm161x2UtPb7/5CCN5oQWGi1MVAYm
LD0VC8n/K2SYYFauhDRsMan+T971MBuYZ2c/pnrEsrAY6E1CGPb38y8apFi8Jx175pJyeoY9Pl5V
L9QLBBfYHeUOqn6pDrVxU3d2UMvgHlr/uaMwqu320/iTorg+i7Zjm4qly/JHZz7aKFMDDJTrWR8b
cydncggPLewzCwOgvasLpOquBKYsvN9GZKiILtak4D4Mlc6YS3kN6Nzz1GmnTyNX3zT2KRig5AHC
kwkUNG2kw+L+9Y2eIPfVBu/hPum57LNMLUX2p2eP6MwjbZY82GfJ7/Chky0jw5LYLx607/WQW6oy
1UdUhHoo1ztGGZ4TBZ+tHGtjabcvHfL3r7z23oJpKYQOj7fk5LjDp86Rhqncc8HySPspjcCEjcJE
giKCE9JYxrw9eIlMNr5Wlm3Tz51qHSR3fZOSAwhk304tiTEBkv80WeTPOJTPTr938Ru62kOvdQmq
kmnrry4UeWnq4bf0Hu6iQWmyGhTPxpfeCH5j+wJfSHMysqxZpa4Wv+X4Jg0r86hGEYEMdqW0g6vq
xRTZFyl8P32KyoC6MYAgRA4r4knn7DA/RMxefSrQRl5R8tntSj815W+6WuGfBdSLS6/JcwqImeet
qzoU/paD6d9iZZQd6Nkyb+ESKcK1+XQ20XP8EI5drVetB/Vwh9Gjd4/K2z0TYNdq3oh97pOTX3FX
QTVx43ymG0LnKA9aB6isoGjrR3O75ZUecdIgKl/VA4jY7u2JLMpwJuOUVpWjt4ENsUDvQ00hT2H6
TtR+Y9P0meef8GYN8vsr3JN/F4j/VAdYc9psE6c4rtF3GYQRkEH01bt3Xo2VHaWp5GQQwOzGIb6v
c3+UDaSxaURSZkj4WCxozDh42r2L6cBEs8KIpzNLmMM8FTKaQGNxoCbRjuFkAYzgDcpo7nWQg9m3
VeeVulusLwI9P8FtKfKlUtGeIbyRIjLL/AWAK6e6tXJ6/3B7Ppl2qgjFUBlekKhZbOy2dMksbq/o
htLLoHxMNRAk/FO6t7wcBRrt2mx5Neuom6SApiR9kfVYBIFKn4q1FbCqe6Tk9rf23dvCHanTilvc
5BaugFhVubqvbWk3k0B7Y6afmslKrvN1i815qb+DWtu/R2Y5ErZJ475e5QOTbOeuiZpOoPG2F7D4
Tq0Osbdcu62YnbDZJCRmtIxQYZ2rTv4ABmp0UINlRPESnNqx27OBRSKG7eNohZ6PSFjQJHpUspuT
9b9Tq1GEwxOrRzIfOvKdeY71xMFUesxO0EYUTAdAmiXy2tQClXup6zBEw7aTUyta67GpzVVYxdv8
+KiYuE2HU6jEkToY2lXdD/JJjfdEfp8o9CrWmet1gaLs2L1QPGnZl79ETq3D+seSCjrdZtWCbf2c
g0HQb0UTL9L3xFcKJd2eip+fvFRqKVcNTiIRh4LNqkdrooTJ8l1CPDgkkbEc1hbDutDwD9ieRwrq
mwUP3XUc3XZYV4G41RZoVEX94lH2RK44hy3MDjSViEXhiciKQZPM+Z1RAkUJe5hvHPIug6i5TH7G
xlWy2hxDvw9+i2npbYM4yw9lo/dVaWH0e1nO7EUQD/0VSPoBLggNBLJ8KWvWhMpD5bksWCHTP6XF
Z5PUXu3c2xaCpMoHgXBeSFkrPFCf9XW2ilnl272cut/MvVazDxURPnUxWzp3WOQv72CeuRmosK49
GfFh8mS3pdcgOQDqCK4aubHrQMeCcG3Jj4zsVRAsdltuLRhKXhQRKK4xaH4xKwrsFCIBfHvHZNpp
a/x7U/bLizQBrDyLgXg5qMCDJ54DjjAJMYSMWsYzbMrQeZ6pP4JKxIbi9FVAPhYLSIvplaHSMGBD
pktU2+2H4uts40xreIOAHgcIlimxPd0PQkN6KnEDSbICDVfLZeXdOBi7zxwUw2wQJJEXJFc149nT
248MWxOtw2PpDQFWzMWghmYAJ8Ona+Y6xkrzgSyQ0CFzIe9aRrWlwv+ODyRelAku07494yMdNQJG
5dyA0rF34Pmc5wEcyRvId74xUPgjmidLlJG9RytFia8pAsu6uihSJymNOlvi85nWq6/esz29OBd8
y23XFT3X1pyMxRBWrudsldiIHDG8wEVIQZE006sdRWTt9ffbTAnAg60ZMdgIYzaQqG53sOeld/wH
j+LcG8QrQK2GBQC3njisokwYebzMMsx8/fhuXYGkfcbjKJhOZpmapyA6FnwKxgZIopaW5U94lX0L
iji4aVzCrzU85OT44+KPGpDAFuPvxer57D6QHke7F6dcErif81qmDPcnqqzqfr02EbtiBA2cGK3P
guGURquT7MNjMP3UdJkKix1Wjjio785DxT7RwCjSs0xUlqTid3RKrVHJfRLTpBrQzv0bc57/YtX/
QLb1iXgVWkqow6ECKQMFBvKQ+bjr/3ifhI0De08cDmCYM+I8Z05Tpj9ymetJxPabPWc5EJu9KFPT
mGJdoeeQf/VzEQqbbeAQ96Ou48Dn3/gaqiRzJ0Uwhb3kWePadNaeJHm6I9+UHIzt3LfcRHTcR5t/
5avpTRPPmzKJ6BpTlb+1+bORMY/4MPyhRLrnJUV8LL43z7NUDjGr7iP7b41sA8yReXzpCLLFaLBk
v1nsOMIsI0LokzQipU4OcLpHT49bpgxfy33kdzKzECROa2XRA9vGkAzanl0/Z9zWxshCOjhz40cE
GTcKaUv1kLO1tY5YyBVSDjKbX467kd9VN/Ph5lQT2DO1/X7eohfVzDoiYRxLt667sjfdHYn/aKa1
OruVOvvsl5LUQKpBKikhPSpz05e5H/ZTkmUFebk1ZNZEM/P1Qk4qGJKSbmjD74aptr3ZSdynGrIJ
1rYWmTgoaBFMiGMF3Pelw8cH8xMI2ub3y/j8UBHIcGooYPscaVsTk7O9+f9DNlnNH8+olDJFgFuG
gJl49tH2Bxipn/uNsXDuSGOka1aqA+9R9mzVDPIQ7CkfGyz6y26ZJvSZKs2afY9XdxrZgP+fnRGw
N2mo2Frmmdqo5+42ecU58jxqMNxVwx2WiGmY26USLxEQERFuBHz3oBPvodtBir9ZYQ7bukdQ10GI
w+wKud2JiJ1oFeoi8a9bOtsL9O179QlSR3T5afygXsS8MViHVJGWWrhs67xx/Y0S/L1NpfMo6kPK
uU+U3HcMhrXLFpF18GCiVqLhG92ZoSL/W+PVQHQ3CYbP5S1DbrsHgfT5PQrbxn9xZ2BIdNrRn+Jw
/3wm52PDNQakl9JwmcHsPQNg6RDC5CNTiX0AEX0givA1c3wmCWuBDKRUIJCozDupUb0ByIE6cpDw
nMF5pmZ1oLbn1KfJIrTvYfZuYaq6gt3g4PIGbKWMixlU7+typeJUpI4XxnIuJG0RzcLqXc/6FRvL
ZriCPf1ZgdV4UcuMzmw3myxDI1q4bHxcX9kRlGCYZEXwjHcpSXgg+phz+CtsUU1FTR1uNVJP7o5J
lYjEnVZ7UKrqvWlDSbe+8kHFKVQgxCe8ye+uzlcCIWKP8ShKMcyKq7RufkhVsoDjHdo6sxQzfsev
/uatxZ+NH6LycTja+FLuPQRhD8BY2g6K2peFlxw6Gfejg5nPcSLHbgbRuk5HpoipJ/7Q3g1qcmyO
cKf5vE/QEDtmokqXEI9pU1k+yB5DLCvRhVd1mvJsUyccPvAaFFHaeBbz+mPshxme6PrMtBCTaSaT
q7YP6cqXHg4RSkBW3lzOQcLaCmX2j2ApeGTh4lKlMRjfxmoAfUsrgyOFD2tT0dUbK06h+j1es64k
6NTkWL6FbYTx02J2gMsMKIO1ZyN4L0dHiiEZBGj3Q13uEHnwa7cKCOJpMfRTbWQsoFrJzifRzVXG
hVbtTSrT1HM/osEsaNw+GCepVFFN+VxHWDvlzmpyYsS+vhKAgtacBo0P21L5d71TKt9FAoeqQ3v4
pvzG6MwOCr5x7/zX8Amu68ONF9ZuARm2Z4+mBdL2PKAx3/1o7e3Ys/2b2psDAzLYhUCwI139vduP
2/fyTdDPXJzLUTzOcAUDGV33HRtsmcZZuJ/+aSrajWl3+QKhdTiGYZo2gG041helF1kn2jr4j6Dh
mK7n3AZgVJP61G1tRAkpA8LWTcAyg5kqWMrztUQg3M7qZKw8ly61iFiidPj+tNFIVtgPZG9OiwXh
OzhjSwGbrbOyUfOlXDyhRfPlABXS374gnxieMJoqilt3DLU0l4iXiUpkCXEZFMNV9YFoWG1lWqQg
5Msbge2Hju/7DJ06e2xDb3JLfFNzfUWt+VNZbqClpIgxydxQMQR3XnYQbZvtJXHc1y9ACG0CWdKz
8JK8ha4bzJtPWY+B1Cf/mknDzgLX6b0BkyfFJlD76Xs1iDrSnkaV028mLykGJU/sVaRqbbsd3i8M
dJ9j0UUKW/tqxJSKVBX8605D5OH6XuFvbFUwdUDSvru9h82jMMTGVz8x6BmtyxBvblMYWrXvXAvO
4EEVGkATyDhs6K+R47nT3TtmgRVuLUJkhC8LSPf43BHEjru6nYrOT+pTja/EDQChYm2s2WGcxxA9
mfrx2l/wklkO1L6z2u8Mma0+tfFgdQYXvCu06Xm3CVu1TVfodPIhw7D0a8ZDu8Dcs5/iHahZzMQl
88XCHzNV24xexQjviAoDTX5f+YYe0DUOHI3qcLlf3MSRaDun4AHaiJcZvP3rmLreWXCAJbOcsIS2
8sFWup3zUpdRrLMnTWdrk+e+fYy3id7Oq10l6xqGbN3NzsUzlDwG7oO8EoJm9VWK4MBr8hPCa9Kg
SUmm6QdZ5R3OvBtu323G5PovB0QOnHfTnqNLZOZYaikiZTOvLpEW8l2ipoNrtGnOHA5cYT8LtuLP
KC2cN1rcq3cr5NlGoFpA5xFYdwOsSsNt8O6B4nIutkzdi7Fyp1sHu48LDLaZ4QOkcY1+DY0gIKFo
I5m2Jrytk27vT5451W9MWzT7tPns4/LjLVG3yygicYW5gGWMs6hVZlAuffJF78Ahwgq5SY/ljWZW
HmmKDdQBKgmHIOQVEjjTEfquoNZOSqI11SA1KJQMYYlBv3k82Kb5WexSfxogN41VrPI4kS5cLGbq
IxF2ylb08JpCmDaE6kMmZvZPx5NKSAdaIdyHwX9Pp6+mjFgWE1ZukMbKaG6QLZrC2CfD6W/rYfKc
WXWMHbfigX0GwkSgIyBLKteZbVsI69cBWnLnXB5jHzdreC9ps0eewoLmibcP6Vsm693oWOUkhqkP
zXEVZScQG4HYvi+apj7A8qt+3xV0VDfBvMLIhrNKa38juY5K+6lISLdhJP9KdA/uANrghPwSMJN4
1CEzr9AWgRIu6ijMf7MmvwkqignwOy8nRmL3tQyP882//iKLc86tY5ohXaZDAXIznDM2sBVWuaTQ
gq1846GdcEv/Zc+Bz8IMe/RLvB7leaD27C9m5jlkNWeLfAnxmAoUoFOVu9nmz59EJUJdAeu+G/SL
7PuCRyCYBOtGI38bDmcAMyYsDhDSnQoismyMlJRo+7rSdmegblfE59Fdi4Ord2om3UFRngZtezSJ
jK4ccl4GrCuIa6ZbRg3Gf19vystWXPSFnpBpC6OX+1YmL+7RgX/Kqs3mgDs6xwEDLxr6cRpklbUw
4VCPn1+CSUDIKgpGTqvLoeh8MCkzvEbbRbswJ2MKjqO8uJVA9VFadKt4MoW9MP2CKSIGIz/obouU
hFfxfnYTJl1BXQCbbaP9UK0kLErQG+wNdi15RFQzNkUYTdTvOxEke71AYCj8N31T0KEfPql+HIXp
oEeLwfDmLbjUyQ+0Sro3zz+AAKdluqKnX9/axc7cTnHCBhwenPqRw6zscox2lV/DQbLIESgwwc4Z
dY7u535WGHjCPDWUzKvQf2udscO0hL37KVukmwo0DXXAZq5jDzJ0HxYv4DQPyW+RWhokDRnrpAsp
eOrmErgSYMwvlB38Or6WJ/PPTtFcSITOk0APjPDexFnVswJ1ytwES17LJ2Bzwf58YkemilNUtE0/
M4RkyJU7/s++uyiuUQmMyDwOgI/Yk2FTEvvKjJL1CZYwwn1wOlZVCffpu8yj+T1ChtVY6I0gtItX
q0wmh/TcFntxPJvZmjjpqxD1TD0cGhhs7kTOcvKOWtApGznQIqeSz4WICNX688LH4CLXPUhO0vfy
6E5fxf5QK72dMTVs6zBSxb1EzlTgqwVhGIYDefbcd1/FMhie8EuUiSNosoMnhIK/dykjWCIRJlCi
lM1ZSVtZE2R4T8Kx+19B1E5+UbxjvnXCIk04dSAIVCfUNxwsORpPaCLBtjkCOmjraDMV1/osC0v2
7bVfXeUhcBE3UJP2cpW8bRRvW9k9emnkOlxCAcVaUxNmPMZIDCMLGocK3EBnCblz/KHJ6bL+fEIP
7fH4tdLibc9q56gcLm4nE4V2SRHaCXy0UGlFv6DTc2GV9pofIEu4IVtCB3vA3/VAw2EYdH1N2ocX
INk8xplHJqAJNzpqWnzXFEpwxGxSPq3V0klNgyh7Xb8DXBSJDfN2Rgmnov5OnkR66aMqoh4ISq7G
Z5W9ccW3n9gJrrEv2pHhJWAjAD5VLea9bHoJVlbTXEAd8SrQSdA3NZ7qP5OXCQqArGAQ6Z/yJCO8
uZJItWjlZhHdqnH4fB6kjCuzUN4/QgD10ZkvAwlN0c3ynghmeN8hwlORfd2DCvEwz3pF2bceRToc
9vWXTm3apAfwcX8I2VkkjppOIBhubb5Dfg1YPxTej0KTUD3ZAnioIvKjk9K9CSa1bh1f0bIOIlGQ
64bO4uNWzIT2uo7+RssJkNjoogYAl9rus83OW1EnE8owAyxvTUA9vv2zL4JNSawSw/bEZS5L8F+5
k7qjNKgucnSGdzFL/Xphq2ID+HtWObMWv5Zc0pk23beqQzKB7/P10JPLevZ3ZJwxeSP0ZJix/ezc
oPg745K0E43FhMAfG2N16HKCnNFU+kbMC+l+WWtFBJ3hyYs8O2dbafUMDf0Mlj8fuQUtbXAl5CIb
9N7TdipQNjBsPjyAXjmPq0NCWGkvV8213lFjeLZNRz4NwztVaA5a56baBxwReXR+rVw3eHWITT/o
DjrKQpMbbRlU5YjL8Xhi1ZlgGCvBozbeSD9+AV6toyr77D/QlHQx2HEqTPe3t7wmP+Sc8FddlBKL
7Oa7qwsisGggztINc6b/cbunEysS4rUVyWf+YSanrggOQBwRGfmfSD//SSQhcJrnN2NUXG38SxuV
xKqTIXf4BHR0LXmAuOaR1v/AI7fLn9LJkhQ8FZvdO+M2o638A17BI3iltXlCYG332rwYFqQ9n0oc
MkAopqDuyino0HF9ZTalrLoIyGD37OUqXsx46i8M52iomYUmi4x2oIF9qHCOLea/USpwSE19gFrF
PHlTXqTzRAjN7Ee/aZdAyUwtuPLyWTcGcArG8e22e2u3sUtUUsCipdDfCjujoALMOAOjdOdYaplO
qk+2hcF7507CBjCF1HAW38M5COK0mYPIjJEIXAE5G0q+6G65T21cnbLKPZKif+G6/myqXqH1E36N
rxiVBUOSpVIp1Pe0rywy3+AboFdots7xIKWkUGeWElQNgrXRgNg8VjSxPUKXy0/tqH8byLOjI6Ju
dPLoVtB3Jv9TsuXHrGyzYUHGhNPscl1t7dBrbvJc8Nt51vzFmwqjq2nokp3hv4JnS0hF8d1DRr9b
2RYb7BqgMnALX8SSWY9dAo8e6FTGonEEjVvsHy9bfi+xj7DFFciw+VfVAc4ntotyffTRF10ORpse
Rty7mvenzszHb2ipOYWjSqUJEzZr8NzNIrmmV/PtvpHLXV38aVh2hFnRQLouA1cofsWx3yre7B4b
ADzmocrjFim/9BjWLCa6MIz0spR3WytN0PRDtmAR/zxh/v1xISuyOj0Fa37jXKgem7ff5mbPbxuf
E4rtYQL4br+JOfjNqYhGAgd5vt6JRZYUTPPs+Fa0eEglKtZfCpFnmB+VNKdo5eQj3FjONfFzyqff
LEl2esCiovwlYIvxiMuX11v6FH6lV7VyJOak2tks+BH9ZX7xIm2sB0uv+9A54Gfm/mfGhimZEe7h
zkTQkFSOYc/RDLo0p8EE9Tc5fjShb4S7o+471v3x7FHQCC4Ty7GpDVHLRdJ0LzSb6ApMcjTnNwVT
qf/rTQ4NOxx96vKgwGx4BJjn31iYFcxjwZsKcs6p4CcBipT0aRTCKbwwXEs6sfG1+JhTFXOa7Qss
smLUX39MvhZCVRYrBxRvn9zXKHO8IMok31i5ClMVeenx8Jv0y/9imEBiEAahLoQxRzfeTUD2BUao
woGbAqSALWONOWxMKSO88XnSBIcuwLieMgwpQ/G8uU+ycpW/HJ+WEb5Xi36cmXjL3aa7Gz64n+bS
gebaBB0LLC4UoBMpzO4YoGlZiEkEHb70mzK+aeho6/89zgYvMGZOOzGSn/gDAd2xjG9b5yUpDDa9
4ROr3ilY8Ue7tSJlXGqjscrKNePUQUp7GIuo0ZlFTrZxpKAB9/s6v8x+WzILZBQZJSG6hUog+Wo/
UrQyMml+hmujdgCRZ164tViTqMLfhJk5MiI3VJZ4qLmZKPQclov/lPT+K1SzbZ7JzDeZgLQRcq17
yP7CdfkyJBa29+be2FY4AEDAUbfMC2pdXVHKC8cE06phsOkS0epeZ10IKXGjWHGxIHFPSYP19FQ4
PnV6CfAIz6RcYtVz6tebSsPoTSxEYwWm8AWStncg2D8qpkO43GdznfZbsSbVyrRLSxZepBPZQsBj
VNUWbNmd3gRd3Ln14AHHfuC4krI9xRUBV0EtvFpN7jY6igtRfgbm46zJb13WXfDtubJ9kxMO09Wn
p6lV+GmG3h7YrWnhOsAKnhJEIeayoAPdQG52S5D2/2UTfQ+ecTCc0iN425Sa3Q0Ck6qncTCJn6J3
Skw0k8GtQO9MwR/G46bru+uITQ/bqkykrqSBVfU86+tJLxD24CJFUIlmeZpDEzgkYkftWkbfMtfH
49zi1nSrY3wqCJ1+v+0CIk2dUOBmsvlMKVQ9XPwrlCOc5V4u7bTXBzhRvVxdWkVsM4fwWB5biin4
DHxYHOZ5+7ZSGN03IAazxfG8um2tpPD8tbvo1q3cJndp1164OmJmUv19ML+P/ilRURx2XH6Ttps4
ASJlrtMiGFOL/xE8RbedtIEtoijKzj6vS237E4A5epv7xqALuT0DSnjbNkE6XLCvflrMFzoI9JuI
QREnaQ8c9fvUiyoMxI63LCsS/lvNcAzaYcukEO1fJ0urjXRpagDL9CzdLy4mI2Tyt9o5e4m6RLXj
k+Y4S6/1yNfwBC25PvnIWDypfabRrmkbhNXQG2M9dRPFhQXoUrm8tqzCaRC/BE7/eewglz2MB9/F
XwXct8CXGlFKIIplaIq7EETlI3h+FRo6bJHfgQQTV/0hTOTew6t+1JPPRluOizuh4MbMI15czE2A
Gsg0lsrz4xvYyAXRJQ2EavBBQ0jLrPecHUCI4pe5sd8MrYLmDAAu0/azysVGoojtm9YBIOhiDthA
O0RJTOQXmib9lsy0qAecdHCMvjo9Y5jKkizsLepI4ydIewS8Ya4tqCjywxr0mSG6z/I0SjLHmJa1
lJIUFgFLGWYH4RJq2/yO8W+ReJ2LlrcEEE6HUU9aF0ycalqAEbLa2hoMxwsjfsp4oo5nsN/pTQds
2avVwhs0xm4QoTjXOFzK9Zj2w7HwgKrTGWo/dJrkdkekcuMYY06Z0PpB1gkT9gxrj+yKWr3BuWWp
b7wEA9+/MVTmXSkRdJ0MrDZRyW3Foj51sU5fIcbiHRVWjbUKKyiKosuYW57oNE6iQjqNSfVf7vT5
o9M/c0aJGHhphnAve79dv6pS9Mgf5UBUFWBcjQhQwYUDLG1kEO/kTd5IZ8cCip9nGn6gAnIPaWk/
jAztJ4O6NJxB+ddli0K2mC9xwBLoCwHRAg3ElqofaLnizL6Amj0rqKvPhFoctPueUwoDDAvfuDE6
PktvjfHzPGY9xgHuf88Urk/GRxLgb6W4Eo5dy8Z8KHwVEpDlVwLwtRJGLKN2FDcJKTF0lymG3ExP
mMYVEAdbm8tHb2mRpHu5WwmVC0oRSwG/nIbFCIthp72wQU2266MdgFcLFACleu2NxXwBf85Hdzh9
SWuhpiYQG6tKq4bie9aOGnlZ9nUfCfDpbo2T4KC7VErWo0Be3W7I0apl9dSvEU82QZD3YImTSD8i
9YO3R4tAnPc0Bcyng/zRTUvfDrc0MOtRJWnRuWHJcFAiPlMpxkzWIcSAvEll0wSOzhIgnf8xJ8r5
P1+HIshLZFetrk4csvFo60pLHGz6nrBLusf6Wpb/N5LvTO+K5KH8oJyujCNbn+EN5Cw3MO8+0rtD
WTmOSlkrwTi1LkC7hw78KaVFk4ibvQ10ZDVNppH9LsbuTF3eroARk0AM+Jtmf93mOtfTZ3G66MVN
OxCs/R+EU6YZB7xGa3kUA+ChIxqlK2he89Gcz4NSOhAq7HcqiaRx2FVsf9rGy4LvQ0Ykjs3gDEhj
n+oK0YgLhs0m0HqXfG2zdqwV6G/FbtfoL+hHCAFVQbeb7IW2HnRCBC8VcwK7lIlUC+/+6ebpSH1e
DF+51mKd8/04DTPL9UySvelADtBmXBx5/0T2iO/i5maZUrFvZcG6Qbg7BkKSWaOoOd7cH+5Jgn+f
rdpoe5T6VHdwavkADq7pH+gUulzds6c0znqjfTXvPNp0yOT5EFspj60a+0LzJ8X9Z24JHD96oMT1
cWmy9rlZ5nrX8qNYYnXdIl5LSgqkxGL+ZQbyUkBGZwXk4oHMK1DLLru/wuHrMlF9k2Ao5Bd2pzQK
IvOppXGy1YsBBVMgHV2aLjvpOXfq00/91FfsMtk5pqC4NbPRUIRQjuPorJuVUDVGPECZn/6BjaMM
TpNZ0GJRbo/uvK0yZn91fttCtmaKvJoC2tKFmDVsmLRliE4iX/uwrQlHqbbC9+lt8w1iSO24GJUP
GyP+UWAvvfTzaPvYKLjJEMBTMrWl1hFjsC1DYX7F1ALh4dvBaq1TGvT6LQhPOA+vBcMBJ0ay2btM
KJegQUqEuFDKIgjKXZkbOEdNdLm2y1tvHkfXdHfhhP6g4dcH+HBXXvM+RrNsAfwPc44RurLC8m0a
t2U4QvDbEUq9UwnaOkSJ9cy1/kwfrgM+Wuyygi5F66hd3EIWtjfDMcNc/bhTf8bJB7PyWBT0IROS
00OnzMi26T3KVuXkqOOIEeIaaBhQb9MbpUxc0XsFCxlWIuk0nV/6zfvkmdlR8B9QU52xo8JKEI/X
2JXP0ju2G6gwJUTJQscMzAfLtldM9pMwvoML/LbXrj6z/jARbc5cwjQNC8FemD396ihFfr3Y0Lfj
PlkCeH47ScaPkOHqGicDmxvaLNkhjifcMuNCojqCfIu5M6Gsqelb5+n8t8DXsxNHURFmazmr/MvB
1pkn6Cone3i0/qgkluavDqS+oAQmxLNJc/E42AE9ZY2JNa8hGOdLfvfFl0F6CNXFiftqHDopgMKk
tnV/NbsHRleroIwt8ooKJMS1q6kyCxco9u3duc/n5J5fG32Ei5/hJwapqsY2Z2O6GBBYFecwlO7G
NNdqi4HUU3xAAhjtgvg+5oFg4MK5PJoFl8HFg1vUtp3ihOY7CjDI/GyD6oknPsrZTdQ1Os1RYVGS
fJM4JpjQZV1fqXFMXny9tT+T0wjTiBV5SNj2cXg6tnBKQe20e1gq2CDBA0EDK6sZalOmHn2Y/6eB
lj0X52OhrRN2ioP3Fi/qLd5YALLpsNCEv6kb8JEsEgByycvlEWwZ3I49hmfYgY79krzsOmCE2L33
VQiaTAd/78PT7f4yjywUBcOCb8ek4TsepWcB+lCWlNJPpIk6UIXMOf1pump8Wo0uhQ9USuD9Cogc
riqfkE2uJjPbjMXdvUtizxPvmHrkKFl2Fu+3X7FmC3JiCwlZ+SzMZKarV47esR2G3kqKtlL7KYLw
T39hCegqG3gYkWGsqQeKqMeuFPkXXEzvudvHl2kfCm4D+uQGIZmCVSgNjk/JPXkE0OK29F3kY9mQ
QwmWjXhAwAJMQJcetl96rT6mPmKiUmVSxU1XbaR4FP11nb+y3EgZ0h0QXpLpOkF03MMk2QR5C+tM
WwLclNU906gMylEiZ2hx6azUMvTPBR4nBVl+BAM3Bq8EdpG1yCP3V36s/qH9ewCueDyRic0ZZukm
UADLuiRrX2srTC3wbSQa869qIUviq2Gqg7x8OQmTxBUuhbmLxPcS5/JDDqDsjkHexghtTY1iL1Vc
Zp1ej9mre5pxhZvhvPCZ0+o9BnaxF/63B3scl2iaoLbknx1JxGEst4lC9IF/tizJkaQajr+S65Ji
s3KMZcLi4I25icdgA55AqoCl2XCEXuroIjVbHFrlnhVT+S9RrqZx9akUsWiBvgyhlCoV/gEMymoj
gCCvTemfZQULurXr96BTzCGt5WVLEj62XJRubS0K7RsG5V99QFXRq/cX7hEH6h6wAa+hY+sH9OVv
caG9XIKRnqVCrSSCVKb6gUwUdbDAtdWnahxkKIJR9XILqgQOIPrOZLzzcYg2+nz0eF/+03M+yUjR
hqcf2Vf1SRW/pyBIxxIMXC1GKJFyn75ggwpHyYfLqyiT510y9SCKoT7VX4tY/L06garrVTW97NgU
+zSylhY5Bxz3D6YoV2qjm08SXPpy8BtMh5UpFkwbvE3R7nDifGl95dR8IzY8VVND5xhjHhpAOcA4
YLRtmgqSaHSs1dJX+049AWRs3YlBY0tJ7hbZ/k58QrdhTe7LzgvDLL0Nok/3A7oA6cIpJlkyduY/
8BtJItIh5JcK39TQleiLSH3NNipdDrSt4shNsA5mYX78J6A4vio5HmFGl/X9JSzUEgIsjyGIBC3Q
2KlVoZiVGXM7plWNbAgsctv55xHSQlBr7b1SlRvGMv0pV9g2dxRd2hNgRcVx1AWrHPOTMI+NGMbX
PeJ8o14eL59B2DehusTp9T4QLgFgFm6eOgheZM0FYgng9M18+ujxk44RN99rU1yiZgM7tsh4jG+V
DDJ+8tjbonc1e8dhjh0QgKF+/6BQjt+KEdhgAOrFdHmrA6IO0kf6n96ncTyADf2HLbyGrgjipGYc
P1X0qVhJzraG6Vv+FD/Fy2Fn6xS5RcqMMg6C9JO3OAE0as+7ijeu9PEez6CL1LiFBn7LBVo7xueZ
7Os0CyegQLD94hxPfJDZ90F/H/oH1SmPhhWX5T2aZGP5B5DT+GVC54ewfXTUByejS4atuMa8cZVz
cAdTyFyPdwE/GCD16SDlAuPSkQIeIZi9EjkYJUg4VodcRq55DTvU1FZVMcclQd/jdzWsQqmLs14D
fcYulAN80z8Vz7AzkhFu7hBtRTJqJJg0G7vOtEAOjYvnIUyYf/NDmcc+tsqDm2Canpn5xzPbxHSs
tnq8awMnWSBQlAGoLS96vjuxgBzfCaiJSnEqOrdy4zmqHGHGV6Z43PmTsxSgKApOZkjpn4jXrfkm
diPtkJoH3cRdJUMS0uXTDD3mb6XzhgmLopewsMiJDOEhlIMfk5aKyGMTs51BhelLS/HgL+Hsf4yy
wRCqiANjrYZi+Q5GiFUKETPg2LzotlY473T2PGFWmRKOB+yfyY38ijo+6TZcgQ25O/fLIv4g64n0
GCKBMIGlwVBZNy9tkUv/9UpAJFUZGFSBcUzG/OkxdFpS0BvNpCVptCAJtkTG239PpIHs+zk++E7q
4xyUUWmtzA3OrrwYlgTrF2gLbfBqyU3oIKJY3ptTybNoyk5XQt6FmvO9DBo/l8aDMStu4bFRFqBZ
MKJ0bhhDHxWoN3ODoWgEuhcGidy2YLWFuXzw39ZVGMZySuGFHc2WTnqTnXynitj1q+86zyFN13cb
vBeucpNP0I7nome+55E2JGOnalHzhsgC120fukvHiCot+2qvIzYFSirVE2RoPIYXiZm8eNKVLqIB
SF3pEKMvysNu4ZrdDI1icc/2qb35u+Lc9RfhHzQmGIBQTwigRvRioEeY/N00BY0ghs5VP/pEYCCd
+/ui3oEShzpPz6oAH8ZhfweEl4phusQJMHJ5ryVWhIVwdtuazrkRKQaiE+hsDR2Btm9g0NG2r/Hg
Er+/Nk/vCiv7a4E6Ik+nMNUVxLBgziQ/7NXkzGZndswwFrHId/k+UHeCukYV+SdC2MSSeUNCND0w
mgdPJ3YsDtq5GSldRo02vdTX6w8aiU8/Cc2Pa4MrFlbMYNcZRpfjJXuCTgkdr59X9wuQzLrmEK7P
yT/FM5h2QHeMzEZT4l6E45cLQNlInidtjsYCrE4qxOT5fn+X9xMHHw85tAUirKMeTjuL5WQfFHi3
TH6m5rDvM9C41b7KCC/pN9yrny7tQhjJVZHNXEoGkENVvSrmDqEDRZfyAOP3cpVyYk5u+VQSo1C7
51G9Pl5D62TWB5RFlSXg2HIxa9LMocUVB81GFfdwyyF3w+KLGWRuj6SSnAOgfzqMk14bx9JI021k
pF46km5xVgsomKv+obt2+K93KZNfnnFpyQIBAJrwmR3e2kf9kL5r8HxgVD7XirA2uGNNwSZuTMnV
6atMoYGagnIFYbNladkvNc7Nfh1hEL/dEVfqU1XNhRONYhLOyDcZXgFySN0fX07YsRV6in0R+8ce
BtjXh17oZKqCwlkPSuNcloNvBUHFWJoRDYpZ75VYGDdzvfbXgDgeCFcLRxfn9V7z25+jEiHdLN8r
RS8DVtJzp+IDQLpZjrWHA1iQYYI1geDEeW1dZWdGkAWBra6NcvnMcJVlh+i0lPDn1gELNv3yUTE8
sIYOCp8UAaJuGUPZ6ONlClV/xiNxAALkXILPMGVb9peDdbul/2+PKd6kE5Z5XiI1j8iAz0I37VRO
HesUngF+m2p4LzILx5lzjqej8A35O8nwlIk86NEVhsjsHlSqolzXlH3E/wY67OEMKr30VFbkp2DK
HdZblrqVjemvhUQmX0raMJFO+e3M57cQr7Nafp8wKc9vdFT6L36TFwWNSNtrLQZRXgxCRA/plVjk
JTKMOaJPTdgLxyMZHhqxmbSvAyHPyBqXKSOdag24rbJvKPHmaVFvHA2WnLkwWe3kMnMjY+DkHwRT
MHFdxzB5Q/d6PJQmDgvZaRsejeYyk1cuUdbKB+AQs2SedCznzJ8/IcH2s4P4g+Y8qY11fmzH91zh
OfbCRWq/6L9g3AEhTURmyzuME54FzkF55RzR7QlD84aTj01Ue5+r68wa4BxSJOQRGXDKAY+XgKGn
lDdw7h/vM18hPef5++nvk4MlBpWSfMSkcSKHU66k46Sl7z87M/HQgqn91qhlHebBdnHP9u8nrcq3
Aijr1S/4UEfBhjAPN60PBUytFtBeRMhdyolQITtxi+W8m86Ea8hiWaqc5drL3iD9QWoiBrzvXvHp
VWhx2GsOfKdS/yDUYZtLCSk+hzGG2JtXKpq4FWg4vLj0kS7lD/g9U1MnnCH06BcfSvxaB5/O9UMT
9JrQlSSq5k5vt72eY6ucUACri3DE+jIFp7+a+zv5+EfYhCbLjZgElQ2XYMGghHimLpBsIX4V6avJ
q0t18ajJX/GHqM29tP+DQJdzhHQsvwrjn9BYeyDyXbrVqiXRT3wZkyIxXL1yIJu1EmQEE4e1SLXB
2vO+dX7xCxa7GvyFWq98nXLphgfQ08MQmzT7zmKFX3mj/tHw69649iL5Riis9NFm+sdCOUYaw8Kf
pICNqGzDGBq1MAhj0lEvlpKhkvvNezyKk/6PxEu90UvrT0vPYj8/jTkVlLShwKfsu7xgBtB44784
cW+VaKCzzLf5UZcG94K6hLQOhieHqMeKmT5CA/OT4Sq2vDmksvVb3mMKmIbNyOc3op9gg7Vzi3qg
aoNE01D0ndq8mdsjzVgI9GhdFMhXhSwAX2m2biJDqBcMdJs3nRovnnxYZNJQwDuUjKK1l3J+NGxs
jfLflfB9hXn9/PP+6O6gskhGka0BKGUfTLmW7YK7YI/Gt7Q6DwCiearhrrq23Kg/IUE/9MzcKQ55
2FqrNGrrKtkQQS1tohr43UK0O8m4vi20GafuzK/KFyqs6Y5oaENOPxiZ5COtScNjsBXdxorVM3vC
Hl04F2f3OV46L7D6+cFonliquTMNthh2wveLlVyJ1u4uZDhz/n++Sbu5gb8nAmXwb48bLHmSBHjl
O/QpoqRfzY54Zcbaex5XmYIHwAnbUM/mFs/2X6iHVazYBS22RtrIFnZW4BiW1EB5N9Xs1orEAFKN
1DwCV4AnFDiQ3/OThnx3y/P7HsK/QNuCa6b0/rOkCorfd2tpTGN2qqYcAlQ67uZ3A68S94xxfdf7
6anmzgUum8kQ1lvnWVmiLbwMuG5u80SUlZcoH7t6l6c8kF4ftcmszEEDYBX//riVdaPV4EYLyQfr
Vwb/FC+JkokMeII9tc92M11oGDYnhWh9RmEI+Hm9LEi5FEqVm4ovxfO/lXGzDuXAqua6yREazLTY
hkpqnrm4bVTI/1nJbTrFHz5AhmAEMYnGGIjY6zoBCgq2J1cKQsxLR5K83OHdJ0UYto/ap7vxOzxx
BiW07vV45xwWmysLDY8vzJqg/P268QTJCwZzLlgLZfBhfqTneMtDLTxgJHa23Q1ktFWTF7vrLGMD
AMqHCEdaUeC4RGwt4uD1PZaBFqzsncjmbV4NdfGgig0I2c7r7+hS0MPyOXnb/ne1JZdP7tqzxI1O
iUNqAlyT/XnNWGB+QaE8thDjD0VrDbmkp5XYOv02M9UqdscG/GIeDQ3IIdhCX3sa72HRQay8reLW
iDZUfwCH64sQ05Ts75m+gsjLheBRiP6OQEG2mPoW40tmolulnTAq/HpF4pB/W4scxJQ8iYpW0SCo
u5Av+caTabaiC/WGW0RJcYVywIfaGzTjMpv+gUc3eQGfddN91PAXVCwx6kdUnZUbuGJbSqt/IRzw
kHKMA37xS0MFfQevqJTw18TGiBS56+Ppe6N4cQiFHcTMVjKQJJxYmppsgvaRb+Zs8+vmfUTogvmK
xhterof3A02HINdOQw/kG111uo21ArcPc3Ksi5+80ZHv7zF0HxNqDRRXLAsTu5LUwd/gR2cOX3NF
BgWLDXUwwfUd4pmvTDhS0AR6M0V+BhFkRPkrozgRkJXXKTdnQeUev9pmUZw7I0h7/Q1gYMCRtPyv
obBz0SAj+2z7eGcggLFhH6Ur2e1vIYtTe2SkSVRkyxfsJMMg1HJ1n5DxiI3LVw34Bf3M8S6j3n91
pjkLsZQlTsPr6TO/m4zzgM8dEboxOmzSgEbjTnJTl9LroIDFKQLFO2zRsJrZvnHvrc6BNOukKh4V
n4flG0vDIPoaoz/+003tkxpzd9T9bWiRm/sLaRPr/QRLycE/yrh+L4RDI//UUQc7i7GCcNFYZxND
UG4J3bmKsgR0uu7QGos4AGTMLFg/uThjqso1j05VbvQ8VIexMdfOYerz0qXl+5250f9JXeyq3Huf
yE65soB9RpJfFc9AdPpAIRQOsZ1FYc1mMHhlKUlMJqlSUZJh0pikB/PP127WJizE3aA9EAbl1gEh
PM24EqVDkepLZjurPUSFo6D4asOpEHP5ttjUOHHWASD5yptsM1ReF7hkNVUxQay9b1A87uhFMU0p
zCG014uyPIfSoriuvusc6QLyqOZ94eqtZ5dIqxoWOLmlfq5oIBw6+lCGi0xwEuxIosZty4e+hvIz
6gpDpP4+dV1C7RYT2htwoq3TnvzcptmJSqZ5uX5UlYa+5Cpt0MJ5P6JrwKqRtJpwy8bG9bHh3CJ4
jyUhSV5AmzA5N6XPyNxkFuYLYznGl1X7AiBM2ip2B1S1KgCD1w8nSHHjLsHitSNQnaK+CWy73ZD4
XJWABasY0JriT8ZrgQM5BCatiUemI64o8TDmxxhOwVzcWnboPssapg7Vrq+rnqO5lgg9NpJQA2Gg
qIVOHUyiyKnAKcNNUpon8sqVWwIkGowNFvJ/HYqUbZtqqKQvkju35srkxLN7ukNdMKgXqYWeKIlf
Hg0rQ3rOVFk7FSEfBerPwq1BZXxhTLLzbCOvX85mrqmP9bh91DMPZtndQ/M+4aZBnc1kJeB3EoV/
pOKH/W9dg3lghtTsI4u1YABSGeCdZaNVQ+NdxBNgctxdL5EES/AZf6GEeyoOVDlKlp0AUCptEjDn
KnMTgkKg7EFJyc+PiN3AiY4dJa9C0nKu/wx2Y8xNrK7/FDHEUeW3Gtw+GZsIhZfiipy7r4lt5Udt
suxipnzWhOniS0NRVWifJdFWd0vKy9JbdCGaKxHfXY0NXbMmq4e8MP2wyMdR7sGI3acdK92Y6ouM
CkEKCPHYnr4BVEvdZ6q79ml/gNb3TxCtjmM1uDS3WZGm3y4WV5cDvxRDcLhLAqS4IxLnYK5MocDY
QKF0718yLeKjNzxmj6X/IhyermqhepG50tUIqSo2bL94Hkb0d9uUKYsrHo7IY6TluWl5Ru1ghu8v
/aBorYmrzkYF4qA7QfAaKjN0wgY4VIPKs3MyVmPhqkavv2LaPc+82My/3xhLnrviNn9Jr8IBkT9i
MOJRbHRwJ2epXImmFic236XnX0/0JSMHtndSN5BEyWMuOWAN5jxGjP93OrrEm4QVOTZCcZ28RBHz
NFmsRtL/g4wZwDRhhcwFGW+ovSPHW6WBxhNt3MMvchmDVNs8KNbcz9wxOdiUgEBlOe8iYRHE3PRN
rvyx6VNeRzKBapHJ/vV7Nr464KAtBlVwvGH0/mE7C8dEYSpUp/M97mqx8paXetjwtDcyORxpdpfr
arnDKlfConuQ74b4teeLBj7EeVfycRzuj1vSxZNO+e4pVKKxJedsD7Mbzn5cuY3UlJ8s9eJd/3Yk
CRM5VZYp93TOJ282jHtDxcKmKHoz8txtv1LFvBGANZTGmp1P+OSVnhB0ShuD3R8EmPNdzj5o9N03
Rhgn4SlRc0fxzHGtP8Dr14+jvH9MtRUqSjt1j7J/s/i84Ppm+uPmhWIR9O4/q0zA2i5qk8QKNNOu
EaBtUKaIvPY6g9b0oE/riR4Gi9zwj2RTw7ZPS89nVzwNPb0m6FOHzgsJ+84w/3MmU366IpwRpPMc
rfH2Z4FW4CB9EeU2mFSmbfUdmbnnyrluNDX33JuOkm8y+rp5kBoJIs6uMviVSIB375ZuBMU1D0zj
d89XV4zUf/Mq/bHviiFbdiUUMsXT0fXlmCPki5RUOJKlBQk+lMnGRz06S5h1ZSfdiTP3QWMZHn3r
gVGjELLGCta7S93GQCoi8VW8wYiT3fl55UlHgIHa3W+f1x6o1L5mtNQQTrbQVrhtnz2kCZUOVxCZ
IaiUigYI/gK1HfM9bk73udgNVwiSsE7Tnzi+z9uacE3S3vGRd5r8MtoFSkjPvXTV1+GCTSl5Ply9
Zm87pe8Xb/4pATTz9n2tpIVsMF3mCjJmRdM0n/OKHhfbE2SbmqZnRhKOl3M+enP/ellBdQ1zuM+o
adwu0rrHAHENbYvXI/cLkrcwkk1Y8T+C7afDAETf62ZLJAtDx5ytKxmaeePINdvqHZEqBOMc1mLU
GYrrihJRr5krG/Q1zeCE0arLxdLGhjtnIZKIMN5YUBuLMybTe0XSP1X0HSSlp63SiIDJcwGH71CF
7aE3nvOfqk7YjC3u9Kj+lL0TwpMmKofKm/0HSiy/yYh7rW5fH+Di9R7T5YLvZuJ27fiFU0J8HPwu
FjtXu0hNFPLsMLC4gs8YbufIkcCsuj3Y9PgJQ17ahioxvrFks3uIlvudSh08cIRVC8JcY1rszieB
9DZaV07qr2PnF2kuL3vm6X8fuolkUYizFhUqOcn2XNPSE+Jqb4Jph05Dk5rah3KP0VkZVXza/gDI
7vPui67nh0l+xReGPNF9f4g6zqSTX+Dle8gynqeKscQMN6zNpaDOUo4MXGzsNP4sjTznS0WpCqTV
DvoqxQWL1HiHOMfaWsII1mmzaFtqFKjbgzhttH81hLJ5otKDYE3sKP6/d0i6WwldF1nI3xoPoZtD
U0DDHtGspTP3F4e0bJPoELAYBAiI7gB/B5/Ntp0iOA8+5T9qerFdRr6erthzE/fu1JXby702anaC
bcw4WfQBzb0q4JT4yfo3vcpDHRZTByQOJr/9Z+gaZOcF09Xm4PY6Rcl/Wv/Zzyxb1aRk0jvDEvU/
AdCBtwIKCwd07FErIGciCSLSDO6E8UerRBKLgUgAwI4OsCUtYca+ZEvCwnVf0ihyB8ItK6qUdZ+v
6jn8gGVyLsPvfy3voOU4sC3H/HXIWSHjrM96i8Wm0N7SeeArDyqtYwTP8v21yZm01U3EcLXP/SzA
oexOObunFMqe3q00cIjwpnW5pl9+JOQ3dEf34I4O/nYWo9858iD9coCEvl2kEHyfV6hEpLwH0RDR
+UbVlatfwKnnSnP2LXDAO7xL4VbOanj9mAz0tRqx5H9juZC5d4O83M8q5jX0J7eWuZDY/eS0kdnb
OzjFUTKFgJt2TT8gF37yR/FD1guUjzmHfHkYEN2W2Oa4DHKhkKodCWKFJfbN2QZ1izgRavnFaStx
BshhmB7FT2QWnVi6nOuqZqegWV/8xYjBzROLh1yRxV9vQqvWqrmVCXisbZTGhW1kmkHG39mziddf
H/bzN9l69dvVxdQ9yrCVbmmzZMIrlJJs4T6XujtHtq3JGMNDwgZUUgC44suKyNwPylsqKKBltv6g
Ht+33IxyM/pMldVVcngezM1hcPXV78YRyxVpX177RAu0fJcpxksmdZQfs4jDl5iGPzzHiIb99kNR
+D3UuBrZOs+jncABW24IvRGsb3d6EdPFF3u2yzV5bi98M8AtSrJ/YUq1V1MpxU1Vi9n+7IT4xJe5
rJKCpCpSUambQFAcRCyXJ1FV03ZYeU6B4VV/Y1pE5LMWGSSHZNZmiLwQIKGQziQIAFWN7YyWxuWk
Z3/KQnUOdHWzkz6KendGQOyUmffSBd2193sqBj1nTyvlgPmtp/cWzuqwM6IxnIrE4j/ccl9zm5/2
2cDMVr/jb85nlM6AthjE412hmmuaCihDXH+6Lv/adej2/hpyM0rMTaQgcEN83/zooRTYMNnfpIz1
lbFIlJb+YB0JQ3cNGe5/rsnoUCXXugp99IEso7/BiVU3x4hi7a0mf0qr4ryVW3pyw7ZSf+wCW5sl
MHnJYrJfaCgx+VDmq6F96vA9KSJsOKoqGwJyp4ToTo27OSt1j0Ziggrm60o2HbhseOzU1Kf5+KaF
65dIbHAjPrKSxYlPdjxEfRy6EddA9PdmUsy115NskjUz51SY/AsQD/HoOmGIsZaBIgcFEnvlAlkB
aKwVnsnp8yZbWF5DZnHNZz0JV2F4PwzvjCMtI2pLmO9GnMxLCKsSzdsHVyA/2i/cDr/V0+VLKxyt
AeKz4/BprTQpQJX6M+F9qVeMgvzGdw06bqPngE6+Z1sy5X38oHl1wVsoDwGn5mGDov9/HcM0SS89
bzC1dLYqrHKb9T19B/irlUlaYe1WbGgIKGHNXdbf8J6gyi81O98GQM4z96pOXDyEmmKevAsoPBY+
LzBprnx99lnx+cQSsoyJ4lE686Ci+BWiuMIurg3MBdXuXCSTaT/IZgxsx7+OeO4o5SzWoZXInnfQ
h9MMKCc02YoIeYN1rY5qFJ4M0eSstEOQSdxVplIRFRxyUJOgeh/3qaiCbWgoFoxg5R6jbhIx4zlR
LNEzWT8+8wNRmSeaEhgrUXAffk77SszUDxgqH7P4r/C2g3RmMAELdrL4qFs98diOQ0xO8Hq6yimu
zukH3OUlot6/58cU7dyNc9+F6gTIvXkMzOqYOp2gfwOLX7jwlQEuuxkYYbPTawD6YFYep9FqSWG5
QIFKuADGhyTAKLHyVj4CwmehtKreKt8RtLMhlpfkBXBMgq8ydylCJufqgkJ4NiJGpTollyOIHQr4
1boVWpemPYin6n25IH1yBiDLL6JVbc+DgEuR0noJ4JGEIdGXChuaKSs+3SM+TpAAaIxW+89zgogr
7zQWy5vASbprb73XsAZaGdWObcNePPPaxNV2NBz1lglO1LOLPxOJNNE/oLU9qN/IIAywg0WcaHVe
1Zljb4WdvgmCTRPRqVk5LEM7P2TRtd65rWF/oEksKS+tFHoetuv1u4Sy37xl1w4JgSqfr+yxpos5
fgSTH4+3exkcSFG/DwEpnZ+P//XBueFpssbwdpN6HPGc6efidDozxtNicPU16GapqVZIUPNtGAY1
khTFF3peyvihnkJg/yXfinXK70QSUYWZ2us6Bo12XVLwicejH9Unq3V2eKRY2HzGVFG4L8qaO7WC
mS8TgjbJScK7hnT8xLfZ02g695eGCJPfsrFBcUz0vKjgkcVvM7jwVya3ServUQFnlS+NkKEl4t1D
pJA8RgHcdRNVK2eFO0w6HRgHuT9bIADboXS6vE8VP+0C9S2Lnl6RtUeMstBzrFoLRgj6jibeDqks
Rpxo7v8r4ByACZrMYBOuUH70Ba/bbiS6idjTbw/LKmd+8hSQCtHgYJIfDpnkFG3KvYjhMO3ttMMJ
GSo1fi5++B8B3cejimYp3tegwc80H1tqy5OhiKB236YfPX7W05e9AYJKpgbCPOEmItgbUv+epfTu
a0s2FTdqT6XDLH+8YGNLMWZ9YRopMKhOQIlfxEKeLQbeuEG7UTgSo6GCmDinHlDR0p879lkx2i57
KUZVqDbAsiw+EUNTRVKAvxdmqHF50NZWli8hUgcPngOWKnUs8bxtj0EZdGpFC6jNEnnIJ+dr/rRA
DT47zrL69azmpIUIMZPvVJFbgyWuqGJkXTvodEBXvjQvO8ZBC9qzaR+oonzRBksziCCw4Is3INxO
R5mMu5hpZs+DaTZSwHzNb0xcNSFXP7R/029zjL5ONZO0n81SAAPBq9eIW5w/DacfFxJ9/XTr6YOY
BB+QqVo/wQpVSfe5GIU7YVay+O9+W13D+ddp5tqy2n0/WDAPtt7MOqzsJu0bjqLg+r22UJy9385a
tLooNLi9mhpkECPw958z9ZLXjIL2r+l8NrpzkFlOIJqRYyOkYLQwMutJn5AVTMDW5a/jG96fUxjt
Toess+/bjs0b80oC/mjoHLDmiv0ANnNT8MP2i8yYwPtMiWvZKsUIQDjrUtMDPm7+yW7i32L9oNYG
qSrQ+IqUe6WtoIkiBybAjhG9imnSrF4w8+XXDxhLSCAm76vqpNMuqX83arsFxdSwRIKjbyZL+D6m
/S3lpz4gLkMrD2KUvt6OSyD0x92HCm3WnTlNIAeqW4Q0cd/eG9ZnZqld0dpDIpojD21pUDBbntY1
y91powkWBGP0kSrFUOIT+gs0zPw/bUJsz6S2VagauwyrQK/i9yd8k7B12xS6cAS4dBYateAaPFUq
HWqxrlR7hlX+vpk9Chb7z5BPSgm4d8A+ReQNHquvx5hwlaKl81oEBSo5tz30DCaAIz4nBUYY2Uij
UiANTdilnHmOEw6+hlDYuqiRB6z+aciEUDPsFGC+/AqGuQuMZEyQ6lM9peQDx31KeT8c6iXF3vVF
Ys3Ru7JIDbvTOc3gEwAfrD1cYCVvN7Q0Rv9H4giR/ITWpfRCFAsMw6mY+s+HUcUVvjj1eQKbv3sP
99D9aS9Aeq5HRewC2G/PhlDBS028J6GlTStBNrpOTeUApbts+miR405gSozLCz4e1xQTNLteca8z
B4FsHMAUUH9V/FVJR8AXX7rIAIF9RXCD65rMrHFIONubvZtb82yjL84/DdyCYTcnfwP4wtexRiOs
A/Tcf6aPCsvLO7cR7nvPEwUhHKIoXNCCKbdRz+ujqCSPel5FNH8qKN6himSzWxfaRGHfWfIJ2Sxb
lJPBAOLMi3YlDRjudBIkmuyuLsqhCcjsc2u6BRjv9qFoqQHghCSFjsD0luHyxfZf9SfemfJD8d1s
OaLyxQfAzRO9SlEO1MfSF1Rd0VmZ+xLbd/PGHEd/dFCLnmhX9jKpearh9sV2PMr4krqdj4bUdpk4
cTfob7Uk2sRZtjmVgvOTfgj4v7v87YoV6zcrDQy3DeZoHBBotqOVpWiXbrFq0w7iwsVsNPzJxZnc
9G/O63CMjDNKTMnr+wy66SYYgMdzReq8Lij4VMCoVy8DPBbGw7yTPHFKgwTg5VbgF9ICUF5oJKlc
pvf8920Z2allwT//dzxJhn/sgVfnAK0bMXHPtgjiDLBCcPkoBUBXewa/EOfxEcZeUf3S7d9X4Phb
z3CO5f2LfiPcLZmTNOrh+bjyHDPN9Zs+1+KuhdKkJ5jwdvZ0TlnoWaZPXF3udaYEkv63f2mtEdAl
W4oyIZtzVTmnfy09lEkh8aUx9bL77mrx1IgwqoOsR81WMqTy7k53hn4SID/g/L5IOd2iRIOWRhaL
qoZDNwFmvaC7zvYAadgi0AHNLMZS4rTj+DSqHGXiwhzT7Wkq4qA5hmRR6JBy/cefQKrSNN4kya/J
OTMcM11McXnq2Yo1nNITSWhflHtQ6UR4kROGe47KcInTC8P9mutX+ipzdBPzjZOGT6Ng95TAHVsW
wUhneJZ3hZyNuoidUDjfNlCEZBFBmtm2fmj41/OzBXJAjHuUd4O0W8QV3idtZH5OzEFFpQ4PDivQ
LbuX7/Dn6GgcbWwa5vn88nbxlkVkmi7moTOkrZA/V9cGr77pUuzDrKY2IzJoxwp/3rrqSm5UqxP8
U/DMPiMwqSZyMZxYNIvMcXoFGsncH/HC1PMxhZw44u0ekqsQCLA53uai9ESmpXHHMR39RC1GzSsH
eHolYVOQreb6mSfebdVNfnlFg5TNE9raR37vnd6b18iMOjxx/cgxOD4AzeMjLQs7XjNiF7lDwdRD
c5SUhkUzkeoyMkJr1oWCw4Pdro6q4Mx3Pz3k94SRjx13Cw1Q5MmHM4gFJNN171oVqn4/+WreVX3D
rNdTI7bXdljfS3BFr7lM0ORJwvYewAeMw+1nKO/ItOSQ1FSEoCpfPPYXvxwKleznCWTna3CO96XV
yau6hD76U1xWd08uCqioe99AcEnADKR/O7J89k6qU6NKPKM+gGSYrUBF9I2vdRY3Nr+wdserbkZS
4R6usSHg+FF0/uP7K9kIk3RemZzI+VpFXK+x1zCXMXfEC4ghJWFZ4uOk2YOaTiNbdycTGJ6mH05X
l6vAHXqWbK8zHBX288ruD3fT0x1tbqOzsaoy110rZ5prjEipMqZEs+zITFGuBt/rflmW8YXZAaGq
v1ecvGXKBgZiVnmTiNto1cCBFtZlPkF2Wv+08sC1GgauhQds3mt+OkQPNol4tWVkvbEGIuOoideU
iZDY0EzO6raevtiOWtrQDWah6GTt2BZLLZsBTHoYy1WJnuCkH1DukaGFXkjzK5I3MJjwGNR/Zg5V
F74IF+qlNnB6Wo4hGnDb4J/YJq4JGlpoC2Zwx3UvafpmPUgFjLo1C5yYrdVLcFKFIlpBC3W0eXxn
z3C1cBXcxjTj/rE0tNf1BZj67lDx0kyE4l6VTMEk3hfBRn16WriBcG6KNVdFN0shDwVSI+THXggU
viYEaABGg/fjjL0r0c3qfkkufkIEaWyezNhYDGVcohtIDYzLSfJywBN5hFc4zm8OTgDxMJ8Jfv7w
KwNAbaaRIxBU24uT0Xb/oO7uCmMKyr6Lo3/614WWq77WVUSJ/bhYW9AdRZfuOPLHbF8hQJ3jGwqD
oS70ebmv2/1/Np0lB7ehVmZgg5yWBywC7ADxjjE+UUoBT7IzLJKY3p+0eH1GJP3y/bUXTxAYpkxi
nJowr26xBczMETzELRr1OH4fnxZzBA3OQXHfENa0O9wCXdE2/mG1Swdf0/fuutouDlABlJZXdh/n
wHVQsMHci1/NyuTGqqa/eljT3tWWXVy4u0xzfcf2SECTzZ1qmJTbjmdsQhC8KVsDBeueFLSWWJWg
nr0dr9ZS2ZfRFHTjRi3MtNZT7g+tiwSulHVFmGQADhKtJ3xYXQ1avmVoDBk7kxNBiBu6C+QnT9Vp
qcCY1zFkqY4Lyk3EKrKCYTE2MAKCY5o8bhjsxNrauXoS+NAp3BqfsTd6l7+baZdM5r/88ih/sxPG
H8TihlzDVnXatuzzWMYLCLEt0D0agsxgkcC+MzmRbU5ZWlujTWdL1yCtPKBbDS1e28hlrNUGV/Re
lsjLeE7zs8H2PJgjYtWLjgyiSe2ohaX0sef/uNf5yTVte08aGQaCfgVgWQYTJTCPPuUT9TPQaFVu
FQGXcjSN9s8PrEPUtI1LRH9vMtLnNSGa2jyV/sho64yPWd4A3u3oTDgE1FwXBBGjTjaJvcSWByGz
kUil9cU5P0Wl1rJqMdOyZTBuLhbnkRgKWNp0+ikZy3OSpFRs76bTJOuKbf+GSpGvrjAbYpXqFA6c
hY6f6J2xfaPFG5d7CByky4ql3UOuHWVEYSrbJSbP7oQrwfdwE3VpgzkJo+23aZFfDCeYcvCexg7G
uv1dK8EwmUXOAUvRBGnMaWYnxxARb5sH7iBCKl5/1eiNVLlmFDMxJT7VdstAMcZ1k54HjX4iQReZ
AN49CGVRXLqzxqaM0fA53qe/PWv5P/JEQodgw59ZClGCI73QXpxYwVqLeTy7ucCg9rYzJeWgQTCn
nhhD0uknsrGK0pB6dypf+hYnisWu+xBH/W7U9YEeyo2Rtpd/vL/Jjm7qQnxqPf952VG1SMzlUsIY
qtR3eE2Vrw793xwQJx5ULi+R/SyF0kkf30H+lLs2G5fXyIcUrIcfx/zS0mvp8/0stekIZMSresAS
hPnJahDCWRTpArL4wVkEdzU+HTll7X9VQmgSJSEXd3Wk7aw7ZBygBDWUwp2cgY9dfbkfv8bEBNY6
UmwczuQOsWMbOqqXUPJdTbF7DMO+Ct/uiDdsmGTRY/04GBhITnuuvs2eSBG6bC9JNTq8ffbIaO/t
hVsGPOMBG+qxyTNMpCOs0bXafwMIhD5sndQdaRozWoWAEc+nCrxkvuvg0fkFciTbFYdPJvn9+X6Y
PcViB9B4W15POpTR89t0aKKMcXU63L2YifsK5d54PGIwByowxBDR++axqsQ/jlD4myoKt3aYFiGS
TRCV49FcGHioeOUDPIWk1qrdB2b++xi9qxTZe1GRkF+yo+A7i8pNgPtrLHikb+plRY+pYH9X/B81
uNd9u9U8mNzPhRTBZbAorN09zNMLpjdptfa1FjSDivOn4MAgOithCycdjkAwNR5C15GYVtDITkzK
ebtNAYLU35O6S/8/A9X8UE/k98TwwifQCDOG5wyAIf+QVzi8y4hwoBXrHnNxm2LShh6HaUh+5jcj
ybX87R0PQmB5D9gy08xW7WFgnSbaTH35MrYHHFh7tOdE+BmGnTdCjUErnuPrOcoScDlYLkbzrdQq
+cYsrFIxroCvXDq0fsY2Tmp0DBSv7mIrkisJuO1ZrVRQN9ZQjrn7Fna/Q+Cyb1ra0YeaKSfZZSsz
Q6sUMFLHQ3VQ8+PQWBxIrXQV6p12EKiKidSAfTrxXCZPb9qhppBuOslUsuJUkxWJcIvQAv2xPvgK
05jP8tPajEqvE9A2rBVpQ1fPkk9/jQwv+W1pqNNZt+Nw32apxRNyhPoPjijdYhceJnBpu/aZ4Z5s
P2lLzgZgOlnS7BAvzteaIGpqxDC6g93P/Umv3ZosnaSzixK67yjAPWQ7UaTqk///Cibo6qEkwPiy
tmZcbz+/KxIUSFmeXKPTm/h0s6xTPu1z/lodQmdF6c5aFbm8cqNYD3ZHnO9izNK5+4RA3jB1y+R5
1RltxZp10jcYln66YBJm/XfOb0/xKiA1DK/06r4v7KUrDreKhrp0+mwxBKlz1gJRolBCeLYnJmzm
bc0yScKGcge7Ojh1VwKi1qcsqopKsxhxLnxzhxTBlnR5ZUasrLc4WLrYV3cGGqIoqp0tph99pdTw
/RIUv32VzJOfuiKheS3wsE6tvUZsZdvEHsaej301DSAU37+naM7tSQ6ya8ViXGA8Bi95z6mgeXlB
it+dwnHCTF/HOvjyJ1D10qnnrnG7neu6zZ9B9Zc6L7y+OdTOzX1GvaTurdCwdyntpqlWQF0xRZO0
xDfc8kBWIXkieiax4BWaNaOjDCkfcMY6fHZ2Hvaxc0Wi8gX3mkasaBLTBRdKbHXBPqvcCSR9W/cG
esIAAF8ZPlWYpHwqByuJs1BAq4J1N0HbKfl/RjSIeXujqcB2jhBmdsUP6ydIcPUCp8BTXDvIUyPo
ocwk+QUakF+TfoSvW+TPWpqQMglQE6IpEMzXK/ySNbeh/K/x4/31EZKSM8Nv/4sjIXLo/mxA6QSt
Goy+JUzRSgGzBMpOOCEnKR7NdfJdaywNn58NXa7Eec8IXB/tazHv+MWA1s3aFarK0KdK1jg73VZa
uH1hT/ujveHOhb4gujANaDqjISgLBGtnpGEE4VFTSvGI2ntrAViREhGimt+m+D4G4xy9c2Zdtiv/
iUag1LV9xUYSa9wvTG+08Y3ii2caizlrnisfXtPr96FCQpgDv9FvoraXhstrUgXsBmKmMwYTkVR5
f8+Tgpotvwkl8wqm51a2VaAn2LgBI1yqCxoZ6PJLbRKzYvip6PPjJlnwSHHDvdJKnZu/uhqeF12N
Ap/1m8M2qS/SaFmxsNQqbZoTxbM5dV/JBfa7b3TN3L5sV18cW54DlmDVl+qEL3bBF/mNGIK0yRRr
AwViHg6aro+w0fONG8Z2oNm35tmR3dQGDfGdDOPY0d51bD/hjrIcRgzwSmup01nnF2g2JBfKV8Pl
J6Szl0wSwnNcPycqekshwyRhf00fuG7pnA1mHH+ydJr5m1WCr0Kixz7lL1pbQQVABY8O7MHL6gNC
15dPENymhQmA2d6+hEvIcRnvUb0LTvwoxcJ6pEmk+qAp3c5+mNLutyGbZQX0WI63nxLJO1NHiaq1
TF6b5XcTi1k31xhUcyCAl42BA31K7SB0fVxqarhEGic8t2O67jtrh41FnjLB3/JfhJQ7NQbgaoaB
JaziGDvffEit7jgGhdLSQdIJUEpuSB4FDUsGSKAPnNmoObtMYpM0h4s9pNXKWY/enLqsm38DA8uy
c65KhVQsRLqc98XjGWtVVMNVecnO5UHX06pd/OFN5JHXCzobITRCCnXpOvCOB6xBgH6L+umFK60u
LkFnX84Q6IMbxFDdVI5w/6Xflko54oIFFpV1QwpZzrYtpKNUx6eLtU1S6bp2xqdaZYGTmJMB6z6F
dDzwTKwSQ8cosw0DVWHkH3eLXvLAwPK9rwIXjv015pw8M3Gnx8DMBH29Y12fos7VZEsloymWI69N
TYSgKq+deEcyEHoVgSEmPKuFxBmkidmEkSGWTT3LAuoGO6t1Y1Xb0wfZ+BRpVPRjhhQQkBGfz5b6
YwwcyL5SYJHyZMqjPLOVns4cW1k42wyNmCR2YPuIflkFr7p9W7LaNBaZmXXuUpilzBTWZmLX4dmA
cZPn5xpPaU8BfFLxWpyv1ZpvR1X/WSgXKHkkzl3SDLZpzARUSLFAUbji4JSP8zgB+d+du3RiNdWZ
hXHZKPSqiZjgoyyzlVzYtaVP+Mk1u2D9FcOqk0V2H7UlGz3+dDFQZenm0E5kFHmiNgy41MYbZrju
rbJomFdklOAYSNm1M8FZQlQRQ+mKU6R3sr0mrtpbQu/QXBnSS6omJG3GHEHWtsoSMUJezJ26ccHD
PEQtjg4XRaPX8pysYzJf+YU5Y1g/wcz/NZGuK9L6tzzX65NBk0GSvj+zAoZZWqtkg5OrxcWy+ZA5
ZYa8p2WQOudnLrxI3fvmATAeTi+e9l8a2KL2WxHIX95s9YOBRmysSNn/p7l73fMb9mEfd77d/Jpb
3eqQ0Idig0hml8oY+8Y1HhRRSWmn5GE+qTSna/1ahuO3IAxRuKzP2hfs2x+mqUnWEnQY8TDqdExs
8YfKdptn1nRqf0fR0s8V3i2awaKqTndK+wnA8iUnq3NlAFnbzbMH9gmm1mwICgzGEKtNPYcJFHkn
vXIGveubSOL2kTybs7JI7wLDKH7mTh1KRIL6Z0WULgpnOKMcP8XneZKXuv9MkSZXT5RkoF3HHCyK
bC4+Pcd8crteuaAr8FHV0QKgknd4hI6EDTN1l3eDWq1FXRpKuMqKGyx0OG5LThk3qEiUfMxv+wpL
tq5Dm5OnKRxb179f5HJ5H+Nu5G3yhQG59UTB2cz7SPqmAH7NfJqd8+LZU2OO61WxOPh2q9rQilE7
/1mlyAbedjyBQvdSC/Rt5X3husjBlluhIjFmZwJaV5Lcp6F9tLvN3JbZROVbQ4EmrElbIqKRtscf
wiq6r3La5RMJE40wwrq/pAwA5j+XNGvH93al9CNiX4u08d/P8k7OkMHfH68JIk8RqNVYCYyeVmCu
4octWqGY6Y4INiYpTAdix9fM5U88ZL/8W4biVLJRxCWbqoaGUJycerJt53+U6Z3JSkyG8MPwKrwj
+A8ES4B10kic6rBvESOM4WeWXXcexGR/rXpgFQsc6pA+eW7NjJMxaNOeU1nSu+FR35HQnSD+Uszd
Mfu6F1hIEFub52o3SuiOIm6uhWgDujGl+wWDtFXbmgQCrSm8DKZGCjW8tTcyruD2fOiRe+EI8REY
EiBhHohnccZ02tTqUgeOh/Rrhb8PugCOxixzsaw8JcObpo7KKiqRR9hlcC+Zs7NtD0Kqwj8bS+z+
MXOl/B9OsMixGFKlJVyLtiiagnNfSlYOSREOE/b6aWfXf6z0uCq9/LAopGjLQcd4wGNU4Kb3F5P2
ux/eXmGnEh4qESExsFVveNqzABEhgFIz0ibD4Lk8VuhGg8bJ6DoSMuz9XeEib43XCrVrNcMIxN7E
tFFTvEQtbJwHz0vnF1LUcgK8iqEkcPjC8ilva1cApEMk7deiJMOMTxDfGYVVi+N9em0JSUNgukef
oKtOrO9XNRKQ4CZg3nLlhJp4597dbdFltLE96jrZkpCZuAci2pd9WLDjTVaLvhiSuijDzTOuct2V
ZNiHggjFvhxrG2k1ySQhMtOWw9A3s3I4gEdX2Mx75cm+XPW03mzJ++zfPPi18OPnHQxkm6kXcPUS
cwgf+JFEKe2v5nn6kzgLawzhiUyKC5Rc6c4NpsNDRv0lgCovMECKLZgr1HkTWmqI3CSN4/sT+/Fh
85iehe495vAl6ws+CjyNUapaqcgjJe6OQmCG+oqAp+ZHEyRGqpQ2gZ2FBD6JZz6G1JhNMmMEpl2S
3A1qrcvDWxhkFL3QnljqS6hHOYhU48kfvhhjfDTGJXx8qgWdncjvUIsU5G6Wa4yORSTI+vBW5064
iCjL5twvXxJopRt+OO+IffasiAbicCfS0qDDtbQgFoMN/YnCuqf0yppinqitvvpqDyOKOjqNL+ig
JOLjamrllsWRFN8UuLlnH6MEQx33o86yBKTOmvUj6fGEoGA1XDmBZEBqhzwqzjr7FI4GD8xuxS2H
mSQW0VgYD9seB9/8AprKLAyxlhs6Y3jQtJz81rUb9LoJ0cjIDinbzyuAdGMW10imA05H0U/C4sw1
YDGG3Vm72gP7UJqCqA2qR4imLJy1yTCy33vShMNeXSqbhCXB8DqC+HxP+/+5BhihHmEC0gFdcVQ0
vOmlVZc8UVglo4QOzn6Qxj4Du8Hr8ZFc/tFcPFVb9qsyJ1NHjVbvS5IGFLx/M0QNZ47/MdyY12Co
MZWyGTWlixc1LIBGUK0gHEQWnwgViJfpMcLp7DroQ3ZT2xzM5FciLojsKrcUDEfZ7WZxexQkJ7uX
gKs9RoGiEa+KAXYeL0qKudV7R0bo3U6ECSN2E0bzmkeEL2qMoy3KMQ79kDkTH9AZyZb48Yxvq9Pg
6TNBfHALMolRWkF1XUYcpED+uOIhWAmjw7EbgBhzPvl3dHWedNKq4KZW0upGgqRSJO23uiJC+xW3
nmsktIUioWHDGmUieG1y4ekMZA7K2MZweW/JY/RUfJ/SuLWaiuFsWJCOm0vWMKE330pt91bQ8B9w
PiZP5oKGh6TGFHTu8NYNdA1yTBDX42fKE7bFjB5s/Z7G1HxDKSBbezwTvXOrV/sfbi5p8+YtRbgJ
1MH7yyLMnt6q0zWSwU+36ENAIfV0EtbtK166GAUv2J2oo5bpMqiRYbw2g6i/SvsjoZYmpaLZNU6u
aCLPIM01r4GYMeDFXAuP0nFaDYvuvRk0pjGdDph4Tk6c7PMyi4Ik0zSvecjgvAj0WmVwpTUnFMML
+5w/qaM1uKoD9acqTb0h/W4sixaNwHFw7QGYkS8mi/xgq2dLlq/P/K+B5Eyv3m9rHtyoCbEHVYvq
pk/FReFc5Pxt2SPLCbJNK7PEwP83/SFvU8o8jy+04qwzZRsKAX3WgfOTldFicXIT6Jbhi+6eqs7G
auSd2CqS+UNXTqQEqGQJjxw+7Jo9ZHoyPgPMl4yol6mnnRuULuhhRKcgQqisjcmlt2tZ5iBUIhYg
KWviYsUogw9mk+1iEHbZt5B6TzyVp66yPOFJv0fQSyKk0Db8sV20P5UFxKbQgfZWM4utlASMJZSf
xEhCpH1pcCDXnwgQYV1GMtl5LpusEVrWYDymC0G5ADKh3CiYyD34gBrI+9rcdfvM5ApnKDVzuycW
EB3rb5BXRt212R4A0sDr8Pkxf3GEkZjHyriw5bS6TRPkCbPeV5KvymUZ0Mfvs4KtXBlEpM9v0oMc
u36nejlgOHGi1nvpJFSOjVvAbuK7UzlhawS67N8f2UN9kYxAJ5GiX8p3ASKDRHw/U/ycXagKXHj/
Q7FjT3chlBepxv7M1Dpt+bgqOqDTJqRgqtvSnnxOoS0bajsOpHENgrq2cOCStHzoWFyofj7lZrOj
g4TGJKtxXJWvQmjZWkb/yzDpH8OPCib9fL6y9mA6vXUG77abcyH8kgBApSHFwnrWNO+n/Fxw/Xc2
Tqv+NRd2mD1ZVbywGrB3selju2Z6iz95Gd6Ezs+GTG1BIcKXQi6vMpdbHbdTaS7Fey+jPIKGShJ7
Vsk1eKxSamq/2wEe41GgUgOsMHLcfZTP1lY7ofSQ/PHCVL5WM05hJWm9Bgy87K11gF2S/acaP9JU
MkXr5J9kkVE2LVXfCmDQTlfSDmZSjiN0l6ylBWTRqpRF0nFVSfnqBVLo791TTahRRW6LIzjtMtHQ
wuuISQJgRe4h2b6ZNY+ar/4hsUud12cIyPQaLpsk2aYACgLKO7XkvxjeGU/nKKmeC8fuuvhnYWDM
ON3yZpgf3veUWAl78cc9sxfdoylJCxwpV2jYuQwPWyoBDg2BfaGN0EErqqgB7PUyj1j70ug9V4OS
MB5ddG7mqIc+t5RnXNEa1+GIpG4Lki0dRumwvm4Q7Fd42jzrmV1R1kBcr5j/ynGydZiXgQru3uM5
7Sw7cIbj34iduemJcDyBPmK97PE2V5P0k6L0MHZB4MSz26E5g+9ZiJTe85Pinkhu2/e2q+A/j4jN
MG8O3SLfHInuUfjiFze+aT0FpeYoaIrMrsCTEsdOGUOhwaEcSsWVbDKVupZLkyk78EwC3IWYoS3L
QFIoTo5oqSQw163xTtdNmyjB+yRcyCUBDh2xS90IDZLSEeQnttCyaroItB1rkyv9tGwUt57yg+uK
oMfiU7XEk8pYztfmTA9ZIlW5w9/bc72ZFHENlDkWCwH1LHY8HrQGJJODAt00TiF3KPDs4vRvOWIo
lC37wZLHqPKOnZppeMFOGXgIEWo2Bpd2piPLIwwr2C/x7WfoOyt/IOdatKJiR6SuDENn4NGFYjSd
HADtq0b/d4q40ndEIV0e8tDoHRncaKROJX7ZQ+4hxF9rtChMmQqq3wk6Qjuy4GQcGtd/gdxYKoc7
zrEh2GhFLFO4t5Biw7xtPJmfVO/EViJO+eT6lgRiwgfR3njjBZk+2GQz46GrVosIGeFn2zO/ER9P
SwNb0WNCzEJT17m6eLlRHo/+268Q046mf14YlWU7lSKUCzcystKXxwUjPqPRRTKfbGl1QXalvoTu
4Tds5VRh1twzCU2i8yRU45Oo3g1GUpem2tioSPrFGttCJlTpQTqHAgx9cDfIHbmX6SBFwyqctrSM
wvWLy1vLUhV5RpMsGwZqKt19IKhcXHyUkFe6RsKQJPG6RZi/uDDdwYvGub4cmk7CUMt3d9SPuuh5
6xu5XYz/HVe+LGG8JPCGRTz1TFFgWeBZW4Z98IPh6IukWUxfG3ajLF3RtDAbN8pPYLsnGqLBEUee
KLDxoGTvxHFVBpf9bkQZ/bkHzlZiDAk35+a8GDi3Z2RyHj7OSDDI7aZzO04Q8Ck/DyROvlZQKeri
P6jcsIqQRB2CmhfaKLW+ULb+txhi4qmDV93CQGOoe8qtnlypWSiVxARXDChliAbQN8eGfAFNnvkG
JnMaCQphrBZ1ugKJwIUZ+NXlaqQn2ZuCdWy4oMU7OlgL5sLFRSToeWgujAB0ykprZ0eNExokzi0y
xn8BK5qm2eGIzkzUqtJn71YDteonis8d3oezrlozzcZn2oPJIBhsc+uGDpgTCJUMt4zdXOHY3LbL
u4TFx476+ao6Fb69P+Lf1RSsmkvjoL7gUjn/eAmZZ91o8EQbnG7Z2UM8CxElSfn/d7vUqtbj6SS/
cuFZ8zfgg9KXaSjqS79yyyMttcq6/Nikw8x38vFpKhePFk9rVFIgeQGipnqXCf2fOTSKzvUG4riO
yJ6q5KNNHVqT7bKR9U8Yf9PI0HGxelZDdClUqUZulB43zbUBYWzv5qLHXj8c9c5eVtGZ36HLcxyi
OcgxU95ZVVo4mOSKTR/VpPpiljR0iegVfj9JOLwwMkhlOG+dQhf4WhWrwYaVT/cp1MY78OH70bYx
73RE5HQLWgLXZpV+7S8XpzK042+2XmhD68v90xEPjJs42dSE5FfADIVrFT9zjf9JWd8bxy0SrZdJ
aqgNJfXgjWPCO3wUtf6djFqSyjvLO0zFE1ucnJQCjbTgEQFplbaSi8et33z6zu8YyhUYrzfeZTiG
wlBRq9pxFFTbUdb4Py5DUkUTuXXE+uxkzaQBQMYDW4R8qrac0ti9yQLxTWEEmvxy9eDQSM7FWOuL
vGEItWr1RPQ+t4eHPrXE7k1sYgdvXVWrLwmCzSxkBxPZ2Dp+bVigglE+mToHhtaWqvgPjjv10+P7
m9Lhc8H+SGSH/FhW31PNU5B2PPksJmDBKQhkTkzUdR2clhwUpsMgkmpW6ZYSRx85MDAobFw8xk/7
DKdcAHR6ZDVJXaGpw7A9/f8czoZw729TvsFw18tUPs3OieKQR+6hy3UMAEfWJUhCxTD76nZk9v9w
55jfzQaED3oBWR8v6NdVLtaxMpdqlloAhXoqqIa7c7YC5S9SEzOZTZ1SX2TgU5hCtTVLzxcJwzqP
CkYlcbvtw4AP6j/Ks/YKUJ8mOKleiH75fC+JtMJ/IBuuiwS7qhHSypS9eRJtNGIJv4lQTyGltg3U
VFqzVPbSS1X0oNK1+UL7acks+PRfPrTJT7H6cvSrUry0TGr5zEK1W2Vie8YIhsA21UfhkMzHwVQl
RLIWeqaK8nW91h1RFRIlx4swqJuZF4fzp7u88dWiqz8Tjc0Z0jxYjVYlo59+PYqLhLhKVsuWuGs6
+xTAlAweh8B2qq1lT2zvQ0oIA/u8v/+jyjvKi4BuuUmfodjAW1yKyU6q79jr64gESLaOfZNF2I88
9F7qYxPrtMTk2zpWkc/g/m5GSC5T+SwwJawfOLp7Uw3iRo0+egxYXro2WQj5U5eOPTpA5Hy5xSJu
mdBP+fxHID0BuIHeW4p7T5Coyc1WD7qkFcmfx/G3uNa43fWP31cDEyIzPeLZ379caycfaRin/zqk
mWaDRPI8qj7pTQRHBFTSCserckwNHBoF3pwIBi79pyRu6vi07Amv9yHOgzIHBEW3+FcfHNRYrKzn
QUqTwv1GUMooEOUihdWIlc84MF4neMkjt/C8jtn7+1FXTIyjHNm70Vi52TmFV3aXByiZAZuNRGxR
5wPEZPdIq9q5HWtM3mFB54MrSzsaNYHJFo/mHSuWfKfsYctPzvvBN7QPmTMTooKGxo9PmAIcg4zq
IiV7h+LFoh/HyGJTwkZ3R25UEzzr51yHM2S1cWZCwAY4JPD2BHBTXei0xBdWDzj33zJNNGAmga22
+t9K/ftPUSFNyNI42SMzqrlSgpeoJhq3E8xQbK6Jsk8yMEP3MY0VgkJR3qkKdl9Ud4DGa55D3B16
C+Mtt7lezLLznqmGQ8qQB3oaO+p3FjZpjj5jD/L0hthTEuKo0OmTjaqOhOHAPVnhWzTMg/YFOJD9
PhGgZy5XZ8S6EsL2eWD/AmJoZGCSWssIT7DAGiJ6WBIaD7EiKC/O01FpM3nT42bIhBZbBiKBPX2b
ndnysX7Lvr8smqipcybsApXCM6Jw0aWAWYHMcPZOD85H0WXHo0sWLqh3e6NL1u1OECfxBnTJGI2N
Th7OUK82DuG7Fb4Vfo3czamcCSF8OzNs+YlRoTPzZH5TG+siSz6aP2+FUUiFa5ytXuOaO28ywdQW
frHLDgfHfpLMKX7JG9jcOnSH/M4jnxTUls4G/23VsCNzXdqNTOEnewXYHxh9Crfhes2H7rnvQ3j7
E4G+oPvumK5LP31Jk0sSbacdj7d3q0O5eAuPl7ENF8Td/fOtr5cvlPI0hB82QOyd6zJTgrqm+xj4
X9RjRiyUcceBKjKVSxuWt1saWSlO2okRYk/UZQuJ7GKpBkCt4c6FENKar0U1AlmH1o9YN2QNfnsh
Okh6yr2MeFoYXhAoNbXzpfIi1uplDn4LAF7U8dTKGFiafvpESMXf3euv7MMDgAw031iZ40ordV0A
nO01xFJVSY/sCT3w4qmbayxSiG9/sghSkyifX+OKiJY9T4j50cpaBbTcl/d8Vd+JKMTjzBXSPctU
DwWMMBU/2gCY//o8E7x14iahKhUdDswPgwpgoHYJMNFRwIV4JLeptEmqREBfQyzu2LP0YOOH2Kk9
3Dsbd3+P1ks97Uvd0UExaAZyyEfnJqZ8IX2hxrAyIG9DPcUzeQJSp2cbir2b4eqg9XEeMwXdtqzJ
ZkykG7v/wWKqdEys3M7HuXIkoMcArSg5VpgpZ+qnV4e3zs2ir7PlDpgA+UO0wPqNgDg3HaBue/39
MKC3mvIatgmAXbpET9DY/7kVeB6nramaMpkBWe0+/pQUL9uWwtoSaNpj4jYc1OJDox6Arcrnukcp
yIdWdueVjLwjngKgEnuM4zz39WxK5bf+xXCWH0oq2Isl3GIIJAvUnOp/w7poWLypeDIKVe7w/9WD
axDXJhWpOFRf+/s70QzIfBG3krgZLjSl+RlAC0nux6zCRp6KlD++9Cf7OBFRXfoY8iE4WfokZOmE
z+34WqR8iGNjUH97Cb8eNcS6Bo+E6siNnSJCnTDvQm2Zxch1PSRQ21Ut3tK45WFBGlFHtjfLB+oz
Ev5dO2Bo8eL1ygiLb9KgiMW28zV7gX+7XE/KS+c2IZ7EydfqyneiZfcIhbiLBeeQtskQFuGi7OrA
aZRRn51FYSrQ9CtwHckpsDJU1A3xPZSSMgXhOliX8nO8wwI6/DKfgAGFcaA9f69+qL0POKvGYRyf
3koydEztPBIrlJWmpuYNKWavj5kJc3Rj0U4Dqc6mEPemnlTDzJTJ2WKApd9r1RNsPs4wpFTIFkxR
TSqVQgAjdHkSDhJE0uIyklHFVQXFbALH5nqscHkOanaiXkNkrqYGgh90JaKU0xs8kfP9wU6M/etD
MCMcCjPbFZUhTeYsbJvcD0vS+UZ6ImyAQc7ZBeau9rYXjY9a57bB5EkzKi6nd+qzc9c737iAXLZA
fxQIYN3OWnWac+qANDh3ydRUFdGRgyb3XESBiQWwwT6PyXe0FZG8QaYtcnB4gnc0/pgt4HJ+sv54
N6qADZfiOjjQZXUjAZFC/5uesbRs+dBiEiwi2dUuaNFYDvv1J6A/TsqdORtEuPaT2A0MIp0Ry9F4
Gvza250QmBK15K257wrBjIKNnaGqSrfGE1YHmtgXzQelSPPKr0H1ho1/STO4TXcmIFzO6QlS5tUc
NnwVLDcGpqe6Ss4ZkLt64LLkwxR71Itivxe4KlwA77kcP63KwOlk5X91/xn1+WU0uH+81yBJMmDM
jAYYeLQNuz+2hFqd1h8YDvsv3FofItMcWXXBXh9b/3FqoDJUzcKbkz32Mmr8IMesiqMDiVT6hiuA
EAL3HBg4Q1zaKYVcagmp5mfu9B3ARWfR844JLAx6vcmAzCiFNwhBkLc8Bik29ymgETEVQhd7o18x
9s/YthQ1IrC+2Uwv14cCz0fWjcSuhebGAoeUEAuaGLtsugSY/pK84goGT8IYMF3wRtGGGxLzrU4J
sk9fGUJ0bL9wuT0/junvzGju+yE4c9IbgmM/CYDWHb6p89KT8I9BkNnY+Wz9Ogw8fhFC5lX7uA8L
Q+t0tTqt4n0ga14ohedUiUsQakrEQ35QnNBP9gwrNtDUKqIBylPPe66tXJCiEXycnHes4ESCWBVS
M5WetYMmN38NxaiapX07ospQWRCua0WV8ziTr96lYFxXGfqbjD8SKe2mksXnNmC1Otxu1Wyjk6+P
2EoOVJZvCE9l7jP9pp0RgY+q0F91+AUGn+nfsXsmNPBYajFVZSntjpHoBR/2ec39oYYz3cX8ZjMz
reKmAiz9mM/KLoyh31ESxJKCskU2T9GBexbpZ3/aFqq+5gE1UIdQFpw2OMfD1jC/p85F4BDw+MnI
xEFxlh8K85uce0ZOB2dhnNF7EJ4y/V/ns2ci/1b2x9gYhQXAGMKLE9wfApv/Vi+JVLpfXcW/nyjV
mGxfWflkHovxG47Y2vSVvKQQG3ysOTwB39N+BptKd8TTglXIVk7zPv5KyhrzmmuhsAwBnbW+v1U4
C125hMAuTGlyXS3o1CA6DOG18QjlPUUA9Z5otMppto9m53J9E77zYo45FHhBRJ/WPYvFBe31rjva
7Ot7Cz6n+6/c8JOcuOa/Zlbo1hZGozE8+HhLjQt8+gn7N+QkBt7ixUwjq2PLGJcGzprGcgDaH9ee
S0D+Fd8gqt7yHG/SAXSDMBGxne2wizLYFzCLJwSEtyYb4QISlGxPhUwDCyG0mRVvwHvS6DXGEC2i
k+YTh3LtaICIxt2r7kaEDDLSGkQ+tJbAz8eLD8D3Iux4l8tbFAAoT6e/3ERA6NGCf2XkB4JKVlec
5YAef10GugmGNonZoJuEwWEH75vG3HZbCfxjtT6v0cbeeD3H0w3q5kA01J8+wEnUIRhjvptVNieQ
C3gRvcKIBNogxym8KYASVCYEecCXzb8crmhGRAvvhwcqr3I9KXDlIQAhtOQQyoXgijN4IjQoAr6B
5yr9cEN43kSOPvYfAZfraxezUPJ1RaGnb7zhukKEU4Cuo7WUdV1jhFyD/YylSeI0p4FgsUqLHR7I
/1pXVxzzw1zPJ3oFfZl3of54Y49Sx6M4aEc2gVOUMvWTr3dV57LK1PT7wVViZUsbxmPS4F0Y1q1M
Dqp6j5wH2pETRz3jPkl8cGXH7OhJ+o/iQk8NCdZcuEyVs39PgNXdlzY0al8Ice25HSYiOtcGfi4Q
mP4vpCo/FesLPhaL/TJaltc6/9DY9vquMry9EfFfWWdbpC+l/BUVTj84+4gApuzedF5Ee4hRQ5AX
GMadYuLc/tA+CWWp+CYj2PEVVQR94puMQQLXz2eEsAqqxtnVlgW49PPOPOg3TcWf80sxHDWbnQM8
v1Q5dXXPdKTgNb1Zx6d4HaBGdpt2f1hzOmiGq3T8K12JDiwvdilerI9HZBidpvWMowcKQ/rsRp60
i+gbP6c9S61+/Jt2Rj8Nx75famcxzwRz+mxT8iacAUI4yb4Z9Ek6m8wfOopn5zrdWgOsUfaYahdJ
/qAPJrwMyKlsmm9e1d9VgiODBiWENrZW3K9qVhx4fWy01ibgv6ENyYXUKyRS0jxDwl16oZd2rdSF
+ddB/cT0QyLLyWSgKhBc5Pub5PATdDNJSwE7YIODuhfFERu0XVZwC2w8/P6/HZ0E1G4JrkGy4DXd
UWCzcG0utAfPngg4grx+uKPxfeu5cDPa+F1kwSr5JXYSXkLGGbri3tRItfYCinqcIaRjeOOkyDpb
BVSPVBLUa3Ge6inn3LBQddocqUWk6IrxvevyICAcdViMg04GLs21DG5ZamDT+FSS5hVWqMV0YlBZ
dOOCDUSeebp9hmq4BgX1mXyaPaZn7375vhou+Qh7flBdgTjYkFCzA8tsP/nulKVMPhTotR0uXLwL
cX0r04OQOMcqJ3u5U3mGMz3rdib3RCVfmUz3L13osfKtdceBmUz2rIZt3ffq/Y6FUcPEhJL0uWRt
4i2QJij2Abf5Xb6YVPekNGY3jFctqLYWexz0/7XcHCvmuNbZ4KhCPAOQv4ENcVYhrqQ7yMD85Kj0
xzcod5+MmiRLiYEGHc8ca3w2tUrA5MPRbpPaiaINNLpBOKAm4R7s8515ehwbFdQqjlf3xlKZ1qqN
KkNN77h9cx0IzXVdm6PkkCrRIw4us7/a3nkGzxi97Kw+tRGpcX7Z1HPrTExurEZBPhaOlKy9033W
PHQlUs6zjUPcOa1QrOQ4POeQu+4Rwpu0HqPqFmcYgLnG10c/oFzLP4QYBZh1Vl9KzwMyi7nh2Qh3
u7+Na920SRD42+dFhB14NuljVMo/WNo3KJB1uEvWBDNgA7b5epE+RluXZMXguqB0WBDBwY8+0M70
d5CBQhTGxs5ayBc9DmkK30UAriZd8XbV4cIaLQtMzh/B5/j1xV86jzRVmOYaKKd0B+s96hBYWis7
38399OksMslJxwHPAHf3YfaRCmUTavYxY9GBzRPcwy0+upH9zU52SnR43bLR76r54otgpESKISk3
1kTq9snbvTe3/v6TPYUBzakWZFCAZPL617XMu+ReDX1nec6ZaFazfi24yEWxlz2hRepKF2ls8+N2
q46+aW5U3HDAiuod3SQ+KC0RJz4G7e3hvDUBR40bQIYiSPdgICg0aOlXGhmd27YfenKmoLObxc4n
sQpg+DTFTRBoXTGP2ZqeMprD0KYsu+SIZTtUMcCLfrBjkj4TCPIGcRI+DhJHc0ZtWvp7yk5XLBmR
bcKZDpuIkTKiDoHeGiZ3ouBIJWWYg8edWDCPYfhgrFVy9pikRlfD/sc4rjr8IwLE5KkBqJiM6uCL
JcoEZU9PaJSsEzd5Gr/7KSI779uGg8HLuwjd6w4g1ofcZzpOmDQlBKYdd4imvGa2L12O6dINdaia
04XpSs8GEYAi048u8vvqfZZDwdSIwQpeVMJ128dSThcPvpI/T6qi+RNJnp+33LSSZb0HBiOpiEqC
84oOxtnODe4XCFCBJVCG8ozXgLXnalg2rcDDZ2NbXh7cMpqDaWyve3g4QqjkXcrdo5aZetr11FFD
Lvc9WLHDlYPDVcWRbrcqNK9DjcMyUSh/hqf+ApxOOUhhFBfpeeOHhJTVBFB8hHBXgJ1IIBXTQua3
cwRsPslWAfKRATS0X7ekDdGfuyQqCJMWIrEDBAC+kSgRirlpvQZ9DFYF69LqG7mLBtGMNvlvhdNy
QRBdjt0bwDA7Htgptd2PeWAYBLbvYMHrsq2FPTQaa55HVOpP+92NM3D1Kjpy7J+0CB5nKQw+Xxl7
vrwY5MET1TqokHmFp5KliYFnIsCMGloXG94d2pBbI2YTaMYNQYUM92T2Xn35S9PR1utMSVsFFftf
PFmsJz3uvBjCe+wJwfTddLqvXIb7GDh7stPQDX5x8pUgtyWh2cTWBkipcucBRKXW6x1Wg49fE/kl
gg1kZFV3pZ1vjZphAE8som51rqSbbwrbI1VR19XMm7P2Sb0L7etpPvwIcsbS9Ba8WzlqDF9J9tJZ
6JjIz2tEviQzyPb37HPxS9qDfOs3NvJx2U/ISyaoTZzEKO8LZ7k9wpaY1s+GZfWh6//lXbr3QlOD
HPqtEVsGM9At2mbRJmD0V6K2ElbCTz24laAv8HA1mmGagtirjPJnptze708q9WFSoU+1aGm2CeW8
i7rS/gBmj/Z61Bm3/qF2b5ZdKZkyTWefRe5klvwdvNzCfx8wgmJe/gf0HeFMHsdkrvuO9qi/QOSu
DyjSXFHgNetnljlWhhQ1YW2qoM+utICURSUTDssWz+w9IGdjlAV5ytrCvVQgytPxh27hdQyHxw9Z
KkfEMlWid+PT6ZsF6lUFJN4jfWDfy5hXbT0gtevy+vUcSwl4ySukgcb4BO38Qog5ryHuwt1OXtKh
s4BSzDgwpXrxOPIV6PrYSnM16M8BjLCRPguJBWPos80qeBtlCPyVe8vreKwKOdODfwfaPY9nFJ4s
OZZ+CdgRHuYVT4SjuBYeMPRgPQYUBcIoHjjy1s9hBXxHtjzuxP1nSf3g/NNgBQXbR5ABbSF80VP5
uYJDsXCTTfFPfvgPr56djrxX8EVg71lpADWCnL8JP26MTmI2qmUw0R+6AR4mt6wRjsRnMPqyYUYO
rZ38jPynVXjsCucBXMg9pWGRSoKAkMBrEbRrmcKG8lN8ed4di51nb1Y3VPQDrVPJinOWzKPnHRX/
YBoURDLeXCpAqcfirjGZmlgyc43B+p6YbLxfy7OdJEEujE1CWWyLlQpA1bmN555jR/VAgHM9C7KD
/YAaJmuHm0H5YCG59zOBiTr9Ns2Wz75K4C1esNbLDK+Nu6eXyFHz4qSzxeS57xlnykFtb99nU0L5
VVi0lHr690byzJGkjXMDM40LjTg+fBKrlcV23v1Na+quT0sZbbznVLRaAx0wYF226dNTSjRElL78
UrJLkhTFqelZ03i+kKIa2McyFLGUDQoxeAawWGM+mKr1lZrPai6E3dtrXW88I2wD+8v2fylFsXZo
RI54fv0rg5ztQdkfPvk4u94SYytqjHq7ClxEIbVAluvakSIvk04jyof0tSpSVnctvTk1iaSJvA3f
4yXFX49yUuvpZvWFm/sJ03We3+Iv3NQlhCi1U7eRIhotv17dIYYe+XafFyharAZwnKDaiOUeeW/F
ChC+dBRe8LEjG7YnPfNH+//ARLp0mtfh1dT+MhLREM6ELwBfash9vKdECdh2GXHOB1i6wjYuGoyN
vLcUW5xd6WTju9jgjFF/ouCIE7GXHY1jX1yn4qdhPwH7agwUi/c2K3ncC2rBoHIjKJzSihZzCnJ3
ncOemlw7M26dBYETgtxGymAIKQE0tBigdWWUGm5TSJxrGNwkS58U9oZ2yyRNbOEUUT9f43ieoOWr
9FO28/8PwDecrJtXfJJ0L6DFIyPlo2Ebq90EQfdLCm7yx/Teo9Y9s2qhPGAqNS7GaNckzThMgyHi
O2Pc/jUy0F92iHwFLKFO5I6nnkaaPyhdA4CO0jCNl/c5ErTJHtUthZ7vaIXYEKD2qHu+LFGyZT5U
lVf8P2ee6sU0nn4Y+kCGdEvmBoFgcb9sU3ZDEa7FmChpQT+wqKqhK3HdovZ/geyI0O73KgrfhouE
DjdJhVX/UNF41OROs9Ar0S5nWX3j/MG5fkIP275nLLUJD3ky5ExWxKvrql91iGQC5BLgR7wjQRJ9
hjLTKLkeDvcVb5MSGb4h2BiDVk2c6hY+w3yik/Xo/+pe4LGCkfe7dR1swzeE4lBu9lmgoUH6gpEb
adKmj5R6LpXULNy3BUwB0MmtgmZPyOOwRlK0KsG9QCSX9JhX9ePe3UySv9DdgkNKT32/gNYGT2MB
lZJC5ALk77l5kl8S1TVxP9331ozwI6I9nA7h93tdlryA95p4U/V7+1ctaVvykcP+VIFO9H2qBX73
heO0vreeqDC+KrID2uluOKvh7A0jMBJZ155nHU4kOWL8ynkdQGB14reezgxR/lqgtpuybBi/mvZo
wVMGCPOOY/7pfnPsHSKwX7aN83gNTFYyhtVwbz81pBoIhqiFqdx2gnLYwu6Ekitz37KPdz4J2EKx
fpe373nUTW+6SYJ2sKDVXQ3uGH2AsbVLjrJEiENQ7VRSZwdVvXhYJHY5xwEOTN2RaubxiUktoyld
ngEe40pj4JO4LnfjrQIwgQwCYsisk2kgPoAoY4hwU61ac2jayw0K8ZwwXrvL/JGi6XDQ/vz1MCLu
R6BvF4E56QhvcCUK2kLHvoyuDMMLezHQ9fE6Pfq4DkTS/FX2JBPr5f16PFJEFZzU15CeWOvmOifL
q7MsrszHLLkvfpKZHSnPaIqXQUP/I1D3DA3FAiPRNQH76hXVg43lG16IvyeY/QJeJ7dZF91MsP5S
KCN1zsPodKV6v2YnSMCfx5nfrSAmIai8IPppBkO68ejMw+X/iIA53unN0dHad69TGiwTAnqt+93X
D2lZmTZZzD/AiCdbTS5xlJMy4njRDC1pceS/Tg+ryivdAnNh4XfS2p7OHBwD2HRcp/+O3SzJzkZ7
KI4GQSGTbFU4HlsGLVFONgF2V8Qe7ZuhTfSuSLISvJ8ZNGVPUABJBTmBAXI9AMdzbFq97OiciHJr
v9l5NJYgScM78BFgcn5aga/da1iiO0qhCYLHQqZZ33ZIXjdTU6w1nXF+25Z9rehU8XpBbAjxh5nB
3YDpnAsVFvOXaSsuysVp/f5gPLW6OnyvWdOb/T5P8LtJEA5ozYU5ee6p4CB63o3Km6mcJesxR831
je1I8iuJakN1i0QAD/1w68gUt0QkFasDCyZyfJROS5CzQloBgLzVt8mVWFnko43L2L0qsUw5fK+N
DEgwuyaixI+jUUvDi3rvJWSelEOT0nMxdfsNwdlUbUxFYE5dr1VrVtGIiht1Z7vQBffStSfuVfxB
Ambe1dZk9kWFH1gmG98pxAVKOaGGrRGVsWUj4vMhsLfSOhlNspXCisGgfNay6Ehlw9QonNDLItoG
IcVl9tDU7M9JtpyAtJkYueD+zaz9LScfDlyhPwEv4/L+Md1uvr64Ze75fA15PBD6lsKvCYk6/GcS
W0k++P1w0QMgqfAxCLWw1kD3VKKwa30a+kyboRfYYCnlE1b3XEpsmIEsMsrIE2thSPqA5dFYt98h
e2KNfqvAiiWVNMGxDjMM2+QkM5CFPYAPoOPtXkozlYDweJYlkb953ypTtfAHXMoQhy3D+Of5F3YY
6dbCwkZDFEpgLF6NuDY9MkaUDIskT33ZVC92yyfU/AfWkYKrOtMuRV3K58MAMF6HZh0NmX1PNoH1
WUPoifiYNeLTAQ9Y0TZD5SlYOC102E8HovA89lwfMC6JuLzopsQJ8esS6NWy5wZQy5TFVEMnhgKG
JD+BPjaW/aehJ0S2bfQa0mYowGTV3fQ6rVKgQrSN0zpE+bYYj0BDjThWXJi9TjwxVrFGMqH7S/TM
ohPNzMnkk/XF1Zfkj1ONCuEOwgeFMlCbn5drbIR2a4apNZGf7NlrgqbSN+TBcnf1+DJhbBLXcUeW
CNNQj9TDMXwtfRWsFMI7y5onL+Co/v3spaDf/7t/EndASYwnD8s8HgwecrO7eKx3+/9Ba2PbZYtk
9gBpWTy5aI7iAfaEVw+Wlu+r37+kQ6OfaRwQI3nYD/z1vRz/UDQ40VP6QZ+dpXNu6pHem+zOjcfE
+YG0zm4O2kPXcKx0pUZCwR55EkAIUgO5n3W6zlvbZUo02LCpz+E5NPcW/sojCtNTMik/+GvkVk8h
A9e93DemXmiEXoDMe32DDxu/DqFHZnGJjbZFYZMCggrWShMxjszjOXJ21OduvVTVkDM2t3bUwY+v
Cmx63mbXPD3uNLQ9qDUVkA3R2Oca2RAEfHixVfz+8i2foVxxGS64jYxy5PXrXN+ABOFZr5gvVPdz
yS8ETz/nIj1BKOnsqXTnkMjPFguvZLxndOikfuIxOHRDhNpO8QI2GAr5hzAmbwZVXtU/AAcHv4VY
eVRszDUiGLEe+OVNHmhkz3fhcaMuDHhD1uZacesvwi0YJfkdeYiXpxgYU/KLr24dndMQnT3xRD9Q
5mhW9Ys9azHpWnGTY2KdtuvjNDJbpJbCm9WCDkCzs2mywQTTuzvfsCr/12tySF8A2B2y50wssz6f
40vb+X5V1/MsJrIrktEgogOXVxsZ2HiIkFMAQGQNknIpWv7xDFIgg0wmWapTBd2jJSn/7f3Lc0Yn
2RqN+76cuVmsdN6xEcOWTFyu5PNnrH4qfXA25aXMrID7BgiGekLqiIkcH/Zu99pM+pM/qBfwWVKP
twwbfBduqrLLQSww9CX3jFTQz+m29LXrqjiMy/j6V4YsC+JII04ESL6X4vAoFT3jFJweGTmsrsqT
Sv2PanHiOx2N/2cJauczEdp2PoSQBiPJF1VufUGYuCwuJua3saiQb3qO4MXphx1hFv1zXGLk9maT
Hn0jpfeg4hI0VuacaoELvfyNTI9mNNK5pFXb9Nea2ITdqgzrYUJlOot8Mn6HWqVElkxS2avLETfb
Gq9VYlunXB7bOOUyT0lVkuVwzoYiCj8TsqvcVklF1AyR64462yDfDJ+CspXvhrZbWZNQBm5opIgz
acIqJqfNIeIhs2JDoh7gFplAkxjb8NJAHtucYJqVMN0Xhr2T2t40QHmV7QJ/PK5sDOiSaf4dUFmJ
gonDd9pycN0p4DpjEHG/ux13/jS0fb3aP9YhkpsMHrEWkPdRwnvn1CyBJxrut3GK1PlSHa4cDRwb
v4Y0778M2V620HQoBc1YcV4Obe/eSVpNUVjHrDBawcSYU4VALwzcO/j1/4Nz6tT8lmFHsfbEn/Rr
/SxZg5L2PTf+d20M3GqtqBICi/74a0clCDhTSO/hYxAa0+nyZKcC+xbnjIQt8yh4gmx87oozPRUw
kV5pl16fF721UVcppFAtD52GXXqaC0yR19t0V8NdqpF9/7+Bd2MIGSa62EJeR+pekGyZdkyYTPpl
W3L0XHaR9/Y99m4WTNgqTed6t7k/7zMUaH8XdA7ReHKqHRAAZU6EKGjuyWXsgZrLDyMHtYHCD8py
K+Dt0iaD23rh+p808wLsSZw64bfmj22T+FYM8s9ApHwKFugewX1QSvG65M4xfUDSJgLMeUf7IC8j
kUusYwfSmfC07HZlL1RX5g3NzWjIP9m718sG95OvqRNDH+5r35qPHGrAbpzz5HMZGBo/3CjuH4f9
mMNKNmMxlIOPk1yLaD+gwtFnfY80ydJxnUGFHMOIlkPODWPuCkD0ooEEV4Svsn+QLDSMTPuf0oWT
ndsiac0ZdpVMNKpxefwnnVWmHsYWmFUY1eVlB5BxZHDbAXLP8F+954SCSGSwGwTmy9NkthUX0Iqi
299EAESlRcZpLYfhN4UPG1XWwUuUd316WlPYc5+P+801X1dydi1pnLFhQ7mzpPftioh9w5hz4gfE
QeLOmLca0QtBmZ0A8E939JxgQYParVB/g6rl+7cCB6xSPGlZQ57kdyd9FMUQkN7k478yyt+Nv00y
y0A2eY/993mBGPk4Ya85ilLyitt9cLb23fLYCftHyutjajbbg9YkPIt9E4RlcKKz//tImykCkdXi
9YGCx8JsKeHF3VfiaruTZDZ2i9wK4HsI9Me8GnENelKEWECYP8S8HfyKMrAZU6f3QPBbiusxMBba
XMXmQCDcyYvtSNeN2kLKmX8QP10UP6aB+tuzRAt0QGybNuBT4dcwkv6f5iuV8ars5h/9YI8v1R02
m9z3H1xIw6LraRxjrI6a96eWo3Xj+TLDdS1zrjLsjAff4bpQopWKvSokLju4Nrb7YGGZeNMgykdS
jO2s6p0XjkAHEwHtBpZdfB1n29fEIMlqjbnTAS7NrnyFCvlt2y8GsouN0uVllrsLKqdYUzQPcKmh
swGYxyDsRe53DMYYAQaiuCyWPflzJqtnpB2poeYjYwkuFcrWeLTJJKzbEEOw4npyUTivkOpPBP15
hk3eH5p+12RfyznXY9lH88tiGqJ/JcoJ2c7NGpD74tFWALh6L3YahpWuHdqgxPBVBMIx3UO4dcsX
Fc/nDKYCa7jPAss+8NH+C0qygnqOZIa5UA3/4bNQdvif9SSoUtOhZ87dCua1MO1rvBWgCaMIIMmN
VibyKzB1Uf93G3KNtf1nB0M142UoJVF7eVWDc3OmRbzv68EvTYu/hgWv0oeuhLZbBGpLPOiVRbM3
vQRhYiD9eYAreXWSZymVLBIuHDCUJ5V1Dc9uY4QzGOTCwjjxEpprvFKIvY8msNLq0uPxHLfG0OfJ
hO3XQAYrBgdbb5KXLF0q8QB+lmblG35104lQzKTaf72vKhN44YUcBDepYb/Pa6r14LECaiadeXRP
ero0cP2m5uC8AI64Qt7o1LamsZi9C0I3e4y6yq8+sknXMvq/7Z+fT8NU+SLn/F2vyyEXUsxxHod9
roSk1MIzoLnTbsHc1lDq5RHY7SN/tHm7PcvZF90n3bQLuvIzgcEYJz/loGRt00ZlnmNpE6zW0TNn
feOmgXanXVZgizEhCp+JfP3+hNC6RfE8qXXRJi5Av1g5VuVg2ERmOwM3LEaTkyp21lw6AC+m1Wb3
q7tfk6zZlnA7lb4ijVgbKkhzBRchI18ReRXzvjFQZCRDyBpvs83yAe5ZUOa79BWLzDIQeN/jzDIC
YaEdqtRZ5cJWqM5jB/FVi+h38n5Ff0VTg5RvZZypWOSfKPsSUYRwzs8mrQGKPlkEj8sqUNI2WctJ
FezHWcHhTmgCAB7XqSmV+zBHTTfzJpgmKuw02og1+cwUA+i+lxqxXlrehs2DFgSPKX+r3+4ChzSF
dRXgi1IG+1UT6hwMRuifkpF3orz7fQOlj8PDLG6vOElnLCYi/2+e3os9dUAXUywip32DrH9rXjlC
iHgcQ/GYYPTmv46Ry0BOSQJP1K4hx7yJTHX1uD2GZfKHXuECtoLzvrYV90zDIZSclpnUgmdX85/P
E6/zboUsIR2WwZrWi8U/BFi/OLE2ZhaNeA1PZCFr7pU6sNUkzyov7O7pNePo0O3vNBdx5aZqaYUs
FslNvd7vqPlOshJmroVKLf+ZV2sj3aN4aqSSluPX04bu8QdUKW/nxPl8vO8A2xv0XY/ESg4HzZJf
l4KisdUX4/Gr9JE98UzsG/dLIPr7AG6fYuThiTcaSEvYnz6xXw9gBjiZLqU0oT3qrtmd1YbkHEp0
7Hl2Usqd18F+/GLgEWq7acAQK0rIZ/pJ2BAJ67/CntG302G4tRcwvXwumVfWs1VyVoJ6kDyVKtOC
QUS9xW6UY1HNeoiwdFvr4OQVn13LlIN9dgO6GlC5r0o2hvMGDQ31tm7VhjkBkhpU/ex2MLq+03XP
f6cZthPhGiosJcTizTGKPqtIX8esx8rRCrLcTwgIekCmLVcDPKQJkEVWYhd8+drQi4gO/B5/dihg
f7BChMGiHvW02xMfvMeT4CeC9FW0m4DDSUMAOlpBRmgdZRkAm+IVvcS4wUhoPRMrSvXfroLiZH+E
q1Els0rBaCKr8LW8yAEtpnWNarbeR1HaQXHgN2534qDQv6uXmXWs+2l+1Gc0oWECsy9Er8c374G7
JQplo8tfPM/0GcTA9xCGCukVXAAEoRkcSLsVKMF/GsDQ/TJHXwHF+uiiit79SmBnCtVxXT08WMm0
QNh8FnflH8zMys7mbKDiw+9/8aOt0Wx6R8gaFbOog/tDuMkyXNK+RxiX63bJ/lO3K4ERq9NNB1/L
MiLJySvwIGEcHo53fErmn2eiuj3GyhGsg/3T2FffFlzunIhIIp7VA49Ksar9vibkMS2WfHH9zcu4
x4hdrn2BSlqeIE9X0DdVdJ3xNL4CaXjy8IFS+dkxne89du0G0n/C9J7fUygyueKnJKgNg4f2rq9d
5fD80AMbOu2LM5swlZtXN97fDoQsRhDtG3QG1bcFbOm2QfRCsT331kkL+6lzvp/X+itcLzBDILxl
tC2HKTo0ke5jw6DQXPYBD3U3eu4K+W7sP8BtqA3MAoGnQA8u4soiPWN4mB9ff3FjJR6JSK//Q/E9
XGjLohve8taJNCoUbbk4UFwhx6bw1lu1C16ZRz7ZGu9uDsdYzL36JX6NzoBNYpN7rwwKz31sI0wM
22M1SAy/2vvzqyOsv5Oyoqav75MIfsLkrxRIrWr1Ga8OzLS8OFdM0VZuszggqg4s2gw/TvA+m68G
smCgUi+C3Ny+y1uIOmyUGH0xHgLKwr2hjpNJeUnx70qDfMRIJHImj1RP9YMjNoTSuk2wO/RlccP9
u/gRTZEoClpkX5ZYt/8FZqEGX9YTN2O9HclZGwEVrNac5V/cM+irXEBlD6xO/Ghaj7meoQcMT4WK
mziDjKuciLo4mlsSdqLuThKE85cBHmanHK9a+j/2cGDAeSSvBdJGIqBhRCJE9EPSSsJmdSXXzG9k
EuSYD/oEehnlU4qrJURmTIRcGiqHpuUeMfUSiii+7+rbTSsW7Q3xqQ7M8OIQHZbhrpUdXWPE4G9/
QKEP3cpt2jHEl33jlFxpckJqH44RGofkORJ62KU4mgYIiowe2Mm/KshOOt+4U89I04W9FCbJJQM9
bxsWuw1sRdUZXEI86rgEoWy9h96t/NoILQ6vMVrDIhblsWtY6k2c4fQFujn6GXvVXWNn43tVLBrC
KYULD0SRT1YjFCbJL46mHUzjYt4gbV99BRyTDYlDV/JQusy7RqlEnMADsLSnwOXpUSWumBnCE4Op
JB/cnY1ag+/cIFrdqIp97VZTLNiSENHbLltrUS5P8Ql8nMmYWrx64bIwbQXEAceJrX1sGbY2x9Ht
mNuuuE1pNxL8zVfzNHSIsspwsw48U2r/VfDGclpt1g6h3tSkRcAKejQ6tFo7Q2QBb0bk6S3IFc/9
eLRcB0SV7gFoXpnnzNqEJG3ZDiE8gVsWeKQnxQDHhNc4PoqBCPLDvkz3HzlegBAa3ls8IGB0Ts9q
6856PgYU1vkb9fxkt0GFpJMv+1ynH+cgy+uWhAKZ02CeIQv8vQcDySDHLCoARNDnaz7LgoIQ4aEi
ScKiPR032lyLNeTQre9H8ZRXQCoOpXZCMjxNvkSwckJYcYWfyA/2gAFYcAYVkuqQq2Ys2kBEcAnY
lHg/q/wFilm6s51ilRyqxiDQcNPEPmGfrnZLEcRo+UZTYAPcAUMaH/buNm7rczSWN/sXiEF7iYjy
wxqiwtui+yXvwz4Uid77w0hJKEySVI2OB327925fgH2csIUmu5SAbhxLRsxLfjBJIs8ZYkesJd6d
U1YZ9QombIagOLtSTYGleWkPhJX4F7ckXz0xu2NHFqcQ6coAtK+oFkbKyiUg57/Ty8Xy1pRbztkm
JjnbPihxop4TKMDcke5yuKORbV9KaF9NkIhDS4ILckXEExucAi3/QKHkQQ4RAYxanuP5MIyRT6Lt
le44XU5elerw90zilZdGzxNiu96Tb8JrNvC1koKjiDwDjzSf0umH5QdwsTEYyviqkjxgeIVdW5SP
2E1ko3dNTnUjAhwNuzkCNh5PIkEgsgiT5vFQi3kMr+2c6OW8IcGabj7Gkdi86plTYPrhNZ8AVgRh
0O3nQnhis2Jr7+fAmB1fuI/a0zrU7ipEeVo5W+V2EfJTYMp4bO5DLZ/EBt0+PYdXQc4dM2kbhFi7
DZ2Oo1d9H+a/UX9dydpuGVozp+pp3dSWYYoGg69ySXLYB1esIpB8M6Eo0NXRrrzJgX1j9EWdQzhS
D+OsZV+pzaKTBQO83IfNI05nHy0CWEkMTTsF39W/yV56f2aHqqOZMfoPYThQ/isNMsNrKySgBTRf
zo6StItSM/XXMB6rmvnklxxhfzVVyNHd3qMbMQvClALt+FuWhEkiBU4L0Vy3IKW1aa95irSdTODy
nYO9cI5QGG06KEvLn+3sEcSpi16XELLCeE3gLqTPgZbtRsopCak1g1wz7fOfGCDpIiM8+nxcOS6U
f2wci+fWsMc4JLkA8sAIyBHl0AilB5/MtYTk1+Z5uqo8P98VpDn20wA/JpFYsTjy+7J7ikkMZbyP
Gw5J7AxALq5fka4r5xK8jWdGBOsSHqQrscRZINeS4+3vbnhWYJqUlEWSIXapDM8oiQKhavVFxGmf
VcMnggf2KIq+RgjrxnT9jsZ+u4NGNcYqq/UI+GQucivsFFjfWlifFE28HZJvgxNgxEIZG3WOfzvv
EJCqCy6BlpChYsYawLdyOeOW6UAWyGADmgIi+J46R62rPNulj68DP/u/9gBOTxvdBdf3BT1JflbG
1aT+dY6zcidTCaVy9usTBnwe83Cm8F1C2cDlvZHm2s2yjXAD03NHikqOtk9t5C3SHkcU4eVo2211
TIJtIvn3OhQUY2A2UbJA1b3OK2XSaK90Czqpwj/VZHB/xeqkQGgffGca8zrgNieZaB5p+ccSVP+h
+AdzQvbuEsTivomE6PMhG5i/+8ilb6/BWVMJwKQL4TOCzYOI7ZQPrWVY2i2NFPxRuCjJQ2ss94J0
5vcSS31tD2HP3/8dofFSDnpGEkhInYcUhNcpNgo9lFYNWm5x1ldBoLvI2eTr31v2waiuvNRHYTDS
oOeO1ahtl2IZB1aIPYOaLR2c6vHG9kJ2QGocXGyuvUEcVi1S7XXyoXn9lBjnuYSpJS4+0ob2Jn0f
gKDo0dQo3ijxs+A3RVmSlTBE5QcgxLQTWpSRB7yQCYzoA6snvzlq+Az+wyJj1vFeEGE9u41bt3Kx
hUylyn3GTm1qVJZrgAAb7Ge00iFjZLWOr6lc/+/j5vMVrWJLu/nSQktBUrhCbVUnl0x4aTzuz7vA
1OuR5iNJiNuNYB749dOQfFZe5AVZkwamQaaLke/C2Pz8UqjB8XIKWHLXxxoD5VPwT+HuCBI61sWr
614ryiGsfc+bMBzzl9ERXSKv1hOQczFFr8fNIt2SWKTJ44Q+IB2IP64iO8+20Iq/j8R+qTj9VB2e
LpSKWcKOZgL1NZZSZhOskKS1VusOLd1VcbfolRdQuIxaYcL9mKytrcFHtki7cxHmDcBDyz+8YrVW
c8LAVOdzvhygDW7OuV2NgLDLAi9XVU8BSi3o7y/yN+OG+a8XBQcM/0FlEB/ZsHCPj0y/9l2UKz53
ayZRTUOeoKIvNrJAQXOxNztmH8SSWBWZjdnxVh3MV9AiKrwobId6l70a7PGJUO3SkPznEu7voCOh
mMDJ8o3wi1vv7eryer2geTeLVx2FxhHHKQ32sFU0K3ixlhtdoJKxBU/XSE1pirikfURkUAG//av7
HBm3j/cfoulT7kxBwwUBa0LRKhNxqiSQDcAzQovfQr6uW2D/A4isLkLQuZqUuCj+IcSgNlnptwiy
DuRFkTQTz//YJuZ90h8qDiHTB85jzfgJM42B0dGEfSkYNLOCPtBiFdJCvY7mGqVGtOjEESPBNDec
Ji5QewH0TRN7gFciSmB5CWDzVd2uK0/b4BJgbXGZpW2mwQj7jgX7fekd5/A22eUQUwkxUGRKpvYG
+ea9uN/3Xy1+o7DG3fQzF8E1wAvhBK92RLZWVo2eOUenWakddzX869LEyDmNYBeGJn8L8g7n0yiZ
sTMVlhpW+FM7pqHdRpGBmrsfDLrTFKabLmqIOT6PC4oL9RmY/SYQwFDJF+uVJdroEObQm50w4uTk
8+wZeHx1TfxFAwlbC9CIrYVHclSZAknWF1EjwxO1XoXYoqU0wgz2DtzZTC+Sfr7FAfp+CS3aWfOB
Y7e3LUWkJmjSHPl1kAWwrvKjdmhToyCAi+Ma26qcM6b8G4Bcn95cmrQ6n7n3qYgncfsQgXYlYB/g
Xi8pXC55oYmPXNfR6NcLeqVGzHLtIhBm+k826O98KesiAAZEoF688V6OE9TAoPYZACEbUlMf6vAK
4Ot0a/ULyyAGkH9UXrOWPFCZj4t56LORNaLqw7gTLP/hrQijJmfv+KMzyY6Lbg7YwXxFstS+mDe+
K2209IRYzGlhrO/MOmWg7KbnV5HtWzB5uLRPYyqmloWUAV/AdJ5XVTblL9lpOar7OcIhzkM/amcz
H1hExCqODNG/S7Q2Id7Eq+KLBJHwpDJMtk1vOBvm5Dg9NYr51M8SiWO1ahkaFySBveYGsj0zS4tV
mVNCcjqCtO1zUn3XmL9N1HAeYJOfIA0ZWog5alLNKY917btbAdKoW50TkPPnoqFPUwz4DrSkLyiu
DGtwr5bx8Et0w8YjeWsxT/rEb5YRI9qyhG86OlW1mWie24nYuoltaoa/yaVAyCUyw3CwnEG6F7S5
eEuXjZoMuvtHqhTGzx/u2oEBLe1d9WRmqtltW6Usiz1/8gstH4JS9YRaf9PrrB5iGFrXCV5/fQ3C
UWP1+uH+ndXDKYmHMaU8nocLd02PWiRkdtyR4ZXwT9cYC6PUOAqt53SDisiET5bk087NfWEX689K
tdPL7SITBQc1kx3p2LFqF849g9k5BGTA6NVgRTfBX6pcXQucy1DcKFwu4w5IVbIhv0TdGzog+jrl
tRWdDl9m05GLHA+H2cvYTLY1uUSXaGoxcmpsOD25a8H5JwyhHbp4bc8OXmiTiaMjqMRoqbBpeOUr
2Ii1VR4QRlFx5Iswlp6rRenk3Oz1G6U5WLgAKOyBti/+/+TXoCc2lbTkFGURrOgZyw9K/E1r/ikK
DIeAeTqIbyTtFcbXP/usxrhDVA6E6fS0VSzRDQqNPU6aTMn+IPqhM8XAMztIYsOJcs1wL656UcfL
ezEudDNBg5eKlhT51tvuh+QPMF/piYTipw3J4wlfHz2qa/wPTlx6JU5h2dcx+lf3UziZnt6Rdrfs
YC8fOdCZQMOenM0dWkzNlIFlQfhwsWfoJiPZoC9z2fjYnQU7xm5HFWxyFZoBeGfnwC9uEprGJDek
eTT3AyTLX5tz6VR8A3IX8Baku4Ut95fTG5lpV3d+c6XaAybXwn34D+vyBt4wbkyeBUSEO6sQc/9E
RrSN3M3/EiT5GBVNnKAuErGRvFLkOI3QuNLG50WHM0AYjA+GMVFFQMIu3O68cEw8l1xCeH9MtEGw
fRzdvv51UcgjOqEu9K8hW9bNkcf07Fu22AXziS7biGpQAKRvLl6D2dMGLREIFpti+Z5F3aDCjfXL
/FICq7/FtfI08sDfAYXUzFwBcXgsazOCMSeKiRPfz/pDm7oLDmcmRV1zfx/Vgke9u4AmQlwvDcWm
NnizljII/DESpLItL1GtfQ7AsSyQQo7KSfMxUG/i0mM2GrfOvYL4fCRxrVDOQ/RsSswAhMmGz9/o
UEg1Z9vvi07bny+enrRX+ZizXIGVyxQkpmvZXv79Dt1xJn3XYbVtXlNzh8ZmVEz7OPB476lEQQu8
BYHARml+tbNGYhH2qEfyTohTMQyYqbq3XRUGbS6QY3gsQnhcUSmNxo4lXtBeY+OURuktuMY2dEbB
MxDHw+QEq84+21Y7jMAQD6bcC4jQNay7KHLGIOTFdoDhr8yCaVsKSTTeayR1xPfwSH50EsXcRB9Z
eD93QkfmhgFqS+uF8Gd8BaJ7cbvMXMFxKrXT8B+zDMKf781Kk9bvVxFv925IHZZuXzoNV/JTdXoh
cFF9PcuWA4ZD5R0/cW3xCqzJ1xKWSPspp/sphIZzJPc/4cdA00hPGPhsvb07ff5fzzS7pJ3plpXE
YBwre4yKUoclYEgvJ6izkvVOFXO9cHtVMGeIEzkA9fvPUiaO7VoZMJpWxNTyv/9DLNcanTOXbDvy
TgrDO0dFMYZfGRLpHGFisHARtqn4xid8Jy2KJ8bXXUcYji0f34fxo5nzi50Mq1Q5X6hH18udhcJ9
SbjzUvlcZEYoe4mcaRVb2X+jsbzhLsw72FPNSgNmSJ6mnE2Gedcv+I42COrs35tlmpL3o/nx1dBG
JnbkQx1MgW7QRboybRMpY3pSvtdtmkH+OC2jw5lyZBb+SZF/b+mTd4hOkINL4Cap3r5z19RMAfGA
x1Udmq/EgU/UveoQy9QBo8VayqAUdcaWJUFZtbvzPPCZH8KdwlXGcTVq7qiQ0rPSjyU4eAmxu2qV
eAOGc/MzFWmatH50pSB5P10BeufGRyj9IEoqcquDC+hVJO+bNzR9rCFkWIhhMIpOWRQhr+TCNNty
bAFnKGoKwbkcmCJ4heRWcR/GQR1TTBqjo6nAjNLhrLf24HDOmm6sWN2jL0ycabBcDqOpq2K1ThA5
UZU75kvZIIM4khxwUYjtYk8gVA7mh2AzZbnoN83kANjGtLxVOi8mw4HDv+7yVhlgTvhB6zsfNFiR
g1BYM//Yh/1bkfzDdrzCEj4czXI5wxICKEJ7oEP3Nflh3QIXoCa8mv6+1R1wM6ZW+m6QY0OUTZ5A
YlNcWsHyQnPURuRa5bLJbRPy8x3szEaUitGE6Yhr9s/FZIzpzBYlr56iDGyPcPLh+1jLU81tlJNu
73LeG6IYvKHxaYPP1gGWv6Dvhx7ZXvNNWsTj+LXIF0TNsMj7zTIzn8IWEOw9AVxyuU6Y5Mig9DYv
EzN/7HFO0npeaozb9DCEP05+vFLbBMzB9zpWzZ5qSG5HlLRT2bzpXNhCUBPhi5Vqayv9OI3FFLUk
H7Sb8EXkgmg9LgVnMDOYG5b0GD+MHdIeuqjGcc7BueE5dIQssr1Fhcjsa2TQZHSIAiDSJnLBIy2Z
H3ohSI9L9pVFW7rprgTGvrKDSjb9W1QYhie+51noEIkEg4Doxa8S10s0PeRD7MrdlLHnux9E3RHZ
mEFWWOsBqik/2sS6RtxOK6pNt6aF42BtXG5o6zRAknAX/D3iIyb8JNR2GW0u3/z8TjXcwxEaWMkQ
Cw84GxI/iekJcyLdzKAk+HMG7Qtem9GlzsrMd1SF8VI2HDmxhfb6flOQ3dr8ZE6XIUtFO8aLRgi2
koaJWthPews/PVMwkIOh88yHA7QMZgFIUTDye3M4l4xTvWtLB/nH6HpfyiqSTyL9LAcU7oOBX0X+
HJOehSm7jDOxZ7k6LmE7x5FO89fRzrPvR+vA8IAUcryhLM3PuP+M/uLUv5zDtXAkg3lfyjlQz8NC
DdOqk4J8xHmOplTjnDUz3tPfBgCkrfjIqpWsoqqc/AtTKgf/Dg2GBgBcn2zFIffE1WFtPFxu9DLT
GzKLQHj/vTqG4i+l6iubyZTEdBqQfj9Tt5d/yabDn8hFAviUxjYc99RzVqbZKGUI6lCyTwM5idip
ue4U44/IfBbgO+fDbq4fjeAQL6QmSecw+tbKWRcNpav6KN5rkyJfBEgMKblrC3Ni39EHXwO9xjWO
iReelQLMJq2Bkqpc+VunAvGBAK3hA5zuOd/JQoQVDpdjFMjvaysdUMcb2D3/eVl+HTGi4P9aakA5
ngUZz6IwJ8nEWa+sZAdeiyora43LHUGRfgS1zbgIL1WFsffZy66rEM1X5mCKQKdhdL+9ZZ+F0iQH
ftK95tjx9mUBYi0VAimDugE3U9cn3+NbcsnTpJ96oqSUDqmL3yXm3PEJjwZRHmLT1B+fWtEeB91r
pqkhtQ7ro1Cy7R5TISCiHG/ZLK7tOupWsxlKFyhM9SuF67dGl4nNypL7q93GFLnfvMD96ZIQmvWF
ud5M5ov4Kxdrm4s2qmMeBJdn/trCVanaz6NmXbFEqW1YVoFaEJmCe9TBfycGKIe/oMh3gNwH4d7o
cycOXGQfUoaooDq/s1ORZmQ/x66TB1vO/qMopvVFwofyXwCASRYcIosoPRK7o9CP3sYty1iEQ6V5
cTRyy5GjV3yhd23v22lUP1iOhdI5zhtzO5GxZQAKbVi/xtiORC/tFKO0KnJb4AqpbqVXDZKo2YKe
lhby+imvB/SsiQgOrYy4SXW5IFdDGbPDYXse9dkvVwopFDi3Fkisj+CRzM3AZNZwfybuX61HIykF
Z4SKTupDwVt9YCnK5Oc/6l0Wm9sCc6nLyAn2p2H9yU2jXBaTTHyJECkED+rrM1HXPZdKX/XtZyd9
/uaqK60xJXMWVPl/OU/1rwhOS5zEwwNUmBJ0+GqJv1JD3JDBg9AtJX4L9SXC2q59jRreN98QLkxu
E7TARYUG1UY4d6y06012MBtyUSri/NZxw+KtyAV7wK2vm1UegZa0BBTHfCwgIMRW5x2qkWwB6kqJ
xz0jK85NGfm2qvHOWxKakHvCv+lieZVdALmr/ojsQlDWte7P50aI01TsbuwbSeikf/ijOzXphNu5
BAJbNjDOO8/QHGrEBu0vP/LYmSIt3e7PiCtJYtjDtfKlJx3v+6X3VlpQpJzAC8WJKfQpQKLBTnJU
ln4c3gDtpwtHs3bKOXgl8h+8zLk9RQJv3hQuFZs06D3FG3bqITM6rqez+rUAN/5tk9Otr9r8C29a
DNZed25cqXkPIj5MnUmkcsVmpVWiXuxvy/A0OPMwY03ftn0HOM24JKac3I0T3kKuihHuvtfS5B+G
zmt42jHkQQZhOdnb8D1tgaTLgJmms9ZlmhCY9FaZzVe5AFtpQL0P/cubOb/624muZJiGWResb/24
KCxhglImTyjA3/nWNh/1e/ld9utxQZgkZkzWdXEqYSM+XUDRA2h+vdMMb8LoLqcSe5ysKhXwd5lu
MzOfGPXEmCIp7PWlq/0m1KYZepr0g7noQl4to2rDECCO1cDRWCr4co96Vhca4F4X+azCc8sFHOqx
Ff/Z8Y3swyWo/GgFPG56+MibEAsoWLlKJBLBrip15EA0lY8cr72LgPIpQXBIZNKFXEfjTNqyjhPm
IxLeEjqn9+HQd4ThxwKcxPZK8GfJQJ+urGuz/UsWnBkrJZf+M177rOJKJw40pJZpdUxwW5h5es4n
7kOYrMmVCUy6F9BnRxKl0bAEmZMv70jJxi8UQZcmSR7HVOZjU505HmOP+6+Dq6YZc4mjNcOLyRZX
uCi7Z1fE5c7Io3I9iAvoOO2i4ZRFzepyVW2fe0PED/zAsbQs1WDtEug9JNSFmDxth0r8YMi/okV2
52DTq3Bep581DGAHhOQAbO/xMjF6AS0t2ZLNFOiO/6+Kw1Ftbcxmg0pdIWNWhw/uXE97Fijlx3ws
DV9RgdXkTR73bWGwuWVhUccOAJSNyGd5EmVbsiEC0bEoNoRXYQYToAUjLYEv1MST4R58x6bhxwWc
qK/zzeBWKjy90kOcjFEpQHP9Kf1XUkX8EHbvpihh53frXukyj67B3jEj16CXojPz63birtiWvesg
gvvvXMvQghAAW33f+vkght8RSja/AIh0+gkqgwFjxFt29//pctnLklo+0JcUHKXygv1wENwg49c+
B7Bv+CzgP9l8GIooRu/Vo248CK/xZEyW7toTEnAMSWv5BgdKS/+p60yXAyilYWH1B7dxFXqF2Hdk
z6MooIi6Vhmlf3q2UfdwNwwx/qnrjOjBeeiuvmY05pO8jpdab0t3XBEvLyBvbv38L65KXXQbZBNV
AN8wWHBMjN2BiFI7RE2/UYJGz0cJyXTKdmRC1ghCy2Kbzwk9BJUftAAybY1eFpQ6H5qxPmZQQnMS
ZX0gJEkxwFXdpWi/gzwtyT3Vg9lb9N/+MOhHnMEW97kqjHTo8L3alberIwvQGNhAvrPWSTV8w2pS
ZTE0QC0d/AFTwmN5Cha79Ue8BAYGD6rsKO9Hvg5oNVZAwEBZVNCVl1fZ+A2Kgw0roegnxlMYnWd4
g8+PS/hMDyva0KiACXC3lFnVTfYtf3fH0/ulp5q4IZFB7WkHvNlRzH41RqELlIL3xVns+iQShKfI
yh1e4krYczbA4ReYgKfUyyVSL68R8Wxa6RFElfgQC7Mir695M+rpOUGbPEfNh5hHK6/G3u5glyKm
R0O5BOMyIfibIAbKYS0fLh3Ub3Autoz/Vq5HQW1IPD/z5I4ALfn8O71ZQjY1HbXxbgbRaTwuz8+q
T8KVgWYAbALr7RNKwev8X1Zo7QKLAXGh0NWFvIRDKjSwHpHTCuoJSKvZQcOTh7XhhTS4cVTiICRv
iUk2KCZOacecVTRbVOtVEypbauF9/8F5DN0t7+29u8dDwkuW2kq/owyTX7yrXuuarq3ua1go0mw+
sxdqdsugnvVJlHxenB5WShYSxL/fZJSOjTWHxb2Vmc43ZDyxL5yJDwKJHKqP9JNW5OdxbhyN7vSK
ylHSQUx6NxcW8zE93Vro5QKzd2qb+TfayqOf35pHBvBH/qOeXNnQSP6/QO87kB73ZOthRNap4i5w
IdyQHkEqK2GbRQurjOkYB9I85BBJqoefMKWgmxgC96e84j4lxxmWHG6Y1UD1TJ3B60bxVQTmQh51
ZxOHMiwdDrHrgVh3oKcSjBWPg+NIyNyjn3AtJj1k2JQ360bNCtMUhqhjJNYlvk2/fZuJNKfW23Oe
i0z29dRNOGGwpP4MwRcruh7e9b3rzZ/h8MDE42Too6IvOUtKH/FXS+Av755r0lnK8krPvQVCbmNn
EbFSaQEcrJqbZ/Di474D9H7QbESZBwcGa8Prg0v8B0MWwbSGGclNP7J3oiHTj9+Khf5YYc+KxqtT
PiYf8QE2aSFrmoe8YQRXIr0rboXuqdC5MtxvVgpAtBwzvaylqxBT1lqDHLjVL7h9aeX8fJJ/R/rz
fssXJnl8kcS4Ju/E9L6m3cGtEZOdnKmrtZYSJ9PpOG+d3CUApZfyQT+afCec13fCCIX1eHVcNoTJ
HDvOmurgJU/9JRq0q02eRDxluy+wpsP47c7nEQXJDY29YR7UELz1jdP0LV5quHHX+UIBTlYrxyCe
Fqk7v09+D1HNYE2x5lQVd2DnoElFHIqPZNt8ePoDhKgA4arzsw00PlZoAIuQ7y1qxPdyhTND3W1T
cusQQ7Qpzy3KAWo8LkShhRvLdOLWcy4pz8q9b2tRDLoNLSRUy8Oz6aQzv34wEnPYpJSqn3JNkslF
mT1V0voAfX8kd/4lWueIb6Jmq5J37RxqkAmzlUGP4reUYSMihHtDMXo8f6rSwPK07ePIs8JbydMz
wiL8mcn4EqFE4aj8BMm42xszxRjfxTRH4TKmayf1olkc+sD/4nuBZpNbxNILCVZ6MkrlV2hr+4dv
5afxaXRJsMC02AmmybvZvgx2cJDCn4d/3C3BHu9BbSIBxZCCXIEFX+A3mWLS+OyKzBXZL8utdQFW
GD+4QfZ1ZhltI3OeFk+vrRbURmFK70yr99Q7xFWfUlfy8MqMawmGfzTpXUkaMvFHgt7EjzqVr1Pc
P3jBH/RZkqG+ZWRK2HhLdpZMBzGF8Prj1RNoq4BgEWXmoXOQyfl1pPAc/vDwQXCKOQ5GTwO9y64d
vZgO2ot1wYSL3tfhBR2M6oJrOEvAHL3wfWWTiPSijrkQkUe1FGXkq/+pwrpvRQyxsbhVG+tLXYLs
iZKzNTh4RGZUPne8vqTDyxBjZjxybKtE+x+pk+VgIGcuYt9l74xUFz+ROkqUVN3eaWo44z1AL2Gu
btbVzTpbvKOD6PnIlWAf+yhpfu3IsUm+8cgQSAOsx6hmJbmLNmQAwnXrT7a6PTF1HKoPPW4+aglQ
qbOsjxtahWtn/CY6izuAx/iu2wAoXWEiLi6X7ZHmYBzBGb/xhHGcLfToNjiRHfijsCurXsaWgwDq
xpbPXRZe307Zdrk92dspY7lMYU9zh+t35rwstcdj4VrP42o9y+4vHI/K2/H3B3NPN5nUXu4nDiWY
rz7uouIZy7weF0/onqMGsqfSB10MY3sKkyW3c7K4spZbHGqo0MZUKhwC09vTwIQE1STiaPZ9sS2a
Rw68odttLgCtWwKeuzgmyMDNB5M8hcZ3+J0PR90yelxp1Ayvi2e9SHCVRoQYdN3OILlVyYpYSPK2
flcAiyAw1UocCuJ9819LOYvM9y8E2C4aWmESckDsdcUaGGzUH0cJdmvY3m2XmWOiJIhSrpk4G/uL
c8uuWotOgv70MM0hRcw4HOXFMY+d9Bj/HqQvzSB12fTKz0xaebm0PUhNS8rVRwYrb6AUd97sylop
Immf/FSgh9ukZMbi6zMedQ9oW/NQHgwrxGadPpL1juH2Lu2+FCazAWDO6Fv10ae+B1ds4V9YuCSD
OqgpoKdLe5Pl2GKgEpG4OXFdXu5rpt0Nk021amT8zYoFhn6dD3173wE/CssxHUKPtEZHl/ZN1cQ1
iJqi9EX0DpXy47ZOOY7Cxa9am71lfyU3M8C+Rg6YB4tqQt/7rtHJPaoZIvPGl2hweQVLcidKq4aS
BobRL91TM5xxaX/onaqvkCknZ46FpcEK6Suvh087VFo/v0TVtPbEEgT5NAQVgqtEZIvRVwsRknls
9aeje0ni7U1NniRSbvtRSMQQp7F+XcXRLcZxD//KM1uffEfNeZ3cmLAgD90xJ+JBV54UOlI+tRMQ
VZp4WuyiDukSU23h9saxwhNwgKfKDzOqnKDll9eNuVXzUUjnYWTOC5SqwTbETey4GgkE+2xtan3d
H/C8CYgRzICAKirZ4EQDFMVjAtiEWA911shjP9c6GL/M7RGRqHDIJS8gsDmISNdCg1+lJpUseX18
4YENQzFsrV5xhkrRVpHz1YnmPG/p9y7c6Rf30mbEMnqmZ9/BocWo1gIeaIsU2ulIquL45Igy9ZPo
rWSfTa/Zu713tonZw4YhkVx6hhgh/vnmNZRYWjeZ6jlZcDgHWmMTmg5yINbHCJoXzwF4NycnJTza
HKhMtgXGGFreMbIu/Nr0IL3C8FL+qemlOaYO0hXpoyxb74miHT2PbmdGW7wFgTGQFDDIL0qo74Dg
E+sAS8rYrxZYZEJvSGkk1GYh/mHBuLJk3b5KV1UE1cuvdX5B0o+VGstEQW2DFQlWF4Z96qlbFdf5
zRwXidWZ8A9zAWzmDCnQiXjX80XYEwIKy7REeF3nVewp7ymi6qpUprr5dcXlf8bXpIhC5nr3dm+0
cO3Cyz8+NPqZgjaXrfn5LNKK2OjXIcDJEdwyKofE/qFKzdl8vU9Mwffdw22PWhNCOICM/ZokVDR5
6etNawRo+e+IIBUf0Nc+ca2lRwW8j9/86qa+16TINdBsTQwVEM7WRFVu/NHhBvrlF/vrCt7jtbNp
qHdP+D5kOPxy/qEhuRybyt4jvdq+xfx5kzhlxJXTGZsGc8UmaG/kjMCuXHOj/iaeqCs+S2nfFoFI
6AGRAn3XgbF3MclK1QuZ4uCvK283pJCcTbHi1WrgfSN8X9EVY0hE2PAR+4Y8KUyyq0sxUDk5ca+j
Gb5L2BaQSARq1G/WRn8rDLNLmPpegVa8h7ZcXwZ4Go6UJUaRB1oEA9vhKbzx8PZyNsg4W/MKDDBJ
wAbsZ4qnkJFaMceKuexLT6fwp2bm79e6GGi0BU4WSpJ4uFLFcSrJh2y6YeXJNLYrt8RPefXw1J/C
Fd+sWlYnaOR0vafd0RPbILZLJ+8ccH6l2ygV5ko+jNtd1mJrPn+BvSw2bidfGChJDtkGmMAHMH6u
M48V1a3LByYbM99lPjgR+qHjeGuzxsMDYNVn2OrordCc9R/+dvHMhM8FNf45Z3e7qPtlBqVP0t+g
WF3v6oKPZR+2RkGQj8I4DwF/owup5slCVpMDsBXDL6sJJNlUZZoqbeS0KsdLxJ9XnQz/n7xxWDLE
XIthMeytLsLHBNtP36BXP1rFYK6IdJGdMPNatBE5E9OrfV0KNqueycBLj5j4xWCcKdWhVP0Mqeyz
Xpj/Vxp+Mbl6hPcc1aIuvdBfN/ThQrJxr9wvB+2GgyGHoPa0qJYOfkJGa3iceglNyM0J+GCN0OgO
yMoi2ErtKc+W8gqlPw0hHSahWEkjEWtJm0ri1LWzASsBzYc1u0fkcfQJNucsb311n7w65fx4Icyo
h1ub7HzHmx575VWPYoylSF5yslhdX1q6ScamBiEMx4ehQiQAe7AvL6A3FOwMrkF3nTOsZyj/Nl7e
ufVx0hTYxLk6q14N9L/z9sD2+PK9/yta0Pv+AsL34iPCnjbn/1Pfra0l+2JRrc9XH3HAVkDluyzT
LAqPObF5EvnSa5NY3ESYlDlrU2mgh8O8ixru2fKUp++3ddPqtbjv9U80Vc6pJaHh0AdUgqy5AEZ5
xefONnB5XTJvKm1gT9g4d5BtchWYDvQmBKUmW0MBEqfXm84Xajkc+Fx9rv13sWQhjxstF3WehF6n
XM19LWDTi8QUez+nehUOGXla6ycDTFCgn6A2iBdL/PplkfIn1hBJpcjSRPATc3U8WkBhG5agzVFz
PRMWNSawmAGaXEPRYkEuH1z+99TJD/O6LpdPnXXhb2BKOFw3R0xReMhM/rdfKN86pSFI8+qHDRbV
lxmzTeYyHrhNDpkTWJUd+chHi3zMCk24dHOKFg/uKRS2kJF96MyKyvhrO3SbcFvj0rbHUbwzxojA
U09nLbSMokwDp+cr5yGdSjNO7i7nGvIkfIh4BYgfU9V83sx76q0tPi+9GT3NmBvXz/XelxFtjkW0
tqxmz1UeTOUnEiWmW8HC23D9S/DtxXaQgXWbKhP8Ho6js2UAP7dwH4XykJOhiSeFSxxZlz9VqQwa
DyC6yq8sLMsUa9spXfrL9ISQzmfXeDMUYkgAk2uaQbGYCiF4GNKgoOWbzqSPHyYANijYxJnaF0ev
9YzEWmPXEeIQ7K6DwffaiPFc4g+pvAwgE8yFvnkdK/NsoN3FgiAd+jp8MEpdhM4TBCyPhYfYoI5o
b4Xes/LuosbtUzt/sZH3rRnec6xf0P0Pwuhzp1rxk1Ec0zXjqUUgtzkf5vG746nDGqEdILTzyT44
pCTCfuebYJeR1/zc3qD7kp61iYhuzssUFvsKjh+n0kN+9QvzOZ4U8bnWPHpvsRd/J4JnJUMtdi+w
0TzUpYcfYgBEJERVR98EOdjVBd3posR/OlERyd1Tt1/m9Bq90IT89MbvKLAssXBdemg0ToehQbMn
00lTXU5P1wiyFfdy5tCbkNY0n44nIr7zHkvU5dv+CSZEmnh5ofyNT0TDg/F10/OoSgldpcHFag2f
bweQqlx/sJXj5+FyfDRxgQXaM4yuTGGmaNAozlz+g+dgGcditZXy0cF+M4edoxs17fBYBGETFoJ7
yJlxRy92/IKmzcMrqpZCXMkzFvrn9dsiMq/nhOEQu5ZLkyuI9TT7X5evZ7hnvyzJjt18bMM7tZp6
CjCCcTTMYDA2sIjRvLEUoodVe8XissRfbp9CqRfJpPp+xZlR4t2X8A2Kop/PFguMd6ujL7fqCnmv
Gw/xzEXitOqkjNxZAAe+EXd/NmkwqsgvV5e03q7N051HPvYNqSQKbGYNF8j8A6SJLl5mMtKuCe55
aEf1w/uuxEudRu3Xcp5qRDHFiTp4xTwhOehg+GN7+QdwxWL98Jbk2v4oloRqPlOStkfcyzXBsn77
ES7h+tNliTAgzBtzM2dM8u98jE5Qb7pGUvThMYOPMD8YIHr8Dst5+BON5GDfp4Kpb6m4IlBwrMSB
1Xg9chyB4mwEDjUMkPqylLyrcKpWswWBqJbP+brkW0K787zWOvB76H0+yLJf39iW+zAiAKVo+/p8
Dz+byhqZPWZ3rjjz3nUHvKCJm6a0JaP/MptSyZAy1MLhPCkxrpcDVIMxuIo7YzSsem0dPkz80Mu4
ip/JIQG/VYvfHSR+a3cj/TJWoxhNxlUZoLCLA4w+aHWFpzkQHfViZS6JuFE2agyaIQCqA8rK8nyf
3miigsSBpWRfHQeQBvmkmhh42xr0LoOHwxPTZfDdoKCIK8fKnhhWRXp2r2vK5c+mSEzWYLouorpv
VszKkzBetnIF8U8ui797CPGiJ7UufY2PtjrCJHBE0AK1E/I4sUY76R0gAq7QHBycyDzzJ4ez0E8o
njt7lJjV5Lzv0ao2VzZ3hPSCTqh6zTaBcPsqoVU4AQ8ob9hudLmeeQbOp/Ur9/sBCtjndNcurKa4
N0+bGB8ukBIgZIU0c+zc2bqTx5n5vIcaGpHXAFH1YvkwFsGcgjK9D+4rCNCtDcPjBDX42HlMQel5
JQ9O+rwBoJ5uEKamWS9jKVYGOqM0fYhqnuKA4PsVT0WDRaJCiDaYAb70ikuN6HRInIYWY5Cw9qnK
W/fA6ZXortsa2ZTzDo19zK7lb8AzOauqnQUR/gOIWFXi7u0zvpGSdeMEfVnuwsde+iOlBdObzNcr
/Emj36p9R1Ruh1qVfBym+WcTiwXfxaCrtPy9mnT1nA8SDELbzlq+YKjIezEpEmgQqqE0k/Y18ArA
gY0cT2H4tE2Fgy+BawBEk5147hSNYEA6zG5HArpt1dp7BNzdv6RaIs4VpcR2xlue0hwKWInyQDXL
GJ0XdukZp6OdZazOt/tJHj9Q+sNQAo5ubvSAbW6RlsTLLXlLJ8rKiqnSRs5bKX3WOcbykASg+pwp
Ou6KmX9/7/ikSQ0GmEAHqzAq6kUaOV/cBB5EqY1rV3EWCxPKKinYri/Qc+UcknyKyREG8vnXEztW
YpFOjulNvCoJP8bX0mfnpXnU8v1YYpdjZycPblTV9wp/zOvehh2Ugmbj9l/sFO5PNjzwrwll5gSQ
MOadZIyXGk465ahr6g714fRxPSKZ4ATf8OKNgxFzTQdNbSxPNW4Qzy7QOxLkLi3OpYdn9AxcjAa4
7H+YiaBqeIxxQxfdkPGXsAEfbTO8dSp+F4E5mPU4NqmL98n4OWqUacLHHNR2jZ5WH4rVf2VOfIvX
Sxd/xUj/oZy2gjrqpWF+lv42RtfN5uOCKOyV6yn/Ln5lfxMEjeItF6q8qG8C1cgjUkiUAm9LMv4R
Bxl8pY1eZFfdVR4E+Y37xVd81W1W5pnnobOxywi/yl7TYlO2Vlyp1Fpb0v2ipiqTnQiqePjBx56l
DxFZ3DXtJEMA6yplbILhzc8mPke3Ao2oE/1C9c5CasAT5wm2g9GT/NtW4ZmHQNHlLGcLk81Bi3dI
Foz7XdCrsZ/8tRhvw4iiGUbvtS4N3TWDmwbMJEjlkR0t1z+zxzixXS7XyFMIijA+XemzMKrKtYCM
fVdtGTeV4BLaHUYQIIdHLAqONOpFKQlOGUulNFeOMOBORCYKnku1bDjNfemIO5vbETiEAAoq0BKF
7KaDXahNd5Lqkxk4lPmt83Kg7IMvxisCfpzYp6LR32ZjnW6U4j2PYrjuobiL4iRZfFfgIlxbpnMP
9o4MlyOoHFQWE0hGcb+VIt2lciOobNqyE0F3Ht4QRlBS6hnpl6PjrKHIr05UZ/VSFhYI5n3ZrCUj
7fKtienmp0wAPNMtGnWqkq7tRCKEGLz4lui6ttEhGi/fsmxD/6WwOSskrz23y5t3goD0Siez17GT
6eNT911CaddZQrk2j3yUccpS4C5GwKL4elxVzdDh/SmghFU+VW8zJ0Hb+jE2Z5esyJpfcihMyhT8
zVn9BDjU0R+rTcA654FLukRYvGcbp1LJbiIJxotktqwZ4b0rAjVc4TGBUXvY3DElSKaMoSUDjZvD
J0Gme7OR+0D9tbkx7znG7HRp4kuhb2lK4odENFdD5S691cyfkgTxCZyB1MLSv9W/4mVQ26neAt8R
6pDpzvpKGVLdCniD4ogZ/UVjQ2diYdPnA+nccEsxvGGLHKDrOvSYEJ2gLYtt6uF1VLjkPqBYwG5S
uxxAdL67Jhjr+OkLMAG4v9e+6xLwqW3enua9HomwDXlXAmq91Z1r2PMkCcYVvty9PJCwW5VyIt8m
UfADOy2Dv19gA7Ju+KAPrNh1HC9/yyOchGIN8NSd4g1bHBmiD2CB9bBLn8o0vn8t6pHKN+jx4uqu
tJc7pZCSqJX2VBlghmlpVPr7PP686V9zkNPLkahqH+ORhU+NIORhurV+mkSJsMfUTYrNJHsqzpRd
3o/tMxbn5Ia+mhncMxO1ULxI0EC2sh5m33jrmRavF+GemEn9HQLQKVVl0ZF4MqS9oxKK5zF/l3lR
L2cER+j+BqlkkjLIC8s2+91ovHVmpt6IxyMIJdu+ukcK4pUgmzfP1IMaC0I46qobgM1brufTplbZ
TEKSYzdEP+TrWBhWL1LrC4kYQWxyO66DZzSARsL9nwZt3HYQ0O2QtP34Cnomh2Fka1FziAXlDpFX
EJotWoQfHOKEQQxsxg1PEUx2YDhFOkgl9zmM66zpYU/DP2pl2K6TyWR3Be+LSGuP5mVQ432Jw6yv
nlJIAPWRVgk+9QmY/CfsEihVe59I/kpqASgi/ZCqOlO2rUYcvNBFIVsByRl8cWSQ7Den6MSvQPL+
HMA0Nndi98xlslHPeKwwxnk9E6zF+atqOA9uvorkklViCjgJvo78UXy3+Co3+vyI8YTLtaBNSkIA
z87NkHZpof3q93c/wWrXhPpU08JC7DdTrATGyYXEQaYpYDY8XGHwemKBHqY9O2/xnq03jja++fzo
ybxX5aOpKGobG3ckOe72cF6mT0m+0AXes39hz1/OzAiQKLo0cf13LVbFYQiyEvUXaipnfrGvJXer
oHFEHaIZf249mZztPpXcPDx3ZgOLOSz5vBoPdO1wPGko9pdeQIvpbtUTqcFUWHTE6QozY9rmA7d4
z3p1+mbbs6QydaYB9CCVNcYLIZznrzxXrIKWAZ2zPRzGycM0BCztavwlGtznW/y7eplb2jfL7cX/
G06v2VhNj2LJlWU60aDHrTSlKoxUUx3Fq+3R9TTHXBFzu1ClVFUf2JSLWAo4d5+DOESqbcK1pK6/
EJVSeMVTRY6zaIM92+iFr8psF0OnKx9o1oBSvwwa787HVoEVVVLdjosJuWFHm2T/RxyuQQ1/0543
ZXTPsJ7JSRSfK0fJy/j4Vs+rpABJjtn/9pxUM01PWAk21pFr3FQ+lhhidLRMesW1I2ozTYBh9CKs
4L0yY+AUtokruVCSHqmAhO4yINCoZv5/x0vPrlYyu0Ve9vMjs7a3JjgyGlS54iSCELTO5eUiOBDp
NcG2F7hTjH05T7s5cJKS/gQJUHrprogVJ/7mdQPpgeTKccSFBj+d4JsDiYAua8qBSUPUYmIjgFxZ
9YKKFoiEF+b/q3t5Ca1ZE/XuS0t+ZjIShB3rr0OCBaQMfcQ3rQ/ygyBJv2OxmGx9kwUZXzXuX7id
OEGneLHh2RsoMbB3rtXWjOhZws1bW55z9snzvMSrP0Sw+Zc2FAo5XKj7prlHs4X+eDpt2oYkkSxv
q8BrutfPeEQ9MHr78z+gaSHmv9Xj0iQzhv68HQFZu/tNAfTme6fqzEi/X7cLiKc4XUw9mN/YQFUd
MquoMxAjFOuIaQtfFqN3Qxqir0F8ohhJCag27tVeViwIAW3LPHNPvAc1Xt7ynVHVC7Nohs04umk9
PK5rVW0VQdr6OmvCE/CkHo3uTqBbgPEfmykb5hl2S05xXcmp0pkB55+i67fdQ6VlTkb1tiy9HGM8
7L4/I3YJO/QGU0L5Mh/fife14+t/n5ZbHz7gEMiZxBHPOEHuMLbC/ULJm6qZESvEIom8OkkUe/2D
FZPZMwhEkUwe4sxVqQNCIAF7djocFnzktdmwoXf2hI4fCDGK8WePV5ibQLMs0l+QDVjNfBzdkIPr
2QLkYfNkll89EVtfjQZNwteG+2R7RlqCRxR494ZGGCzCz63QLumVSs0vedLC2YTRAd4igdp+AZXW
7FBv6GtBj1WJFcpDvsmy9QpwGrO5TJ0sDhtdLrsyGJRcLuvM/f5fQ35L0xaokwEmbGJSDBzSk0tI
CgN1g/l7l/JdrrUMexGUyyob0LEnbBZScQTdA9IcBVJgsR0hKcJ+X+OxIBWfG5v9F7MeFVyzaou/
XtEnOuAvcksit7mDeXw5pq/gjRgOt4miByyrdYXpembRkx8q4raKI7LeSgpfFqRtmqOTwVzrfzfO
Ko7NgP+ujtR8DMZnZJv/p4hkrXe5ViY8/HBT2qPzFlvjIMl8DQL0rmbaMmPSIJSa5KRD+q855EvO
wcQyvAlx7Hr21Gx4F1nrjfeNqHDft9O373b9DWDg8uIx5yGa2tUGz8Oa8E+Dj5VfgRPvO5Xnnp/t
ivbtGjiU2sqgbWvoaLu27XjGnqZAHwGSLQamyLs91ioliMEL1ea4uGo7qicQNpXqgoeiu4I5+8B/
+nu2LXcYzkGDVpHrkFSMGCti9oINA5E39PC4fxKTJHLH85094oTGTd8ePc6+E8RBbfbBBr/4PQV3
oIf5sQ39C3Xpm6XWwLwNpTN4qmi/PhCAxhZ0CanKBzOi6SsRfjDXWHYoL7fMarVoc9oH4HNG7wub
eqAocPZsNYgGitmWCd4cBBgRw5Opm3knRo2FlekACCSWgAR/ZFtSLkvSYeYsivJ1I9B9e69urmuw
WweCvspHsqNbUg4vYUALAx+xMB49pTaS0Gasm0MLjtY+T1EJrF7fQJuArqszzadFtqpUNHrpiMrB
PSTZ3eaQR1HUzFOuUtOvxvst/M7pEFKZtRPJCGGqsJtgdSPB8zvg1/V9ur3JoBOi2eeX3KeRUbFg
gNIFldNZDLkh/U14nuJCiuO5TMrGK8CvhZbYmVAkPpFSiFPlNXlWaxxzFezyVG0HCnTRT7pn4Kdt
W7MskEi2IVbwsSsp4v6rBATHslj4YTQPtE9tOJr39Ww3AgatxSjfnvvP+4WBz69lXmI3Y9LFP18b
FkjGy+PYBhzgcJsorgF61sFIZtSDmNcBo41oyMJakA20fyPLcInoVix5fgj+44GoQMp91KY05JYj
ySY/WilYgJ6g1v7iHG3l7uEIrdAQWXFZ+YZdbOwwWwJQZG8GGPgsxHDxYE0CKlZJjXcO5zEb6X9J
PDeQ05T0cgMMiGUgjqV4E6sKC9Kypq25TPB4KZTh5zTJy0YJ75Q2CDtPSuZySwjSizraUk9ogkKr
wtOC5qzPnNXvaIHbOy3om3AMR94ws2ewU8qA/fKzMFx0qyK7lxc9NNCSodtfdYK43HnugLiwsIsp
zpAEq658QnOb2PTccif/hzM5TgA3nzQlI+lZKe+0TvvBtzA5v6s9NPGNWbUIsM92N08RMGCMf2CM
zMo+iNtzlg++pHGDk6ccOKBtsAwFCUO9DghbtuMVU/vDzLZ4j8nqV3PMz6coPvYcvs/H8cwhOgnN
IVR9e+hAC8jsAkqa6vGzJtmm0aBy2FSuxWXBJYwA8K8d07AN+kP4skddipAUsfY2eN2+l08tpAsn
Tn7T+Lh8sq+LysfvUSoxa3HP/xJNpP8nhg96ngpdqC8L450fusOXGwZLX6AGjN0qHJhZQwTNgCMj
LcQrFsuLCuRm1GMR6vJlTWhpIHjUI4ZPWbjxXMew55jENX+iq0n+Q0DRXwIWqQn7jlhw+VMwSnDi
muLqnrdQtABZ/bUc/8xROzeNQfo3IV0IuczsHpqoLNX7waxNXVkX9tu/MWvYzv4cl18BTebk9qKM
WUK9quiwwDMjjp0SkpNiuQcts/QIeQ2OTJ/Ht8wLMe62W/dtpw1egGlqBkcxLWVGDrL1KxzhU8t0
EfbTMLwabTKjgAYmlJzbL3Kdo9WTZ64+coVz2y2K6eXF178z9D7/TGnzdlNfZFBhGHoBKn1jb0UM
LN4wrFPCmQT8m4N1xMxN1KUaPQUQtdWcvcdfphALNHkrv0GesxXw/+pj9zpjBtKOVfgMd2vWqwR3
TLJmxxKUvwWVLPU6sbaArFPE2My7RSnLcYd9v5VoCADPVJ0QarG1SvodhMBRDT3bu5i0fXHdBkOb
ztfg+UOZjhCONAc74RhyJADx/LjFw6azBRs2sx4zij/tf4xy0RenzpNsBT+C/17o/k+/Ct0FhHor
8Klu6bcekPropNpdcNat1cNszqRU0T9ItKqqgMbtMOVE9/yeFdlpzhCAyGFpPQHDDOLa9TXuYEiP
eCurc4TfnUcn2welQoLWNsuL4pFrBWCYyMB6CJYxZX5GnEgiJf/0nvpfmR9HJFivktuPRJ7lLd6I
zSObTRyEU4zknwjqLLN8zBcPbucalH9TXmAXppoJPSjsewjnpyNWDZBORQpf0rV1YjWuRE+bFNft
dnyFKUOztYp4vpPQlg/6cK1ugk7gDAfvXaf7fwUYimmCXxQzkuw0ERxaA9E6XFaGft2QjRGx3DXM
Vwx1Sj3BlrL8msBwpa6cnNbENo+Wu3En4yhl9DU2yt4OihzC7d+g6SGwJ+jpVh/QpcnB/PKGsb4O
5NHGjysVA6HFv7RODUmuiWDLYptJC3RhnNRUGFFGCm3KSc0UYAcEtJSSnnxh+j5Eb+yzPSEm/uhP
W6UQN9DOqDW/EULs4tbWGLq+WCcw9TyXQDuLl2VbiZ6s5yV4jJJhN4Q0BmBkUswLdmLHK6GPwadM
YqmzVqCLKH9PwFIMM7SEOhJAJ57fKHgGdgZStG0QDnifRp/oFoZGGIpBXFozcbs+8lb4N9OpivsD
sOA5ntel9AU5l809FsypmCvvgSI08q00CEbxdKjRDLycD7o2DaML11zIvVLSGNv6AiLe7fYfa+ih
xO8llmbx81IJ1xs1fNwm3TMCUhxTtBw8MLhP+3NnLxKJmzjEpa2BdxZjMPJDWUi2aZ1xPh90q7ru
pK5d8tUz2Fb54VzbjXDXPFebBKd3EzVXuP0OAdfvGduFKm3WHym7/NxXc3d+2qVz8i2k7YVHt6hw
niVridUPutSLMR1UQqroknx30ecijGKL9lWKTGB3T9gCd5uzrTCNxKNmMj4STSwazCBTB9jeeJrY
0w5ThqKrHonrS3qQcE1acKtRU50Wq6SIPXeHV2tg8XfYGbQ0lnOgEUkIUsXTX3hgs4BPNZzns1QW
YUAbqK5ama+t+xfl0Amu6opZhScn9vBrnrajMeGuZqJJN4MJSmy2zkhjVFYbwBpq4wxCstdKXvKL
V1pnfYK8ZW8ISNVQyrgyrzY+0H7LsrU/cyVODbeb9/L+wdWNbYCtuhR8hT7/3VJ+iWTFgh2OMNMP
XMN9ZkucT2lYIxBjsrG0WIcKEJtX9f2JvlL1c7zqkxzn2Sf6TsPSEslbElHEYbxTyvCG9wQ65XgH
8YAIsdBU2CjP1d8Pjq9dVF/xoQzWlm034f04zolCsGyFJVBh9naW0npRdmEVVsewRhVLjQT7t4e0
+2VypvNrxOfqPzaiWsajyhoyb1ii+uytYq2hxNWm96QTkGm8ViKWyCwW6lWeCsVdx6uo2C3dvpkZ
mdJZC/KchHB+IBqHdBAQb9iDwl/X8d575sEJAlEg8BMLDjR6xuWG8Mviqf/cnnTmx6Cy8T+1aIhc
yq9ewAAUaOy3z7WJcDl5NR4m70Kz2K13g/qe/eJUJheUuYdmDTwvsxibF4UErg2WQVxX1oGSmC1W
P4GUyJ3gWNXfDPOLm1b8lKoWZV9a/u2Xb8a4VoEQZ3k6iBIjzhdL7RVMoYNB7ySvbfHuwqhdBe4q
DAWehiqBgKMGqqxeWKikEc2lUUCa0IkHXAxd42MDaKJ4pW7942Lis785iOmFBNN576DLuBSBZb9O
GAHiqigVWoja+bMaVZH+4DywKSZHhH4DsEMEJqP6Ma3uNkqvKb6UUeqf2VlwiO8DmcmqWgzRwKvi
IKyLOOK2XG8EaMsenWRlPz2CCgK9pML+xPjV0i/iqvylUXQ6FAiiGsEMAxlekdV3PEr5fRGT19V1
Wzx3CJpwoVPmVxbiF3wQn+z+qqWYXZyRV/Ezk/lWWZhZYkxs9nzlQ2oWfzggH/hu+zhlYJHFlU1W
HfuRsGVIo7z63DvrQvVBhZ8PGx10VHkU1knYemwGpRJKCM7oKnbuXQJ6s8+r3BmycRsZw4m+PdXI
guFYrDLqTJBsHXq048XoN0vNOeJ55LWxvOlWNBpdHLvsFkvFFvyTP1OMfbcwUpj/sQLgIA+Nvakb
DrLQDbLowl4HCIT8OEDuC4YRW5se6a2oPgybtZiKIkkqAHnoF7asSLdomzBZKVz2btivSTfQ9W9W
BbTQzAWs5G1TGA8LADndoAdq47niUQtY8+/qTw/Qv1u5QAcdbRCoZ6oumpi13xaHOGbg223/FHFB
Y7iRVWipEoCMFNgYzu9BN9tU8diOpRpVtuAl1HhhUa72qkw7sjrZ32IMLEt5ZWRS9qKkBnvzDGNr
+NcX4TPqI/WH7u6tg58E6ZBZbHTWHRCoUcXeqXWDZ5BNGYM8y60vvbyU6pKYhCw5R2Sv4ZJbB7vY
/jvnsz2vDwqc7HiBrUNRu2IjmWeERcsxE/RsNA5ZGXoAP6egPZM1Cgk9gbAeceYGQWaFwrRln8d4
mpWF2jOgLqPHcrB9r4gn5ovoBYu8U+7XDtKyQ04BXa9wEfZVkJ4r7vIr9ty6XzvMHPtfxbarCYh0
F3Q3+9fU5EIaI2hraJ6qLFxYJDWoc873dj9GAaBdQiwBAnMQzKQJlegMY364KAD3LHGxzwqazaA5
8oZAzLUPx2zwqqse6rhwwM2rCw+4UYTYVY/iy39vrTv++RQtwoWrCfPlm/T8erLvgigPw9ezfyNL
i74CTlrhyEoTmI6WjWoVOHTm7+ZPpXMExDx/zPuXXjc/3oJ3MQKXRSpjfepjec42KSnG/Znkd6hp
TFhOHoXqM6FlI34zaOk14YYZeLGxcogNq2u3lfFIQI2NrJadQzNA9RRdenvEx2XgcG3LwbZpI4s7
H6Axi4Gcuo9M1X18luHFsMq12S08mw97YiWtzVrKIJfrMZvk9++uJLL/vTbjqDSApRdUj7AGevCG
OP8hSoSC1cjin9mM2ni5ItwRdmsIofBMtIaZsuF/nJzoNR9Lgv+t03DTScJ7+mdx1eu+gtYMqi4S
oL8crXtyCgTdSUnyfkid6xthmuODn3VeQmuAOIiJvEZfsmt22Nl26jk+nU4Hirwht7ILeVtDDY0T
WDfbmo8N8NFsoadI4jaLrXCxmT/8NlORPvJxpGGA8MAAw/pjDpihy2pZY7rE8YUssjSGyvMb+N11
kJmJ0pTEaoLA09V9TdxTiWQ2Q78WQYKiUKoGFABsjyvxTjw3E5Yda6XwiCSGcoy4vamWNLnTZ4rV
fP79uZY5S0ywZsLwU2LkV/Hfrx2OhghxgTTgv9bYg+Zv4CQK6vSWuCTzl8VdGT3KmaNVyZ4TYs/f
gupqXX3ETuvjycsgArSWRlZxa1a3ERd454XGqxjPMxzKyBYs01lSiKdlGfhioSHero6CpvZ+ze5d
V7x4D9XM9ORKS+315+UymR7YfkU5SNbgYDzEWrnygV4ranQZStO4+RvgGCgn3YUNldw87FKpykrh
ftRePHviX+RW1PP53IY5jqQ+r8XCPcmK1nMwwtYxZLo8FMhkGD1sBwOJvd5aSo5MdMdJ9Ei4oni3
KBl5kH6ilv6Sgep4WEaPK5QBT7gEXoOwOPURV4j510p/M1fYCSXUsLkwRNY1MFDgevJHMuTa5XZ/
VaG7aS4NzmN6HsxTHib+1GIrnXKy8oijSMnhfvOKONgND+F1e1/fWg9T3cZTGK/mWJ0NfrIljjrF
YnIJS4ikcXr4yLcY9h6flnlBZdpTCVIRfWaiimsoh7cUIZoxr/PwmjI/YoeQL2IlHYDqiBhz89G0
I5CTKrun4I46JHZblVBG3YOXZhQSa+eaBkj3rdGg2ULT7Y5guy28YLlm+geD4MLSO1+tUWKXMMzZ
k9cv9d28JPwQwSTgWHSKx5DP0IFaoTipFOTn+6mOC5x38GpMcmwgxu6cQeTuFos7TyfWJ1z4ncKZ
b8WCcmzJScGU0od0JbzCk9gx8VlHyvsevXuuWDWtg9t/N8t2B2FwgmJHBxYjLRWDfU/iJ+32ovAp
F4iaCZ/DlLtfDjUXlsgI21fbg2kbG8u8dwwhKOHA3gaIDONdweynZekl/Ml+s6vFwDSgVYFHIZb3
g7LQ6bFKzlYqRh3Q/8x/8LpjZU7LT01yYz495HsV1gukcc92qcLRZwhJe7YS2K3p2muwRv/+PEcj
9p/kgBjZYtzyidC0LRI7WywymUFJehq/LJ7+KVqqMbMx77lqowcF3EihZhMWAB6IXolAYMzUvTHB
7Ob3OQpkezYMmUvCw8QC+Ln+kN8CoIcltjdRirsZ2Xcf/fUoeD5K+SH0xYIYD5O57qFjQzbNMsE3
E4CNuy92kO5V5hQZpInKUynkaNF3Mhq/4MOtynBB+lu5GeTdbRzlmNoFHb2Yx3DZcxSM98WwLjvr
10vzHpi+stQY+SM86nn0RJFjQS189nQS7n1/Z+cGfk7Flj2fVZsa27hotRGTG2Vw+Ulb1h7HHXAo
S+zBwmgQKzD9tpcDC2wnyLL3KPPUImMn9XzM+PFDm1EcAc0d+R3QlX8Boz28Y7Vmvo6ZtkZU+dqt
H1fWCsqUx6PCuePZJ8DmomGSbaZzxBpBmPSZxUxG18b9koFW5ZaX0rmZ2DZOy6dsPxrtZTppdDSf
b1A1oXzzM2fB5If3PxQ8TpMhesME3UGyrbNGYtGVUsqVCA8aoruDcLowksquWihrg8awGGFFNxPz
V7SoWvQC4H7+hMkNMvZWFrrvHifZ0FcHA+e5VW/7gV+nvM4RHQNO5JAModPmm/NcHbmqYJgORyc3
q3097Ei1oOW1Uf576ufBuzy8wREXf2Bx8DGGaUV4hBVPc8FtFymgcLe2dvRJWWq+SBLOX+VYvmmw
R2vbXQxu+Ioe/VM4FIdMefgE72rsNBy06joy6LvYp+BrOaMS1pYLBTgkA9iPsZLnxxCiB2NjoxcR
uRZNU1/Owwff/oOXSsblHQjScxFyJiLMRgAhmW8y1pM3f303UmC85l7bOFgx//lTCo0onQS8rQKD
chIh96TcLW1By276bEu9s1NDOE0p60qqUkUOVu8B6C/SQbYS5d8W6aEpdWllluavpGz1vYH9WXBw
UlUuKvUZUUZjOncVqMmmvDUTRNqYYuF+tjRYlBbvKEHqg8PVTJftQ9NtZwuZrEn2/N4kniKodqOC
xaRJAhG8y9QOLSECe8gnqSsRsEvWoVjMSUZ4YpSJyt+EofYgvzHOZjlMhI1ltw96jV4DjktYQhYF
BNx8rOHLabL8suG68Bvt+tL4b8pYTpzdcdJDkjDbDm4dTIoNASBkiOjWZMkS6QIX5cQMqcng3Qq3
LWuuvUKR9Xjdwc3iInnbMNBgcmIQjwaP4Zdyyu3+mOpzLI3PUKmm5MgNZLngjKltIwyezs9aEi3Y
83yoGB+dBcp+tNDv4Wx/dBuWP/ExcgKHvsjxm6eN1HGvtQB1eeKZSEMnwDwEWsJ5XQXvjjY1dFgY
xBPdNFgBVI2iyEKCZyPOLx4mxhYx7J7rRPpo1KUdOdyI4/WCEv3jwRLl3Z5d15iYR6cZAPAkvA8P
2q5ZYM15aa5C64G55FGSPyKuP07Meq7W3qHBIhQVGgpYqPWPZHWB0+LKIIEZxhRXrWUbLoOx9AkD
vc729/BiEsrBZdv9uzj0QIIDDt+NQwqrdoGz+XYgy81PtyDKiKqi7D79jmm9do5GvY/hRaNrwgpP
Ax1aKOKNuNe9jenFmZnlZDmzJ3eb0/4USa4MCEHsDOsEUp77dl9NNkQt2HJM5qNhMUJvUME27G9/
4ooPpGXjlXhYi9IeXyLCrSP607sR0KzSt6nu2Mb4tQBycQ+xp7FpVqvxnQQ81qwbOfzbAJvgWR+k
owd91JzqZbBcfYsD0zGYgJXzgvaCXXu3lAgQFwi34S/mXI35vNknBpePuIVKroE8J1fHt011qrYN
69XHoE0Qm4gAtaWE4m8jMXSf4WF5aySJKwO8lAPDSFAdIEDI8UBM12OVAoXJc5xXzUmLe3aKyLUd
S9kMTmMq9cTTwFD9vOaZ66ndlTOKi0r4HxElWOX4DtKtspV0FCAoO974iCCQJQyG1gL6KtryBdLb
CgEy76z44QcduWPlhPFuj48zR/9ETAyZgt78fW47o6Wv0I+7/0ZKLui+WftcXjrHT+D0cSrdUc94
tOdCk7czTFQ6smEbqAX97KCimbZRF0YDfWeDWB5qtdjjAJgqg6ZEynZWi/9nuk6YzTZfmy5v2AJ7
y/OcVRoInbQrGA/kGGn/EV7H/+TJd0G/nEK7TXYr42lEWA9teL4cc6ebZCwA4ztkMwXIK6d2+XX7
6SMalTqhqbzCGUK97PBqGApXLdX5lbx0vLygGV7GbE5pOnHnzHY0Uhw9JqOSuEq8pBtHiJXaVuef
Qrg5O4qB2WqcGw++88aa1mpAf8XeqpnXEVSxdOnc/hZIQUJrsmi64t++lk8ERJLRwUd+QWUPwOGS
A9rvme6+KeFr5a0bPgKJHN9oP3qf3NLk/aClCoemor0iS7q4PqAH/GlrqdqU5v1f3UU12sTipXZr
IaSFbqfz2JFy7isodFiOl7k8oLLJyuKpvvQ0T3H0ePg0QGR0TvjpDSqPXWh6op05o0S7eusbVFBl
8oElaxVCyvxexGIwSXkkxn3PFjCR1ZzrQC0abVHMDpzmOjLgjifsD3mfIDyF13FoS410LfjrZ70s
C6UExypFYouFbr6doHnDMeogaEOuZ5g1tqlp5l6GSEMqr7JK569YDVHkdBGhyDrT+RWr8tknGuas
CwINyTU42NT825GZ+7qFoW++IagK1JlshePHY4vahKzP0CxAGAGVOUesgDao9ENl1JCWCBDdhznZ
8cNfN83+AWYlnvMfDsix8q2XEh2KIlwz012axRZdb1URaH/0GFqDUZRc7jNXTrkKY2geyx0hcBrz
ZIr90/UZ7smKII/IEh4VsNY0o1uDDE8kc5lNM6bKi4Nk6gAnaqVy7jqzqR/B8qg0rpdDDU4vZOzu
6y6sra2xXf5Y795R2jOTZx50W5gxyeBGqZCv0KEDEgqVFkq7WzpDoCTeb70KZ625wb5Rp2a4CY8T
rTKpI49bYTcg4/KVuciGI/qR4qfvHhD7Z50TVBew7Jz6bF/0rLXx8XlskGYO4bFQ4O3uL497Z9EW
h2nvmE6oTFFj304fyIaBDYN/a7q8zqLx8bOEk4nmr9Co/HhSh9xacUUKglklh/3Quo41U1eCI2cR
BQJ2YrwHPssGGomPmiWZ5CN0C45abeA9JITKyOrfgV/MY1hmAupQBUbeAbslHAF1NIraFR+sCF/v
QGQlgpodJ7qCVLiOm+g/kXfiMpjCwfZIf0tk/xfiFE2RDJjiiOoGhcNsosgTaMsjPcJ06R6d8Vi/
24ztxVYJDW+85AjnZTjtUPsiBbj7jwprPk5Xaz2jcIusRnCUT8PkQqID+2EM9Xlu15+b/JzPxXbZ
ZGVDyQJA+gV8J/vWfOtkjEZzFFYJaZevuv3v3+7mGWXJXFw1u6U/Mw/mhVuVuzJjbTYjA9Pa+NtY
f7wNm9LJIm9JXqxxGr6baF4H/uHsdOG4FRUb6f9O7WS66dumzKihlKolNSpxB6C5jgvxKhv9eUwL
U16yCC8fAKfiKucrLQN5bfVWfjwvFUdK9btBjwGR37EslIYbwYTf9As8Ww94uKMiEOOTVPBNrc8w
gggYOYvp8w64TxAS0H/NQPzrThwu7z8+ctASRPA80bl6OJcXGjuygyQqNn7ibcia4QwNSj7C5szl
Ha16UP8elj+lSHCXKGoUcAOE0ZLL0A9QuHaomRwiKJmCq43oLJ6pH8ED19VA1PI5aHhC0L0Ukzh/
2naODXAZTdqeLiqds5+FJ+KWpmE2HzZHqim0mKjAOMne7LQXR86u5QRLsuIpRMkqlCbj1VGLC4ZW
mhy7dc67qXl/C6t0WWjNoezjc2phjBRHLRptQ+H5LneY2vAXvxjEZER60hHneb5h66pvIvnGUNpK
dN61HZatnNb+3ay0HaBO31Zs29i6P5NboNM08z4FeNSe/3EOhmA/Jc5UuFXzxrT3Su13lVSpurCe
BNd9B+nk1IcDxz9lxvT3BsWXSqpDpsC25qf4Lw1spY6ne+pWbtrcEfrS4A8HGWqwNVQjyKThrb5b
/MuEDerUbGh6Z3DeP2Y047ipXyxJnLH+ZIepN6w0WsuFgi4pyJadlI9PtmDusLgYuhwr3U9QXoey
3DICLjJeQUIwWfncCyRN1UH+EvYnG6n4kvjlWF1907xVEMeCVY+FhxOM/LXlT9SLvFxwj+8El+uW
2ZFYDsl55XlmajA0F0US0qbaEeWEV7LskJR5ROZRCs4c9RaRGbsYTUYN0TBvLV/bDS/FfVcS79QG
0QDC9Ih89hoTLgAENIJ4MO+OJsBhInEo62Ri7HhIOy0uiQGc6L6JThDbcavuf5RbaBupvMafRlij
2nBpHJxWY4MvLmi7kNuTd+7I7CN6nKZvg5tH7CX/XuPkikMrTtCb+qWkDrlF5hCMkI3u56js1BpN
YogHuzTd3ANML/STNir9ILmeQmrPFzhRBlj6KKr66DDSUKEH4Z/n0TsvWcgnD7uoGUADmbQNLejS
c7H3OQ+Syzp3/kOrIgCjP9hKTGzupD4X+0XoshfFDdXCMTGvwxGx2r+yNfaAJj8RnIFg+E5ahtW3
TyyEJ3CT2mhyMg3a3nBJFhEaQd+TC93IZWbVS/57N4bqpoooBaYDKX85DXD+fxJpFHNtbm/XFSGQ
KnUpgv5HjorpXRsJ94KpQVLel65SeZMMJkpYj5rkltQG6R/9rmcei4jtJMwyA++zcltQAkntaz/J
umN31JAG6B74XW9d1rEqyguzpvv3KNOi8bFjUSUHZPxH7KunaRhZMxAGyG5Knj97R1w7hGPvTXr6
sRRKpd3fET08Cb2lkr6BmkziRZsAC/vqgG5HiK1FKmJb3XfrgdByLgodzsaOOZEkjenu1fCH0/gM
fDqsJmIpuLJgkX76m8y3jt0+HVXNxyU+CQCdFcvMZ5Kl6OLTMu6zQBqr/+t2V53E3AJtK080SDsD
VhLT5JPhmPGyRNR6t25t/dYmgJp7LkGqb5j01MrV4gX4l4aHerRHaHD0XJmZSItEElClKNdRO7Ze
pu2zF1eotzqvN/Rha5LLb7nbyD90Si0MQscb7iGrcN2XX5ccxO2nUAbaHnBOzIGi2zpJPDMaEWwO
L8BrwQSbmryUCQ0qYHKImNblmRUhJHM7WjJr43pYL8MfafVDBbEsy9eKSP2VKm+V0q+bPeasi9i2
UPpsh5NF1LbSxcdLJKAbU+Ga+l8fSmDDHJfMSWmyGlrBJZK0dlOppd27SR+ic3ZePYvoTsjiLpRf
e9kiu0qe+Xmv4XzU4xTTDexUNiHC75N6VynuhRyBGWVMr4T0Zh+23rNp9eWu4CW+T3VZ16S/ltqh
m1ypK1nnmD+zipS3DdawOEm+0dAH1tOIp0grp02TIHy0eIuncrKlg8AcEQpoRExoL/KApCaen/dG
CiDsrgoJyv6eY48bqf9x076b5cQseoOZnNwQbhFNMK6hazl+8K4nzbXkC+Pl+HP2AWYZ37z2meEK
/Qh5uUE3siKwMm+3FiKYSrYNGTP+ABLnz4pM+EUexn80qZq0I51vv0LMD+3wxEzCL5e8649Srbuj
YC46j2aUJsKqAzpXtYgwqE3m/to40sR8XA9OP3lSJhAIi0mM6pxsV3GPhne3kJGiKz4k9g6BDMqW
jPmsHjSkwJMT5/o7kBck6Tjgr9nAn8eNGpdmpPN2/fuuoGRrczy7DDhdaDxGP2n4zbvO6axoneMu
hyD3K+UgCwKfu178P8Ym4cPMbv5TT43vKG9oLEmlxQ2A9XWh2AMUhlETLPEtOP1pdDrDWkdPS7xu
oVdkLOiXEE2QgENSyESkCDZZP4WdKQjB18g1MD3UN4r0U3pdaGnAVT7ZwwhLMusCoWxozJDHKlia
wNPv/8rifOAjsxBVdUfNi7wpLYuwC1TemXi1pJo5b6w1Hj9rdFXOzrE0o/ZwfrfmjYZ1CJMAqSyJ
XmMAsQ8wbzEFd1NX8i5fhWqkMtAfdJGf1Iw0u90BwgFoACeEAWfPILPeHjzooj9BEvE1P6CSAEvE
Tip2O7pOfdFwzOmeyrQsHuVcYidnYzgWYiNzswei72FPI5MtE799lgS4laxt2IZuTlaW8P3GJAbo
wPibymmfocTD05v2s1KdZsoZxgOkU1VwVcMiIzm8yN7CniF2WivrMmgt0MUq+5jwlwhsbZd5B0t4
Lc9mp2+c+zJ5jOEi2IOf+Ez2YNmf/IuTVFvrqwmavW+XiNxHj4Of+Prfx5q53FdqBtR8AhKvC7E4
7Fh5HSd4aL0oioNmbyRtIZxJyyhNKJ6H8e2ahBbagXFCBXDTFH9uOKoJ/z0iVlp5osFFzQotR/1U
CeqhaeVzMf/oKN4QZ8q+tERTf1JQpC4n8iUy+59hhZgSh+4gQpr0aNEIDzbNQw57SyXANCULnD5m
TyCeX1Gp6XpgNG0kHYHXI00BST49BoYQ1FxSEAtgWnVXjHXLAEpz+punCs0099F0DQxxEie4cDnY
j1hWEsSEJmrwOmO1+fSFUDAYgfdGSbngHObXfyrPx0iUkbUyQMM789DsjplVJtH0XwDGH8EZzgr7
oGngERvnSiKmX8cyQOTrCAX6oMtW1qQ5k0aQpoY0yOeV0mg1d/c4gL99xsWYVRqvHXYLOLEq6P4I
Lzv2WXCEqSpABQEX6lD3XWUDJT/jAZzFXQ/8VpFdomgxofCvXAlSTSQPsQxwe+Is6lY6E9jEkeSV
45S4Wcyg4v3RFTj6pn7TXKXJfsKns/648Y7FDXr/dZ8ekMdH/8R/3M2EGxXSSqswfrMugZgX/801
CNOeHJpKRpkKYb8sDf5WXpiUhO5RKQF4rImkv004UmyKOTtXkW2/ZcE/tkGXmQkU79Nmq3JMqhmI
s3GV2Cnxwc7eDmdcbovJLrZBrMoU6nPeAnUKd4zKQa0tqnhlYlXxeu//29RYMj/pHgee4feP99v2
Oq5+6QiaR859ex5oSQulWbgbY35WzLIgzVN1d9Kkngm9YG3OpcwanMCbLifFVXYZ15I3RhDiMaZZ
hz01KvTtdHqHKf48kSXrBhUNvoDgdgnsQx/KfX3NgGEeFPoUEnIPsTPZHWgFj19LaKjbC7x66OkQ
to327UcCuo9aTTpocfOee4olaAUDiEQlrdW6TEZ9iVmo/YTrOn/tSWopuTEHC50e5TqapB4RrvAi
U1js60zVgCR7BypKp5AgAT30qfikdE6U88/7dfWjhTCz9KJ4YhkHnhpILMVkJkE/dQenN4ShiR8Q
AB9saKmgw5P0HTyIW6Z2mewMiOpNG+D2DmxUIMxRFFEuUWNYbiwC8eEg2lS+BxR8FqkeGr9WbT5s
X5nO1Rn/enGI1Oj4FIR4rgwe4APCElf24ZD29ub6bH5PVhm668y2ZdR4pwab/V/B1Ihtp9OGfBc/
Z9WUg3CwIg7FW1ifwQCukPkp0MdnHRxyIQ8LOkUTj79E5qO8BEy4Fpe0L8iZUPV+IbB4pk7/lHhO
bniZZV036wNiEj0lpAXajLgKIEmcZzd/dGxwuQhh5XEkenB2y2yDCOpG0y5+1w07RpXThFvIxLNs
7ZzT79xGcVOT8Dr4vV8VRJGldCMRCqQViKu/xyuxfkr5V6xT3EEZh2l3yc+hoc/gUpycYuoHZsAG
JZ1PV608whq44E+tPaMaNiYvKQM7pRNNmLUCpMVCeWzFZ9qBmb0x+u8s9LiF1LQ1utenkuFi24XQ
52lyc9G1cR5E5tbd9dxkT1clLaoCuZU/gJGA7N7l7pJGN3qp592nPNBeBmWa+lJd4i9WIpEDnhv6
MMY+T+jED+lnrO9O+q+9WsF9tl3dnd9qWxopXyI1PaTkgFkBe08bUDJsppFD/aNC1bmTR8oQzcmG
HwXJf/beOyNu3mcnjDb4lePATcyh/KLNURQ0W4XWSbHFmN/UtKDtAYmP4eSbmMgwcaRoTaSnPHm2
QcCMe3uIVQyUWw6wnrqIPXTXnzGhaMOi0pvLTTrWeE/oLg8vL+b/WBVm7jZLLPgq+gKy51L4R1Q2
97OonjA2bsC7qYq6mbJOm+Vr6H/uqAl3EtC2QV9pfYA9H1O9oYqPsYWhM3wJwkFRIHfTkIG7IKv9
RwEMcskid0FBiacvUkGyGvBgaWv8EwOzlyjAL6wJV/5/p8TsquZ7Bj7XZF4JEGy25Ufo9oEo1vEG
8hpEQEShXevN4eKQJTx19jGs19FOSCJXDbwT6cMUAsctB8hFP65Y/FTF1oVOYovhQU3KEBeiKrVS
actVP7yS5J0NAkVStbUjYXraUoaVuCzEKCqvGo3sH2Z2j2sEcf4y+nH/z8SJR8Buje1ESpqurf7/
QRj3qi8jQ8SzA0asCssyLdnuJFZY/QNIxmkpbBCqTrKgBHXJADNpBfzHgk8R0BYhtqpG2U7Uba9/
i54f/6goqWlsXuVb3HbQAlRErsJ5HcIt4TvLim6FQUwskg/BYJK2RPnrDv4d1rKX3bf3AMSYX6GN
+Uy+LRMZ8tf0SuC53FafzWFR0w4hmWpkFGARie+qiuTiq98u9lb9J2thJy3g83s9Ft+JyhgETC/A
qDq3neULTl4UZEOWFzVPfru/Ja2NwKBDusDnDSDsBl2baDi5HEOsC3fcKwbfEOHUvl6QrV1iJZqF
MLT/WHOirzZq+Q7NL+h90+vjLaklxYaGpaLq86zbGPaNXvFzTKTsRwCbkJd3cxw9j2D4ir6kEM9R
UFROesxLgItwgBcHXVpiZ2dYNhrop0Km9ReCUc9igU0vC5j2gysok1qDjs6eM/up/N0zcRCLPo4t
uJPncE6a5eOVM3aB9dBqVkx7kMdqVyPeNSm9L7UFJw1FwrropTch0bVRTRG0xSrA+WGU9HvVXp8V
Eyby/llhFOMAYK0mPzIzCivEwTLO1n1WgtiJY+Hl4pOhWjqYt0IRsgRTx3Jwr0eRU12lfZ4uE5K/
9u8hX+HrTpillFnaRlWMMJZvENNDuukzg/HtHT/QZONvF1CWrCOkUk7YKJPrSj8w6VkRbR/mLDPM
GPYxrqn83rv5N60hOwB/e6b8K2fR2qcPpdh3UR05sPi4gNJI6VtpB3yN8h4kbOGDLoGyZBnECBuj
5vAQ3c5Tk24E9KcL/L+5Xf4aPD7aOXDrtHV+QibfeX2aMVXzNTveRC2TAj0yQgrsTUFmV6HnMjze
St5MS+zpeBc2kcUTVdwEMIXGZeqj9IvQTnUJhxpj5HCQpZfeEI1DcZWCVbzoGa8z8udXuEeBos4v
IUd/hiIfxuQ/E/RDKMtqzdB99t/hftqhVGxvLq7zZmyCf3gG2XQYCFwsZOPJdbBA0xtpyJb4F2IH
vRMPo5QQoD3v/BBDzJQLBZRf8IzmaYVHA+TeeKdAuiglPNd85gVkjo7QdLJvkYKeAiaZgfOMvI7a
ZfYR17q50f+Zgaso7JHVSEJBg5FKqGv58Uz+A9FUCV0dZQWzjB4KhqkRG5N8mVBk/WcKlXOLLPH+
SiEIbrjp7HnciG20AM+7KoOnB4atFlXKB4N6O7oaCKPGHQ8AAp36v/W/VsJyJhXNDJNDyc937F/d
veXSbCK237kBLDsmc2hzuxX+oNf0CdWnMG2bBc43Jp2Q0V4uN7OtJ6JcQxx3/Yz51q4uuxieqNjT
mtw2+A/Y7j25Ddo+TKN81lFq+9DaG0meP2ytfftwhp8yh+DGSNdNIWRgEPKYA531p8tefUlgjdfa
g4RaKmHF1y9yqWSi/jt5jYUQ9YdnUsoOFkPiWhiciQNEWdn6Pk7MpdvSQ+PQgW/NXS9RPhkVBAes
+d9boOeeTaYwAdjTAsJ7YS86+dGBcw1sI5f+A/gIx69nMog9uFDnQVIgJLCQQ37+3JbGLrf/iXfH
3jwkfVVZxWVkeMKkR6pp8bVu+qbGaNwJefWvHmtHKPGcRNtd1Snd3GeAo8pWyh71LLf5oEhu+hV9
NyUkaXlRwnqoXl/nM63j8T65CaPiLdyTDp26lyZzxj8G9qoQEj3L5+aip/AW9UWqh9vX8F12OLM+
PSZK7LwLT7l/j/8Y/OxTEBBhwJWI75klhp1BR27t4okv6wLjwIbt5R1S+qPTnZIYKEPIQ+qQNqdc
VUwxW5XkVq0diC0W+uM4/AMDcTiN4R7Xc1a8g2gkyRJczLB0dylLDCCH+V6myKxG6ryWYv2NRD4t
tUr0WaHcIBminDszilgN3I0/af5tu0PzFAyylBenMUC15ifIwyn6kO6mXmzD+WAfPcujMhDW7jbn
NIaVPg7kjBEAQDrrhBof2I3FoeVagoOI0PISx29cvB6i36rbsVNEMpUbm3dzCE8PXWu+wciu1PnC
N2b2pEmZAllR4GAaCebtUYvSkYJ8yKCyuQJMYdgT4ZWvRTrTFQ0ub+R458KfiW1uaiS7rEyiZcyD
NDI+yjWzhiB3RqpOOaUbWda+CaCcREcwRA2N23YIiuvUQy17sHvsBaCG6onK3a93g0u+srUXSnXy
RK1UKVAmNkIAJ7abSDhuGxjL6HODZ0nB6dPV2IsbQVBG5E3+ClXRn0PvhxAd9pWMugXday5jOWXj
c6DOWy3pxS5704+J9Pw09wbfykGAYunT8o/MZkBflCzhKKsnllKHsndW95bvqxjY7h1qD3GDjJ+d
99UxqWKp9DdxAriPoq6095i9LQXEp1vGf+5VQmY75MgBuGZWYnHyVHE4L6dTFaJKdzq83SEzJMDA
Oj0YVHF/6ui8iRxsTfdX4SaRTWcxMVNF0xE5fn+j7XG5Er5BGshS9y6gWXzT6s3cszTgVu+y6rth
BOKo/zPNAHfc0RrnWrjKy0tD9IwQ9Fhnvy5u7u22d371AFbNFWIP7JeqnMkv6QmGyvbCrDRbzQ+f
e/NRGNaashajBNWOfJuFp5AQM2WklD3ND/W56UuFLcKvbNli2vHeqG+5p/8jBIdKrzvQzolsiHtc
TCJo9yWTytoeUMrRQxdHbLHUPyZ1OFCYPxMAU/eX/FXw28oZTs7wNVcmB/zJqIQqEiAX+zU9LG+A
p7dEfV0rFXblMAUd8E9cMDJhfgffy1+UdNb6kqRmAZvmd2KHuZrfSpIb/Rhg2J4koudfWS73Bb5c
Kym9emXhmhqOdSCc7w7HM42CiXw6mF88NK3XDHoATNIiz+gYfWUr4LucPIBDgQvLP7NIT34IBG/z
yp7L2jyEbwjSPfJSQrz2t6arbqfD6b9MeDd3BGfFPw683FRGqi7/Ip03OEvy5n9YrVxF1rK9SsyF
/12cy630KtzboV5/opZ1pBN2JPR2eRv7lWQ3zvNK72/8WUVrqybGeTEIMLLUWs2fUlD7Ur2dA/Xc
DlRxXDy644giI7Gs/x8D1MbiSrsxk5c4UgUGEPqwiNuL2CnvZPu8RsUSh0QVADIwvVMGgm/Rv1Ji
Ox2cFEDSzXt2sYQSFkmx0SpjVe3piWa6TYOkG+MCXUQ+5sHqMjUDAcihW4tzRtDSBw9PG+NBfXx3
J3QmHO0KkVMVfbJIZxBchauGlZ6KBDVCWbTYBPcrY1qdMvQMG3i/cg9yYSJIWVFmY940qxaDfcrG
HmFrff4TleAb9Ha6PApWWVieebWeQx0TfbTWSMcyL2SHQlTHxeUtd7HJ1M2dO3fpw3CNqktR34nE
LL6MnLsvV9MrOiOvx3v0Fdyw4R6T9Mch6SfWIT7xfYmjA96qRIKCuTfpMQKIl9JQ7ayZErbKFbrA
XPNdOhXaPKx3tgiNGWOjyR13UW5Km8V3qaX66BZmOk7wCh7RU9mjhp/LVU45iPt2oQNV6BtRR/Uc
o58C68O63XSzDZvqF/e0BBTkmLChDVcvCIIRl6QcgCeEAO+Drpyci91XXsI6WuwM8Y46o1yyEqhO
Q44HdMMFcsaamM5pDcM25G3Y9fBceKEGNIiHu2yd1x6vwVvNntnzSnk+/a5WRZ/+mDjfVm5GyE6B
coxhKqD0/n8sv2/t31om0gzPeoxM7n8UdBKWEv+57CoRwKS/3xM18SX/ZvojniAfRHrNJ4hQfpS3
O+/038kQfNw+ha3YZLgEWYbQtcHkzO90CdJuwLZnoIZoEY4STGxsRGf4klzeL7hY94KPJ5iovGb4
H8d9lUDWvIH1ct23DLkKdmRIKv9fkoj+9l27YrgCCU2WiExZ4WWatzH2v6ErdX6WQdgeh3TBoWQW
wFosE/0uSSssbSid83nHSydh/77N4xPgEY1haiSyjILGD/08ROdoNnfHbKXmcParC0dNWpxbXtg9
c3DKMxG/BeQQqa89dAgFrXBfKkNB0YnmtQPoX2e22RgoOui5KwNQ88BwWCE/S4VnpqjfB1Qq727f
t73/Nuz+z6Lk0kSe7rWsdQDSGs53mCuXFxWMvFbINhTXz7NVbMMp/P5HKxrt/EbU9wD7qUKjTOOr
RlXq+3XUctRQBa6s9P7jfpM7vCFUia4zh2XH5Cb7h44ExoACspt5mMQ73cLLmhuVu3/SIrJHqSHf
63bwko7DTLgJ/YKWKL4Fok+nLUzUY2BXrbxFGr4zXQap236VJLGQxcT1kpsQ6I4JcywBbw1MooTA
MHUcd6+YQb+tkctVKWwBN3EpWhMIQrjzz7qaW6alb2MxjrDSYmAc+kcHij9zh+lGCLUC1CWvjB5E
8It2WPZy28IP14cHFBvUlRfuNYOfdaeReZgtx8aIcKzkPTsxwJc7jRtAx1uERR6j4prRcJGWx2ya
aVy432Fd4eqyIRARLM9n2q/AljE9UrEUcrm2QBdIdPZbGwZtF7EqbNNaRlA6U9pTi4V2MUHT9lWi
mdh+zB+qGAWd/cF96jpSGfefCsP5PanqO1DpyYsjrP3HQsDVTGPdx2Xw2RhPqaRZBj+p5WUtROjF
XmvAlWQDnXLDhXsbnJMWPikOsPNj+63XhbRHoEULzngP1pLiSvl22+6c0qRFVs7IRNPHr8B0auHa
C7P6XmTwJZLgOBGkEa6L51GqUTrGCNZ/mVfJQv3DQJK9LwtGxy1FQNdTllm9v5OLNGTHEd5Tx6AO
eYHGkjx0wmE9KrgTGmIWJOg0grEuf2GzPImO4dtcdaT3SUVt9KKkyv32sTp0XWS987JcfGYGogt+
LFDdoHH1gyUk70wQu+tgJ/GaGI2tndE/uihsNKYjyrOV+4M0vma1S3p+XAdHirGLgQ2heA5miVaZ
L775VhyN0mi0TtF1jUjFNCHhHZiLmBupMibxR7ZRSlQ0In71qkWBDSJB8ylebqVgCiv9/34fnbeK
dqYsY8wSg9Mb6+nxDOFR7oDWeq35R+Ll4ad+Z8giytPvlt01wr5maiIEmZuVR0anvcW/EcgmH8qt
GsvntAJzTFUY9HwFkFtFUqBtvxqBKv8jY+9XQQLTTIM9AlMji/KiAQuxv8HAOMRh5vAIoyucOb/u
601s0JdXrSmhdguQgZsiHuVv6tfK7HU0LA7mUMX28aNKQJIaq1vcZHm5MZ1jIFzDICe7modfkQug
0Pi1C2/40aMtBlzVL+NYIy7Eja+LVZi4W23qMvzzFonTQWH+mnRqCwhmp25+vEboC8luFj8P2Gjd
u1Wc2k4eUFWC73N+PsFOApdD9Gcl/YA3ToGt1PWV0B6MLCkmRIqyZrHoxLond3mD60lD+U1W16Ek
kwsGlBv82f2588tN3NdYLvmhFc8j+weR1iK238KaEbdh5CpqIW+Wsbhc6xbDSytKol/iAuajHv5P
8ou8rzZT/U09oWJjWGwD5NLFPbYsG3+hieXjnv+EygL+Lm/6hyiz3qxwLQwl7YMALU1NOuJjQEqd
sKVGl5fvYGdQie79k2xEwGayqcWWqZgOcgerp//JO5hYEhppCOWFx1zFmgs2riZM9mqjVeRt29QV
zQIgLlWqZ2BZAgfkJ6QwGPip7k9TdGXVu5d3ijRSowobrrAOVUIfx4u4b7d0gPisrXElWYTRavdd
Y/v0tt/ARrDuSIqZpkpARffQ6qybXJ3+JckimOf6P4ovzEKMmtCw7tH3fpHRfPftKhpZnWyryBNx
a3rzl+MZV/3U0Z3uZXxNe2GQgYcYu4skcq8rn09hxAAdSx07P2h6cJtdQRhXiZBCXWUIDFz+32au
G9bxDf5hLb0phUHbL48T0ajRcNuBgEMQJ8khIfh3/gSd5iVnLKyq2/9KJu5Vqhe12fxj9B3d/ctf
fJPypSN+IvcBH8lvWyfqQxYikZgbiILYtVCc6ZxZnFeEOhD8bj+v4CiYNoZSHHT7o3kCkm+fOLFX
Tq4HqtrzEtSboMldw57b68rZGoesSQvByXGTYLpAHyDgzuQgIi17ZdHooDGWw7Z9eQSyMxYSh3L2
jESSIMoLqWaZ8lkhYnNWIKL73X9d7E7xgxjvuw5lb10/JO6KA4/dOSlGK+pl5PO+ywQqInsoBzpV
3mFCA192lyrzqy1dOWPkwKiqR9/oWfpOGIDoFKFNAYicIKZv+RjHHMST1QPgx6Ic1xIrxcQZ7znP
30sR2lB0HVtRPUveUsyIPSp3ubjv2q8udzA2JG//+UD3Fb55xHBtUQmFzh5bpckA+OZh8lW0eHld
+KPJNTuo035yaYHS+BijSP4N1/ei3W9o3Rd+hMGZqYZBvWWRtl7eXMG7wIllO8I98pqEl7D+Cqxl
QdgygMzPhYDQqI2grMxEccwq9CW1UkpWshgzAoeG0hS9Z9igcv9M6L9gdOMS7d5rv82f1VvMBdtO
V3CLN4rU/0VsUKFvKms4wBIeHEsN4lIghSmAbL4xf8iw7A0s98v+jDuvOR5+8fzBJHfupm8+3eRy
qeCvOr8frAOVm/vRs9O+vQEt28T1rlk8M4TpP8ZEUCYhfzwKU3qTyLGQmzhajFhGjagOx5bKYnb/
L97B4gvndqMR6OhFauiCvdO+uPhqjG6KgdATJ4+wsyHlGc4xdCBxuV6JbBAI4ulF2XVJrG4QzFB6
yM/A9hC4XYkMbem8OC207i7gd1eZ3YHWjVyrPYy5F4S/B2z67lEXrt62CuTOyPtPap1/jJY64Etx
IQGvWydtuJTCT6ZGufyVFmjT6oYib/xreqp5hIGB9AzRHyO7FJUOlOZhdxph0Pc2DTmdbovQ7hkv
vXxd5TkS0lWAmHJ1e7PnEEveKsJRf2K9j4Ne1L8VHSpbocFTbuTtx1WSQVBWnAl8PE2HRIMsNKrG
wC6FruVMXruGvS9UEuNihMRCQswg1yoC2JLq/sBul/skrpA35Vt5MQEii8xenzYlANoSGek/gWwd
xI0OSPsa04iGc5EwqsaWPA8X7z8IiarqAGPtBBgdMJYSSj5IIYUXYiJqKVD3yaG7D795vx9BrOy+
OxSw9JA1sc3Mdws9sLRKZOEjRHtvyx6gIf78Bp3/6rzUbg5WBHpDkWi5l9/mIxhbwT6421OhLzW/
BQoH+idVLI7G6yNQTOuzxKX9qH88wS0jWyd8osIB/3F0etuPFXA9Q6FasEdxQdewqYY6bRomrRiG
QjanHJZxdseKjeJ96ktmHd0TDJVKJNAe/Oui1J//5mA3ci2iT7HM577ZMTWWB4kzNPLwiyRtE2DT
GkUXG9+MvumYV2jqL9JI6dI9x56nUHsb5ocIIBQwlam4WlvglyOjQIlgpHLUpL5lWBpwOymnSDTE
PueQg94/lINewgRmKLTkmIWxozWd9aHVi26oWlm/VcmY/1EAbSYqQCtdH3tHTu6AgSePBOMN2URR
sZCoYykdGpwK2DYwTbvu8ay8VpkL0YSBC0WwTsgACXzeOXaIhknZNooJHmGUN0R7HMepwoQmQBPE
uxepRD/bacE1QXNaQNqLRX7BsMySKA/pMdhm/3EsI/k7xxKb4pW09Gy0rVTJfPP8b5MTdDJB5/tN
AkTuBjrqk0xaixX/MmL4FRYQsd60MDsDUTPOJOLjd7ure3/mZh0b+/O8lOboFvWUC3KFQxDi04YV
ElGFJXH/kK1uUYCgNx9tjdEiuDVAt6TAA3LWSWcisbfc+1fpJ0sh+/hVBAoL5PIJw1cNggrYFBsx
ReAyVX8O74R1rRH3LHEf8K4uAJA5LIaQ0erIjucujhHcq1cEwZqKc1VUXiwrW4cX6LjLQodRtOtu
mjcgiYpxtGhY+jYJFKG1WwBPw+N9AIF8KG2naGRM5p8dpk0ulZSYMT9AtMMRH+eN0Rq2LcwSBHXy
KSPZj5sJUPVSD9HGRmIcwRB3Fk+cfXsTreZREPuTeaXhjqGKNXSZmyyjbdwg8tr1bdq14Ju5syBx
lONsYZBAcPeFzPtwQBy/GMA2B0x6HmU/Al3Jwd6Vp/3ZH2tquuYw5a/ZJZfLvRiUKhH2j9A7RkFF
/YTt39z+cpbr0eMKvd5sg+IrtkpUrDBjG2KyWHDrYOdv7qfE01EeRyR+nGIsGJMV/3MAc8cjxD3H
MNqf5PO8v4LM2+gMG9eokDGKzPgTSJqiOeKelF+QnxXxJmsIFB+RrYGGSt1VrNP+/2axP3rTtzs4
tMqsJ0e6vTKZ8kyzxMiallGZN+xKkGnVv4gZcC7BE3yjb30n3GzZw8vWs0D+WJ4oLqebren/tVQn
djspXxRA5Q1KiYLvq10ISBndZrL8+8f4NTUZ6F8Xg0c7q5O4jYukYdGExUuexo81tv9X4vyq5k46
Gfr5F+28Ls91bHKN8G1u9GGd4U2JxNV5HvuSobnJtldEodaMChhZJZ3ySVVXKwyKPy5Pm+Hz/gN6
eCXjfXrvpZlt6/gj7e3Ax7lFHdURsj/eyJPbMk3ogHS/2ZuwdmOsvhhwtaVW/jVbNyMJJesFcUhM
FIYA4wcMgz21OfNdVLxkBYAOUpIOd0T36HvIjCkfP5sJxJOdbqPzBICDpovsAT7GAbJhctb0ZdrB
4zTXANeKqIYYL+4tCVgUUFKS4lrt90s5W3Yv7W8OXIiAiZPcFznZEp7y0Ks3OqV40Tjqscy6TNaJ
U2ziZjuFNCIBGcq/ITdMSxRMSzM5jTbjs/2gqpUbfQmnqPr5lXceVGwYQtZZJFVtNqnbvVdpzV0h
vCiLyiIDWQzhFhxbiqCK2k8NwftdMVrGLAaxECdJiPjJl2apoMU3+2zDXiu3fsuTm8PXgil2TuTZ
0Gmzy6OlCHkFRf5rejF/97O5D6juL01ezJSPUUl7zTnzPoQ01fsqa9JPg5H1Eyg49CtHGnvn7xD3
vH7MKQUIBLKbRcUN4Khoi/QJJIV+l6KqzF00B3YpEl2y11AxCDg9vjpGqyYV0Mae7/HJ3sE58b9D
Y7RX3Uyg0Pt83RWLzwblR1TsgFFty2J6/m/7WXf7BczDP/Pp5pBeXyTHiOwJYfhRWNOimoNQ7R8a
lTExDPc/wLoYr1GTVMRI4SoX8lmXv0s4hWAR+Al91omtMWV6jLdO8L63EyozqvaSFDgcki50ySps
YLnaogjORox4f9diim5GH5E/+O3fB+ZlyFWS1mp899U2tDbZVPhDmByZMIrE8oCDoIMSkpjVW8LB
Hbo4lORmj5qMPPbf8PkQouAdVwHr1kJ9amhSx+8NTH/kqfwtpE6ttQ9SL3S/31ZxdMO+0YaD2SPs
QTv4ybuSyT4uwI+6LKnIGTvkPnB8sQlXS/HwjoNy/Ksq5qF6sAYSuIEHAeItmGQwzZ3vbljTGFl4
PMFXaSl0JFLNfVF649mtKaVxLItS80doLPqPX3mSLtPmlx3MImyMCZUCi07L7ma2s4s9hXEUmPk/
GCKqbmk5F5B6goaOHKPoZVOX1CL5tLtZ1+1mZpGQXHxEVlQSaOaak8boe1t1dbyxs1AEkYJnzTdo
D9FF0q7AjAmadn9JtVcVftQEgCgB5zAJkSoRiFqWeX4areM8RCorm5BTzJDV3enbIlWmhsh8Z3wu
XQ+EjxBPUFf7lOHI+KrylUJjtsMkoef1KWxgLB4nkSSFOhtIJuuDvYVYfAKqNKeWVcUrj0tQG+W6
ujAZGidQPk/HM1G4/7gD53W+eDyF27IORe1wDhjAF4vSPfl8OrsWwVgho4qO+2T7qI9EYvAWN1ud
9DyRuuAttvKTz2olIhuLQviiYSq3rr6/GTdPlfP0S4N6uTyMszkdwDvsUqiDJH7w8ctdgfdfqfde
FXs2u3elZvsMHw9EDFd5QQdHl101O+oCEiVN/BNrFXY4BY7SOfFfFXdPDmdND41FUEMdQEdpfXlE
oFaQcboeoHzHEwSQKVcl+21BFWW9um2tXxwZotOdU7qLJUf5cbREDsktEq/Ak3/DFsuydkOyWb5K
nEo7XKXTNIRTQFrhCPRiQwrzqS5oA5dAGfOvpCJEQWBUQG3J7vDv+C6x+hpWEDpz3pato0idS7a0
gDjCoyliG7ge+lERRJc8Z85eWVUNswL2TDRavZadSDkzozn2eQntaYEMyGKvMJnug9lkT0hT/XhP
T4zP8Dyb1W5pVxTw5vcsGE/8WzOfSinrdBX6HetksFGNT0rSMCRlX2k9TlEj+K80O5UX1/0LpRzC
yx6uxHdp5Fd1yd8LyCFfS/NP1v8rgKPuDRUUejgKmG48LZ1k9KvOtBF/kGw9iUre/S9l/DixiPRS
cQrcr0NFEgy79LuOzvkOwK+D+DdXN1wd0M6355Bh4yqDZgkmtHlOl9II0/nedT4r+94cLvLK1iJb
lI6vhvC7ZAvYv1s/vuwkmi7P3th+gTzCEWhICE8GvGHDIW+xges7ENmn5BetWbKGGpMf8XN8AlEH
mRoCwWIF/v9PQZ6KawtgwDqYu5QH4uqAEHI6H47n00tkVcougAYkNx6wVxYil42ho9fWV7STekNG
JXc3dCo7KYvZrJ71wgK8UI02ob7Je4JPQ+f+0+SjaezcUIyiyjRKJnQRM8aWZtV7y8AipvLt2wv5
yvtL/ttbNFAM12IcyFYnYCqTOmO6JoEVjlLQ16ra2y+XHqIqyZUR1oeimrj+7EzbZMkYbqay+isV
Oiv1/ltpfRVROB/F+6doQE/7CuOiu/QGJPMN1aWv6I1N0hX7fU0gK5lm0rtWudGBYMhfyqT4VUaw
RAqNbmouB/CmxH7teNAX0lbh7TCSaA8NQxcRCPPZF3qUjtFJnRlgGEZc26SfkTKXiCeYMGfrIywy
AL8NtF2H6+KRpB0mNT1wgu+4KgX3r0TEdvoO60wA0Qv6ZeFucAE0KADPFBg2Q2b63quNjXYNeu3M
GMe4fYn+2+nXS7LLALyKXxZlFTA9gfKyN0logCoGxi3FGphNwZT8NlPvxBUjL496nbGRU4W+o/wt
Ib/4leUG//ye2VhRDd3cFT2UWnPEQffw5NBystJZee6KTidMpGdrAaR4NEXZNGoN1ED849MquOVt
Ndf4U1u8IAYSaxYvk7WUmfT/oexzJ9n5oyWg2+h7TzVa3VplXV+saIer/XGp4iubIp9oh3nqD7Jn
2+ai4kMP79gk9WsShTb1dCwxHBS5vJrDVdUSiFrjRsInv8UHyCdpvB0CrHZRD6YhswE7KjGh4cdg
R7J4ZK2TS/f5yKh8hzowXQu2IcvRDTOtDkko4/CoII/ZQRCjQz2tj8UGPn9G4ZHPbbvfemCADUSd
SphQKQp/UvnXPB7LE9zWU6iOZj6W9PURe07TqDF+5dtd6spq3GthtG7RDHZmhNq7Vb6YeU714+A8
Q3/EOVe/rUOQf4RztJuADIDVnBKEAQqfQUlWyzUnRZFkJK94seyB9R6/mGIFNJQgESNnLqb27eyp
HA6exZiws3YcXUMmBIkE6xxmeLpliPLSfACPZZoo7+ImArgOIpCi8OWutpKmkEXH8wobc5tmSLZU
StoRKSxD1BBDAeCSR09hm1fiK34hxUqjVYgqT+kfVknN6b77bC0YQ0p3tbvHgufqP7ZV7DGRb59b
hhWpgPNUnBKIxIbJnmbWZHuhGVKUQuRLy/j8g1Ar+GDmJJVZMPtlBYVLDxgslafFFwGu+H9+MnmQ
XL6bCHPirfXxHyPKGxwq4YvpIbu7YhC9vrje402StxKOpGXqXG6JMCEZ94inuyU2HtdNODeupayi
u+i7NYXVXViiTo7KAGaGw8nbpLO38Z9XcoBy/Bto0WMJ6ipoBJPlJFqAEacgQyPjeNd7m8JEu5uE
VZVHqEslHARmoYiCq4/c5no4x8bePr68QpJW6CcdkF7GpEi69gyVtqw75gSUnGrik0ZmwA9WKLag
jTFDa2NWq/WfpSBItWgYh1+2ZviJCUzyGD9a9YB1Q1rVo61aed2ZO6JPXqmMKCPVmeQg/X1eyzYR
3Vi7brlu3ua23DDhXJUOHbawCLSmsjqH/dLo0mTaSrzpGqCAIjipH43/+uIHCgpFJAzp0TKZNQSX
hhNIRP+u1gvt+/oRYho8g16UPHJY2E6tGu22nHAnK7TvXlfJjumKAE4zR/GRQqp4AjMmwUSMrvN1
RQ7ibZrJIuHe6x7z+xq96BsnjP5xMPSPNHi76Y3rwOA80RFPKXSc0oeQH2MLLKYgU9TvvoGTADjI
+iVF+CxsOF4iGTzzTXaRt2Wpc+NsWasC/wH212yT2OzrIVG3eVwYV4Kc0vThGxEXISeq7N+VqrzO
rC+60kyhyUq9NqJ9YYLfxV2EK0iA8sq6g4AeU1wF4akRT+pdb5tGzqv6ujbkqh33OjWsR7MJL7Ij
x6JF/dH4+0SMo6Q92B65hSn4Qdi8R0fgz7LLWoldpnkKtn7wAFu3Zav4q407x0zIaP+A/gpd/pFg
67aVQZrz9UDDmeIgd19hF84VKmSmBPv64MMWAMWbZlvK/iVMBcgP52l6YO263vAFHVV+dFLMqHyz
bs2aRk4rLJcs0/3Ag2TdaSeol/q6FDosnwQ3bX05KIL77eM9ZeshnftyWVRC0HgpSlqDT5tw3SwL
0fDdDOYNcEGyG0dKaZoM7d1vqJLiKP5mVmkJqlVqAmHV6biUlhHn4AuSxu7461lFgvYNX2632piG
GZaiqTuudgGLJ6UCxf45m3Bs3C0BNW/iAMhdgzZQ6UcF3EfsKml6s9ajMJSdhMQtYyi/kuplWmnj
GfDsmNl/QRiZmvmRs8PVngpaC+yK25Txw6QcUhLHFfjRkjVocQYr8sH2MU9mr6ktbay8Hu0gnntB
pjw14FWiVgJL6lkhQiOK5+xNNGGH8GvE7LD7rmpgeO10ZJ2vHEC8ww9xzirz+ea8H8tc3zKSRpyH
t4fUThtR+92kBHH40t0fseb1RT2mFcIT7cLvt/6poiJbEuZu8cDUVSFupACsg7Lq4rk8o79UtBvl
0kXonL3YcmliqfnHlk/BPlNAptKOhcwl3rkflzAL8ughK8Aguaurg7jYBsQ4rVGEc9ea1kTZQcVJ
u0zd7c76cP8CqYbDx6e6nXZwdESkphc2FNjhLJygIfdOlkfk4xzOZ6mQMNpc400yXCUa2kjAKPK9
3jDuSY23A4oVwcbuQ60OMLjd+z/VK+FqZBSQeV139OJXv7UIIat8xoaxyKNfaNZESFWZ/5qH709+
4QSh6jP9eac4pBxf470uyYIZ6DPKoR1i1GtGgGgpZV9FeDH5MtsDQk3ng3E9u57uXZ7mg5jDMOjV
7YvSliVNQrpNxM/YfLO51ugHODc/jp91G82q87ldu/XdJ5rw+I3d9L6cQXAdhAysI5uZS5CKuCxV
ukkwqQjnVrvxSeMGyjUOl/+iIr50Lz9rnSJ8VpBjjDzv8NKKDBLK/E5Z70wNepTwBv+bQeJ+3Kws
6Dt+Cj/4XkBukkUtNLWZQuOHsWsVP1r5OLtWkDvtMv2HxvOLKEtQ4Y8FkKZSmCeyk9kkll8OhPAt
4y7SRE7HfeVbeM75xELYdSYXajK4yCX+k8xNc0y0ZztQoMTTCMXujgXv+NHMR+4Su4MuUJv1+pBk
sAK4TL2/fFNYApXzIYr7uCMtPuUGfYOhk4AiAvYuuRQ1i4Ez81QEpdYFS4ysyXOiY2U1UiUq2AT4
v2lpVstDPnzSyrQqJsaYld/trAA99ejJE40/kDFH5VwhDY27lmlZaWyuhFvUr84oe3oYJgj7iY8q
io5r7cxvwpT4laRIH9ypVvNRi2TBRmiT1mZV92XqIHza4mtOD9x0RaNGhAnegT4XVXjFpehktJcr
gINb0m7/FFhVwBNyS69za+IBaEzpVbLUpTlaa/RIvsIFwxv/zRrlLdapdNazOnPRXeA0QgtLhz2U
SkFJTH8QaDUp+Z+RE1X9q1QTO2VfSrNbWZHpATXlmNyRDwdWljLdVqnUtuqybfioSks4T5mG5+B3
V0pLt98tElgbFt104TLqOYByiTBiCdaW6waHCVWOZ+k8mDTSdqeG/tmHujIkHw7nB1vw3q/1z9Qu
4J3VdC5Ze4E305We+S+WfXA2Lh2bszXiKM9WeFgWbv6yqihY82XiFb/f94I5enSIVDgg9W0gk7m0
t3CRg+3NldlUW0/7LGDz0EJb4ASU2oDy+u2ONDNzZWuKOIeT3w7/juz33nZ/TDOCYOofwasudlXM
8AQcFfDYigIxka2XLd8nhRexZioXX7NstXPzHqPTWzXp5ucAkf8WkbFgxibJr7XkvCeR1K821hsp
NJVoHYyEZuRWirWEURYCbzLfjx8Wl8TKad0dcfmr3TzfKVaa/HLrwh/wD2Lt6E7K6FgGSLmmdeyw
w77zfiBd9xSpq9t3Tah2+QetQMuGeFcyRTYLCgAp/ihqaysoy/J2cCkDgeEdZPKk93ePEZKC90xP
BXdutXmQ4LQtyradYj/vAH624v5SJoLJCJVX8YnzDKYnNFF2ZlNdgTlCJoElzxWsK5fLDb21Il7v
jXbRpInkg/NuJItHKZkkqMMQ6Rn3Bp5SsalFp/0yMwQEzKSh+wINByXht1724ZAC+dYrzQ/W0hMp
hhaaJwmWcEpaDEjSF3ypYcsuuB6ZMlhtLUdX5YictzcHeS2oDPRSYgJ4xxcg4mr2DfXUIcWgvwY7
KCLXxqNw4CfKEGXjtiInIEpUpBf3ijoIpCRrqwYNgsEsU83Yjb+IdPeK1Gh3hNhEDgG+Ibeq9Xx7
xt3/bebNRiZPyWl6so0RqZ1TZbSfuAOuCPTbOF8C/6lTu24of+ppoobvkdenk08Hx9oTZwQgEsjn
mkLZO2G+V+u/SxO/vcPnA8Hsc1VzTQy5f+UkjnQPwUGXlQ1ONJkdfXNnF8rXOeTz4c8gWC/F21Iu
pwj1azhXNEzzsnIxHVImbboFJVUX1djKrZk9XhzMmfFXErqp70yd0z+tBcpmVTeYTfuaKgz6iAwu
DnbRlWlP3uA5ml10VageNbJ/7dZuw4Hn435jobw/gQHnubzbL/s+gnYheO6C8XPGILDePUrM8YC1
3H/2KR8ChQCUtigY8+Vwt8gIa5DmhqhS4xf8O63TxUDEOYArUX7gZsZgJ/Q8UH1sf3m8KO7gAy+5
3uYHTg8pYGt0wBFOlHzpkVoIUf9ZFqomHhyrGPKwbaNZrCJ4J/Y4C0djCkPn4aD9dafJzIyRm7iq
Has8ZQ41mr9ZJzK2PO0FsRKw3Cd3hVXXXEiLNAAVjhog1pYSfopJNcZ4U94wBBNwKC7cqj6LzEoh
bcl+dTfmQWDpyuRzRsurP/XRfaXdt8Vj03RABkL/gsxpaGPdYZJYRRZrHzp7MZnduwD6lzYWz5q0
cN+ev0WQ5MgabQS73td+19mmaOosLBpg27Y7A69VAW/GoaDw9j3bKb0HzBpM0UWeEZVyZjD+xHs5
K1nND0eW4tlHAjAA4FPUgQtpjZKn2b3yIFm99ReGR6YblbsCKXewR0Q3klocUkuco29rkCNLaKXY
TN/Wzi20c08ovHrbDo5OrfYJctSF/i5EYUsrPqb7sp07LHrm1MyA/d9ajCVcymVTktklD4sE6f2B
vYGQPVglo+9b402ozkadOcqtw06diIP2SvkhmFWcDg0noxiX9fePFC0F1wvKtlBtIwV3TiWgg7lM
C1SfsS14OlWpY13anZ+Tq+Gg8NLL8yYjLaCckNKcoHUtGJSQ+1Nt0GE34v5AiRPXcX8gYKPgjF4y
I67hcEZ3k+15/J46ggyC9U/yAaQlQQUI8QtEHL250DTMrIENYGgWE2YBLGTMfNSdr63Z5/GfWvP0
6p4q+hDOrIggYFFSkQ2tcj/NDXH7Bm5ouOQzRbCY7hxv4SFLwDv0nxwKJDDLz1tMtPGSUMaD0KVJ
XTRSwQM9BNAxhYhZOu/j3z6thRxArM86b/m4sWOtkZMoYkMLLJzmQgSsEKGLI1HT3gDIwVCH79XV
p6zffZvkD+f2nm+m4Q5q7R2auaChLkeIR7koVmURU9KUpL1Lx8R6bBssY+1RhMxOmLLhEzC5N2Ra
K9TD4y70G3943GIh/j61hBqDV1nZIFOX8yyaQsaNju6ZOwpN0FG+LXd1hLwWzJwF/m4MkwPXM1bb
n6a/Fz4mtGdRDy9VcWTcUtznxQ107BS12O9pD72woQNjfYdPDGpxqqlUX7ZzInsLXFUxC014LnIG
ZoDyU6tcR5jmuam4kmLiKi74QzDgBpRrkkrtS+/E1CjoHq1k7zQ4BL6CZtaABQgektEixfPPdjep
Y+2IzPXxbMAzl3Kga/MoOlgcN2MhOJmYZR+99DGJwcMRWAiBXLY+RT7Kc5BFA4lIYavS5FBDcZEp
FkKC15PbV1a2V6uWSWNHepkm8Iv71VfeRuGbwAfpgtcmT7a3TeHHmJl2HZxUtzfmSUK6pr8vHnJD
sUsyF1M8TAnoNOQy+kDNAohFLo4PNhBVwD2KjUnuzg7FqQpCbtGVgmRBIX7lkIQ61XNMctEVP05l
ubcxlS73QYixfIF4BTMeb9ALJvY7f2ffVZdzd0zJJKiiOA8j8MB4f8zdyjItyH/y32T2m1yFEu5n
nd3xvO/5LGm6sJavL9oLBKPSBPWHA8+iF+4hudzQAYNgBcYLAHvTc8ulrJ4l/JkMmn5SudEt27L3
QebUj9A5u2VjP9tsnV8+Czt5hARqy8OPJS+Rg82uhv0xw/eTS7YURfsLLg4c6v88S5/3lGB8Tz8X
F8KoHuY1OxsEA72cSY1p/ImkYDL/JNNwa5maC+ZToE10d84pEkwDLfKE+Tmk1RGve5SZTXb92KNS
P4jR7y32qZnbkNmYYoSYD2xucg7EvQn6OoFCfkzP7ynlxvYDhPwbq9s0ijza6ysak3PbIMYGQDpd
kkQVn7PSoUSJuBQZpIyyFAFvXVIbnUVoq9tFT4PxzLepiUy7p3PsPxxf6B4G4bE8kJucVeM9z/XI
pc25I+eB3o6N+u/BZR7Vj9OcOi6qtTy8X0EbhhVuxbGENc0l1YvUOyhjBQL6vL1A3lIOBs1Jzr3O
gMTMJ64KX5jLTTyGs/jEY+SGNA+JZt9q2O/oaiWHrwqPOq3nBjixs8GM5ksgWBtCZ5dTlMxUZU2m
9JWnnpGoq85Y4/UrjKhFKILNHSs9pPwecJZKCrYTWoDY9eN+1KobZPBc1nl/obsJaayd2rK3VDkW
WgkfwXuoBdQb9KSLguqUyF9tKIIyDKJl4GYwgZLDbTlyb//obLEHUnwO/gZImfUsd8JssUhAjPXx
xTTA8xXhx6BUR2fel68RG95tvOiiGB0G2WsUu9LeR34pnhY3iY/+DqenM5OlKQVZyIZNKwcl1axy
XcykSaa0g55f53263+I2iaf3g4fz0S8YYJtDwXmQMdgpGMJBs6m03IpyOwlvaF//03U+dB5pamX9
JxjD0/3MpaN8/dGvpitmoDKDGzje+QP83Ytj5SZV2YVZxJVmYCJBmBEfExytPk2RGgxTT7uZXIuh
iWUE9wh7e+11uP0aPLQqwY1BJFm2xaBdn3hY45VpoaLl65nF+/aikEdpcFJlAvlVNywcuPGg+YYj
huZ13eJ9Kt76iOBDu3ncN9EK4njmGo58UvOr4l0HV1lwzfDSnzRK1YA0Jl63KIv7kj2NR5XYdPc/
idRNKbvQRd+VcMU+OLT9NGkjJ/ZcC/RuKpP/X8jXtSb/OC/CJUHqY/SXjvvvwBnlmZU636hj8NXF
LRG1YAYTjOdU/TH0v+QFCron7WdU3KSXSKSDL3LsZ0uGXCLHkbkyAlsdHixO6tKhPrNl8BFQvegT
EFMOM5slSyIZuyjvAfI8UlqGyrvJIm6Src+5ATKAwT+Pc4Km8omZIl5HGzrbmYh9765pofQuQ7Mp
Wp7ssAtgznxBmEPCg2TffSF8CV5RiGf5IiYh1UIVDwLe+yZRRc+wpcoDInoTXg7bFRWRhbcghZWw
Vdnf56gRRCFygMLGbV+qwljvB0Ss3TTVt3E75MCVMzQChcyQiiCb9a+NXXgCqZn2+LvZ+yD0bSNg
DEFAswATPGSvIwmUE0PjVKpwyKsxZL9ibYF1MPYvOx31Ep+2K5BDkbLBDkRhpvMxhG6eZObmnKY9
ZugVHRwP/a3QqOt7+k2Xo+vIyqUtSj8u9FItV6uKeNVdoT8Z1s9t0WCRK9FbaVcAkFu9Y+zLJZzJ
R2C6KLCTDvJayk+s+QKssbs0PUAhT/MDLa2SaFIyjhkE73428cWZlYJuLtMu7PTY93eLsZKR6uRs
ungCeY7/RBGrjn5WDRkaV90QuyGdQDyIZMfPOst8MPWmm6O+RAKVO1fjhA/sNV7e063R+HYFzepw
4Ix67rukf5uCIVKEBYbD8gaq3PbW5Qmco6whcI+YC3jKODdo3WXC+iKwz+glcd+ETZ+NMs93tKPi
phjeOcAHgNV5ctu2B4dkTk1NIOZrO5IFPk//wd+L8gN+d6cpsEdRw0rC8jshZFfEBciIQMZ8wiEC
7G9ge4oZpUbGnNXg/oTihDcXNSI27od8qaTrF7ZMhF5Ym3vy5ofK5ORBE7Kw4VuB1kvQRfIxOlUZ
U1ZvLHrE3/kgPQEKaEZEHPPKtnuSVcI1fYdYnJj1FhnP/y4BL7i6gK1rNPm2P6maQgJiW3382jqf
RSu77wjREBy6/KmxYQPseIX1jO8qcLAm1WqxKMeiqBjo6L1buUszTzCEMoWosAYiUDI4PSLfmsL8
tG2bCJi+wYtQc/FuPZfY+0YA6vxz4R/MYs/8p4hyANb+a3YoStOLZyAgAPFG2EuGWSB+zhmPe2xg
47j1PCoHGwzFYbUYjOg6vaUf+GF+DB2c/ytfpKQ3Hfpex5B0ojqjxpJxb2ai9L0skwYvJtHRGGuZ
pRAvlsZAWpCvQbEwl0RKvigjKs+Gdhte7UrtPertfWG8gMtHb6/wF7glAJIvEyb/6TSiIwQd/73g
B00s9gwc8A7Pi/ecIP5xXjUcmwZpfTW/4832w3lbZA9odU1lb0sKRUJxvSPmebr/zO9uCJ1gn2W9
C85dQy0Pn+59V9dsZCDJ4f2zyflVBrWlPdwCwOI7/hu0vybmBF1u8/b2Bg5p0zArcKDDDpypNr9F
Pm0HzqWFmKKIntuZaTZ9Ihs32a8jZyBhqhZzcYLq5Dx066vhs8tT2wBUjHSIBGjN85qo60N4/SHT
hgIux3gpqtk+2XpAvpBy30Wo+1HTtvSlTU89TEPRe88ren3m25oVbo/ScdLViy56pQQDd1VknhKu
wX2Vjn4esKucQunCJXpkDNv90GncK5jj7efVRaDIQP0FSKaMAELH/WC6K0SmlY9nD6ZF+H9blnGf
meeOrJVhhPjGsnFt79sJGzKLun5AXhrIb6wJ9NnddnVuOvPr4rRJWGKs5jAEo9sNsr0Qaqymze0c
JnUCE2TBeTmI/6ezFbWMFlVnm39G0mAclWuZA/IMLWU8Z3qc1wXlbYKW42R7AlyiyHhs23DAreRS
d0HEfMw6laNzWWpKjFHvQu4OosmnSOJHqga0ZUJlE3DgaS9PnlX3WSwCqtkasvft0IhJyuHZoHI+
A0adsVeaFlGNIi42bkfSugxQO1aalRdkNRyDEDhHMEqxrB1C/G/yfAHxsNjCdTsn+j1RHw/Ln3Cw
qGIEdlmSlci4C0XnLF/LMxvwf1DJv1A6GDLdliMgc2b1Gqbi82w/XIDtASnYm5D1pWgyZp5bDmlA
PFNuyBF83ASyB0qxZRMCzhOb6CADKVy3ODy0AHc5nJFJYxEFHfZtdz5xBHmx+sosZAxdPq++fPLn
XL02lKf1cD9P3GP4Bpy0aZckOMRtor/gjaJYfA+I8tmDMgnrrtoehZiqcDHH2yoq4Ognju6TepRg
L+60DhoCyUmbgnnG+x+68QnJonVG54GXc0ALJ0lTMGz88b0Up66w05Igsk/YuIijy5I6comSEX2Q
HeLsSyZ3++URrPKW1okAPszcnt6zUe4M8ctzbwNRSr2Nf2SEs69ID3eFG8A0PbuF844OPbDFxGN9
+uVi1gylpqY9ISxrcoRKNTNTCJzoXNamhGSuSGKbFwmIwZ0/I0UGMZwDuNjw6OxjgzJQou8beOaE
nr7tzRmPfqwjS619VAxYeS14+cs+hglEWGZ2ELBYvfGkfcDExfjVg2cYAESHQ1yr1J0XZU1C0kqI
OnJf182Kn66l7E+qjxDmEIrnddiq/cybk1rDZgrU0mteuqBswNAtM3oLabIDrI/s4/f+AgpS53uI
XZapKdAMeolMsiuKXeBUWQqB5O/8iOfCu2m5ZeFAsMqlQYy/xsKRoNF/Bg6xuJf7K72PJt1EzFWz
XEBQwFjiI+J2LbnZ4ymM+J6CmqmJ2Gi78TBg7abh8nOtmGkZTF3HvCnwpdu4L8+f87lvxYjt9vhn
UOg4NoN0x3zE0usjvdmF+xug87SqLfvryxI/q5guOgKy+SLecc4qpVl5nssFDpEY8ZZ269OnMexP
CSzlW2SkTlwE5FAKdpX13O3wBexc2vjRdqdm4dNqs8RVlmTvXOsmEBQ4CNTBhxZ8lo560X24fSHK
55P3ebieIMXM50GG2HS4zrJ9Qt0qnbpgb7KKTGOKNsQGZ3b+XaOIX5nOg4Aw9xs2SYml11+SOTSH
ZhPmkcZ34tEOlOmcFjd2iB6YotpvHiKUL3Q5ct9lsF2cPedPlsaGSrPBZJ4HSwgj6iYVDuSG3bs9
X0c7si1KL2NtD3EYvLPQVGAW3x/9Zvi88Lry6olm4U5zPwcXRCQbWeI/ywew1i6RzDro3PNKZAj+
mEvCz/aBpllC/zKXSuAiV7C9F6ZTSW0HUFqXe7LXFbJzC7S0Q0vlE9bSD/5dqPdRcv0FmK1hm5hF
kdO52AfUAavixHR8dHb8ZZQ0t4TeZ+n/UlZ1BzNpDCNxdx0nyoUvREzI46upgxShDM5oPNR4VaLc
0gw73hMXIe5HYt7+GB3Kv3L4fupB657Kux0NdBLEyHwaJSV5M2CMjKU68wqlfGGy+N/QviUB2IL1
azgIgkzr7bRe65YfiXPd6aqjo6AkKcYgY13SbP8jv1DrsDTJZ+syl16ArLkzoiNIjUBfj2i9KrHI
XtAR/sP+xw5n+A+AP2JZfIVvSmEFQ+zZFC8//5gTJisGltpw7vDHJrf7gted8LtbJ23OX9YUlSAE
gTCox5eGjZ3CxDdfQAT8N58OiPSRm04Fn/nO0HvldIXYM1HNAdvJLES6xqgp5zH8d7ln4WRs83sV
DnICWDJ+gQFcDvIoG4qepT39Qs1Kl8vbqDOaR1Krg4OLpY4BTUSecPEQyT+v/uBzBOb/5J2Z1omH
sl+MHhys86PXmuTj8Ga3rfbhf9agZ9kiZaStASwk6vZznjKMOVzvbweFzBq2aXpHXZ6q3JbSppAf
r/NFKIzMFQ1ajnKpm10+fsefQX2xshD5lfRFZlriq4lZdsakyahl1zkqi0XdmBjSFhEppUAu8jnN
4/z5ZsJ1amUc/1My8LcWdgHESVU37xqVSulVbKvyiPCrKwmRNgl9J3o4VMBsOSWYmfUGWetUjIOd
HrwkYoOABtky0MKw7B5C9xDyRzUi4g2JzoDkrIyQRORseAudJpqLLbuKQpMDukOLIh4Da1ogSJl8
n/JlSVwmPrIuaavEwtbFFttvOx8WYAWCib6ZLtC203Z1Y96sGSaEVYVcKVmcZRL1eRU3EWYFhOHw
kmcDuQf2tZBXu014+RJ7muqTtDzVt8Z/K2vwxbpRWLSP7WrCMgh648us21kODgQXZP9KMnsqyMa9
moUG8PnjaT42iVyMEhGs+f2XQ0B1AvBnxwx0gffU35oQbUrTGjWOBGIxVHSMljgeHFMqfvRnw/HP
5ymwISYQNDcIChopQ5FZx8jhHWD0MqYmXfY9Gp+jAXz6WXNSnJOccgDExFemItI2QJnRUVj/0n1M
hX2JoJ7gR6KCpGmi31ccB0u6jIH8u++vpP7L1JnKJHLHE4PAACZQf2YnsRXOoeF1Q7sH+7qKh5xu
Mng438uEe8RgUElsBFxWIpThm7Nyj4oUA/i/xCcn4hqo5AYVY5ouS+lCwC+symOeEkjWtD9o8mCN
2GiZb7ax3NGxRbIkTpkEmFCRkRCQowOgx9Zog+MfkQSlsuUXflx1urECCCSR8rQ99EI54Ze91MGM
4WGnL5OoR9Zv3bxiy9ie+hM50dfdKjOKRhT66pMNqeUjK2lp5Ao/N6/XGwsN2rpFY5wwno3L325V
J95aseMTO6NFXtxft4obiNg4Td7wIu9sO5CNSYs6qnztXWzT1AJPYwZtz+1BrXmn20oS9+mGmbWl
mqyOr0g0mvw6D1zl2a5Ra/Sr9Sx6OpZfytsQg69M2QXrSXQI1SpZvbA5Z/ZN44UroXsWWPvZrkVa
vjW+UDfVTEcqRKdPc18V1gzKHSxd12LwazppGvJEeFVWHqJxfgoOpiOTTNz0yRSPi4fxjQMQAUMm
+5iqkZWTL2Hki21Ra/zHVRkuW8KoyriZvahba13VAs07Tl74L5CzEfisljV85QzfxwP1RP38ImL1
iafP83PMOQVHHS+aiI1q6Bb0qyGZHkWklKv/8pTBQSjtT7PpDMAyqBDoJUMaZN1MMuwZjZ4UkXo3
RUtrIY0SZzJoxJ/JLgORsnyWFWx0QGcGbqE5w8NaVj9YUocFnXLEgiY2ktgutDyrIqCd+bxx1VFO
L7s7mOor9WD9wd+U2x3dhcqNeaAQRyrNJNhZWBpmQmsRZyUGzjbi0K1TfHMg9BGieB/M/abGprje
/R0kCeuOVehI3bO5J6T0sY5eHBq2gnvWInGJ+bEdH1L4rvc729X7wNEoEq4UDx9kqgkMVV31PABR
FVcdp2wPOycX2OQTT8yRnsuDC3XMAbQVoGaE/nc9Ph/k00Ospkh7Xai14CSpQ8KW2FjyKlBWnbxd
dAPPBT+i+efJdW6lIiDZ3Qz7MbX/Ml7hDRWNRBOVnU8Awi6IhwUt1PDEkf6LYMgQRnYfKC93tWhf
trWqI4IrOKQmg/g/SQ2HUNz9hFflgNlNWKAyQhy5oU9GG9GLI8/0wbezUNbWwKTNpFsm1n9YpsVd
iqm0BosIAJVEzAnFEKzitYA5QBu3byqrjMBTPXpXJMQnuqSolZoe2OaM9cDQ1r3iEvISHEQNZ2Wo
lV9QwbC0eQn1frVjSlbpK72va08eNd12zZ1imNy9Gnh9azNDE3n5+Flwwakr09nviLMwdyw+djMX
8y+1haEcKA/oET3lQ997ChxDliCk4uPpRi2SSXWDRPSVSaDKM1SIuo+uKuigtforlNNKGJYG6JAa
T6BDBhzI5QPwPo9z7o4v2pK+qNkPC0VMaOtEfaNbNHEVReX7q56ix8HUh5nG6NG+4OSCrGdZgCzL
tw1YG/ESgO9kkLx6I0jil2gLFPeu4ohe+4odflzwumhqYCVcg3bo0GejdrXTJrdwrOYxq4PzwX1W
TeU75J9ZwHvki0+FwTS7Yi7SKIG289m68SWfXkLRkp1kddlR+59QLgIyxs3km8oIYO61H1TaII7c
wE2nBPJIHBOqRu0kjxCOKEYoxoPDzCoJl390ooAOIEc18uKEwC5dXqm87TKX+kbhBEmQ1zgev6P9
tAhUBvtHDYT4r7+V68I3GiFTYC5K/+xaf15H2Yf79D/vYNBdBUnx/qD6O21BiiyJL44F22OkRt3l
FwLAs2Npp8BEZDJNpVhc3TzHFGAaMnU1tbNpe6ng9ddCKGTAD2iYnKB3y87mGEWdclbIPAKdt/fE
G9PTrXkJYTQ+7I2KvhPSUC7e2g2+ZYuL9q338oRCgfJgOjdqWBHf/cGBjYL4A3nxU06iwmA2f+ze
8lVoqNohzot8VP1U+but4z4uoBNGSbk0EemxHGCtX/xbS5h1bdy6BnJjw2HYdkKN5JnYG4LAtch7
NHC32FSv+gwpcpSW+NYvkBEzaBVA4WLKiJmwCQuX9v5tDQj194GQd/w4rO2VD86Wjsm9Jv5eyFcI
Ilmz9UgDljKkCIk3f5A262IVaEem8XEVSrgQF/DzVUdQT4Y57kQkZvORFp5OrwMtixJ93hjNDX6R
KzsRY4ChfFQmU5Gnz7WDMcb/wkAmk1foaEEa1BB2Ys4hZmPbL1oXC2jkzykHXhEhm2ChpaKOictA
Obbwzze/99U2STaCPthq2PyxQFB/k9NxCuQoYEwREfILB5ue78sGyy+piVE2ZvXfat3VNCa8kneI
4f+Fi8HTF6q7M/mb334ZcfAUeIigk/0UmLBiPQlZGKyYgpxKZ1T7JyqxaAAnUI52cTPhLOL6DIK5
YiE9ahZTsH7NnVDXMLMIuJNbqz14SXSgqA8mpiY/j+0VIeBeKSzxaW6GTQkYY9PmQi2LFcBAbIlz
9dtOXsuF9RQrbQIAP+tZNkuxOQTTGYccHGkU9eha61OEUqmbqvjwPNkBi83ceCdoIAILhI8ybO2a
AXIWpGYWEL0KWaUtX6vtEQxv55tu2uUK5giaExgMTfWemRBeFSCn0KrMNF/SqoUgmHhKLL/fitsQ
cbg2fuaID2P2fdyioXX8VN7idThEWC3Ayz49uxkQUo7oF3Ms7DqbdbSIrGWM7yWfMRnjw6tYa+jF
QD/3762MDMG0FDZgpKWqaR174sJaP5TG1mnGCH6pKgkq2z4vwj2SGz/KHubN8bCRSyyb6p/DgtN8
5IevoFx/BdDxsnN1jVx/NxlZGuvWdC+Pk5NILRogZ9Z+yXNLnNE6mZzDokXqSdQ6lOD8fQT2WNx3
vWP57AnHiAsGAObe+y4sCxnqo66hAIGjlQmCRrgBTpcHZGgPBsljSpeBLfz+cm4BXeJYzrF6ZoOq
xvu178uIw9xkrPLwNU7t7h9WFqwu24lqEjaUdn+vynIkvc67Ctgvq5WGT/lSVMWyk8iPDuRPWRKT
WWrWfuVY3/TohMH5NAENVpbBzaWhaoCFPbOVJSfhmZIdE3JAbJMZjRc/8iZZSYPrND545ACY3ml4
O87gS7AqmzaI6Z5/s8ht7tH08e5t8NImK78TUz/lbHU2Akn1y0p/7Udz5PpJDiY1pA91VigegVbd
6wGSb3i11s5BEdFhSQHMpfevD+XQ73J8qxsUjlhJ2DicrcYPvPxgzVb59valVqhjuW++StiSzU8x
cpYM7CMMur3qTmKCNAB4zbfViB0Pxgm5fMQZZnvUK10k7tjRPyj7iR6Te81ttCXk2P5bWaqA+jGW
dC3OANXai6j0d8vkWMc7WOfQHBmvl8K2YCLGGOfe6IkQZDmPBMx3Kjp2iVLCc1hEGSFY5CLMqmQT
SweqFSPSlkfLCBRzAfJOKvL0Dc0+8JD5DszULFzrjCd4BYJ9C6SZdmy7a8viDkjdLQrRvd8IG2pr
U7Xpcf8LYI/uXHHXQ+4GO2sUoZt6KXssXNAqSP/NQSuJQ11PV5AwBHyvuxdlarsVbWXYV5Geb/uF
DiqUJRLCGav/z8zOcAl3pefwQm3aTZQ/F+zOtXVRg43Hcec2SgjXT+VyrC1nfE6uGR/lenVN4I1s
ash9ieYdaaQQvADVbO8nFS20F4FUQOC7DQTRtTjganglaJ1YqnQo0PqCbIvQpFDB0JVZi9vAaJf6
t0zUZWG5Fvdj/5MsB4jo+/fSOAdiFk/IOM7pPmQvF2vPqQ67lyoyCTttybX0ZSSwyLsnKOEa/Gtd
7d0++knIf8a0cXsx6pjzP4lNG4j4MxN9HyX93XDySBCc4s/Q+uhtCyj4Yqd++oTJ4qhKi6Mn/zoU
vXUpVfE5KcSzNEUi85UJ6CChbl0y1eHi5l71NQ955Uy0N+ALw0095PMWrl0/8TJjqqGfOWNbZQf/
eXa1bEFVr5mWpudsCcd1KMqBbPeA92EtT2ZJhz/TBqIGTg6q6LMz0TANV9cseIHSBGYzv2NIToaM
RFK29XFh9gdk4DYjMN5oiALPuzQ6oYC6ImJPcMj8Ca0C+0MOvBUoSZtsGVvgry7ukiG9D6Q8bT6y
7AOEyIWKyzZJNo9c5hWexavBoveLIC7OCj3VYi5x3MLIgv93+kHOY0lrPA3w/Jx1RC9/ff+4+gxu
aiMdG1/q203x1ZhPvpVpN3guTSzqZ5b5uNfq8xRAQvTN3YO5lXrwHbwEFcdhxBlmX8GxCF8Dx6sf
7aZfSyvHm4GNtL5dLNMDYgPtQbajGb2qtD+UBCoxJw8yG8I/pO2ijgrMG1x7fij9Y9wtKgZBb7Mw
S/X3LTky4jvPqVj5YkFXMYzEw/3CHy7Rtd6Ux/M75Cms0roHKEHp5UEdTxN8wbocHIB/qeIdwm/C
m/0B/q2yI8kGIicHGP/DpQ6eXADOZKeXTSB9wTh/aTzpqiwlathvY5Y6nKh4LHvxxZpi5FNJWzAJ
m2/aPO1twfbYgW5h1jbHJmkZT5kzZDHgZRqmxpaHbe/Bxi6TN48RKsq8kStxbrA4qo1d54rvgMTZ
aVKK04gIB/LWXI1NKRqrRBUKKQtk7Bw1znuqAZPAoPDqv94LjRl6PhtUC+MpqsWXPrLOY6Uk92+S
nKLGeuLSXq9t1iafc+GaI77F1t/1DyhKS/F6DGsaG7BixwFMrV8GyJdWq7Hz69b2Jgjr7zmogO3s
mCVrSRPkiBxN1NcuY4D9SCuS7x1gGnst01s+drPB3o0Lv232i2B0A8OQoAypc5TuL2QUza8tYm/H
SkNuMK/cfE+ea/Tp3hcOgpoxE1nVl8/8AGHqYTAfRU1dcai2kpNAdcRSTdPXLhMyI1+x5n6s7QmX
/6ia50ZqktHFdNli0L+jFvv3lQk6Jtyescx39wvgStP4901nG/TVt0xL9MtBi6PDNX874kQ/LZKQ
5AXLwj0SumjsodFzXdImR8arQN2AFyNmXdEfGi0xgaMxTR0F/gYz1wKrn60NMOq6cqc7r1eQs2ii
XNB9wQsvysIROomXuv1VFlC8YHpqIlZj83mUBDrBX0EW//05ZScEjXh1jIIoBPtWjcSKI0Hg4kiR
DDoOYIy6oOftAkfZcsIzVuDXTfji5aEVZV6MsNM8UYTIC7w9geYavm5vM33KwDj7ZiQazoC2+gfc
8SjNM1TWL2yZAkWj2MFTYeOF++jRnRG0/7MuCNUvjv7m3oxW3GNzFT5qtosn6Pe0MowDYiNAOOJ+
mAplwnrm1Fgonovtb5GWihMWUOB4ofJJ7gnC27hGN9p5+lORXN4xw4wVq0gH89DBpqMM7HiXI+Pr
x6wjfzHqPT6RnKyUrrMTdoYR+H3BTf7IG+xHxjb2bu9hvGok8j7vcmyQol4tjWR9yvNiTZVu8OwF
FVf1lpR5+xEldbvUtqfmw9sUDO+crQYPnaNLDzePhUEzSw6RGQJM/xjBuI1ecAplAN3gg6y9cFvV
ULjzvAIKbG9VpfGUISEtQ8a92lhBPU+b1Qbc5PPypILwCF+zsPiNnTg8LVoJi4O/SG1WlCMznX1y
JDmsNMcvRDsE/quCNehwuiOutk8D8GdWh4a6BEfT4MTUWF2DqYF2ROcABk4D1nzS3Qdm6ks+DVSY
2Gh1OXP0dlKl77Mz7gBSyOL5eWt1HC3gJkoiTIiJ9mmIYI5ko2WxuwvjqWNWy5Vr7S59C4KnWsGA
G9PV5aUGtnasdHKoyDOb1XaLg18KsXMmC3SemjHrIaFjAkCtLojxfpB4NGIxeJsZVV+yrvzw/EbZ
1QxtKa2qNcP8TTi/+0QFiTQylZAz6CGoE4YlkvR1xdpDGZ1GWXv63dbA3h4QlU2hOVXf48aPIXBZ
fBKUDKpiUpHH/+RHSLNbe97rpYHVe7ijHSpHZJUMth2KDn8ftFkhI3KhF1VPC0s3FMWPPeAOSI1Q
8FkX+LO2V4P5t5Yj9fMk4Ud7iF8BTUa8syaJWKVT9u1J9x9j7dMnBSwCHeEA/tQzbBhQFZ1RZNDO
hvPB4l81u/wxNF+ADkFxy9FQxx/uh+0lggYMY8i1LAF/9OLuewPMUN9mQP4TN6uiAhSJDCPXYgCc
1g52nMlirUt7ws529BGxgUCqhOQ53U7cnG0G2Iy+3gl4KoYIoqVIS95niVc11HuowDnm64gGUh1m
dBDbtGUxHJcoMYINe/GTvbiZtvYimN/+4zTDzUqkza+1qkpPsO8bfLCV/fD5j9RAjblO/JjDfDA5
EGTUwmY8/ycbKjtRpMbxrhkJtwuMKX3OyufSSHIQx0E2o7nlHOAFztJX9KReW6UujG1O63pHaY6p
0vLfVcUMYXxIEqHbqRm7Lk5J6zfB36+/pgkRKv2cOPlWCaFsSoAlDe5s81jTsv6ejddX1upvVG1U
LZ2vmn2WELK7cIPFz17lJmBcZ6heIr3q2h/TR45ECLJSapgoXEzOz8jxM7YG+zEHy8Tljp7++QFU
cWXYXYnrQzI54qJshpeyDU1Aq1RcuBHgJIgL2LfuUpS4Ux7Ru6NaUiA2Wa6YBls19mwFFw0JWlH8
NeeR8Cxkid/aY0jNBfwpmQuybPsIf3/2c6QIJSlNkZ1GWQTGiuLs9Pkn/yuvSZAd8iCXqbWIgNln
A+mqJZBze7xyIH2jCscyHfJSQ1CB0L1vylVpuv9XlVp0ZEKTV7R3r7zCEE/wxoky2vZDCPBAA0dC
thHttvm9eQ1CcN0Q11fV1RPpHDtbOLAJumclyLsnednIpLLNwlIZ31lPQF5j5vAxCZTingChJtul
0wZHGERKXV0sNbCB7+Y/UyvtnQAITIKafuRuBGTw9i4bzyKoTzt7g13sHNvbn+FhDYhRZ95uuZ5m
lfo4vzAobFf/sh0NYim6OSP5cxlhHeGx+hhSGEqGWwxe1SLmr+3KPdUihuiLcMJ+tRSWMtzoTqim
FyRplezdc25y6VxYY5WkQgy0CxEN6VUHSLkgsD8hujQhGWVZUKwED7rp+8130YD93OZUWfFZQnqu
2+SZp/PSmAxVdGSak7rd9h/8v+xiBE3EUkVjZeAnIzj7tOa9qGeHx5Ckq59+pBBLItCBho3SFSMK
6Y3fqVMVLQwoZYSZ0gu3wO0ddmXN806KVmBRbwBe5o5QNReLm6rY78+ox3/G9UlbGE6j/ZUrkq8b
0gJt3qIKH4ODWU+/h7XXL2fyU8HFFp+dfy0z+gUgH8d4QFV1f5/48MdWMAATZsxMO+eF489j5Fbg
eZa4T6ztaDDNwb89CigMCChaG8WW/Df/Aaa+EM3UMbDHnEEc8nqGfeVku2j3wu+DdAUgXCGHISTi
QDjQWHLFsT/NGgbwoKWHOd61Mdr3zKxlBmjbimgIR0vylKIiif8YKsAuX/tcyfQWbiC/dCKufA6D
3DREYesOc1Jbi/y0Ol05AcWn3FzdyoWCFSlbLXVpod2BXCVETxEMxqHdBiXAmPJ/R6w+Zucg/ml3
z/5af1nuq2gIhx4GisTqrRCcOlssPCKMYJOj36CV9hVCcdB26WlsyGIGmpkMQ/VjNHZLDAmzcJQ7
w+T0ndFRA+XKiE8YDeUhcKplxpuuCSi6ttJQL4VLq1ZRQlicSFM5o260hmyxTrivcPYsj3avzxKQ
I7hz4GGl/B1alNS1Afle/MGjCCco0RlUKtyFpkEkF4xtRCCFtXjL7U2K/hUwNLufL8eJLdr94j3U
o5k5+NNdms200G9HxXgt04hxXyUTw1d2gM0tkdRrZ567o4rgDtuAb/w04VbmSGk82B85cP/PcO4/
DMJ7syu5/Ef3oyzHfgUBvHD/40zps6D7S3YnfnZdnAv6NymZ2PL6GWRehCuvMwR/n2E2aFzCnY47
2bXB0uH649TDoF6g3iB++dPU4+B+Emhhhw3H+Zc1+A833dlAbSAPccN+/mmEas/Uo8ZZFj22cLW3
qUmO/+TokqLbWwcKYs+kLLczJd6Q1Ri9TbiSOzG2jOqBTt16XmFekL3X4TyRf9qjZGX8bbh7MP8i
xIS/AHYzBAg8TdqZPip9E+Z6ou3+MNfhIYv1mhIu+sQt2lTC7n91NO5WzH5RdZ5yGEOpRGvzVoXL
B/dbTLZRELRh7NHDophCMkHs5Gq+/tZNEWExKhLFm+61jb+N561eSbCAG4BUMPdLSxbX9xnAys0O
t6lQYKhiw5vtTXfLO5aJhVvg0/t24d8z5W8GdbJSEB+9ZOSOAQ3RsZ14JCmsryW2Muwhp4MLUntj
A2KDZTjqiz9ORUiKTXVNRAU0jvmy2Yfau0pQ0O71tiKf+9elLgObV+iSUxz8iwH8fcKxP9rH/CSY
McK7R7kKSt3YygUuCj55SMQCSJe0Iyb/70VvdeENHl746qjr/dsp5n7ixwyVxuHS25ecdyT09Q4/
k+Xo2rAV6z9vsjXz3BHovuNHoCazILmXjacbetoIcOpI8bfQ+ptSkSw0R4aYC9N89bQLHQFOVYTW
Be5mdX2Kig21ySxvnbOoSav5NiSo2WPhGAa2LOLjlmWUwOk9XO02D4F1yQxJsZPFrVg9jufiM+Ag
M9fhwYxIqBI363weQxUusQ7Gg6nrhhcmSdktOrAerOIS3VeK7pRipf8ywFRtdrGpNPdC6cbw4kP4
Tb6Xgt55jzo7yT8BnMbwSDkkst78bnWIUD7JDptwEfTMEGmBUs2hb3ApT26hhLHW+SGXboIyWbXc
QCazLXdrQLkeMeV9wtfcETAIPW2DuvRxFNCks/3WKSoi1KDioSFAzs1RTUccMZXNQsm9jpApFYJD
nHYEugnXtBsvpYaNBLAFO5VBVvj6OiR5OLpvEPQ8T6daqdeKv2ZQKk20hhmO3zwPnLQQKuXz6+Vp
VUThKAZBTmAxIFz4s7PDsZe9B0DfcHQ7Lbv2qHzPXmw14v/Kd9Qw5ZMTsmbpIBlZfMiEPgkc3j8f
JPRQex0K3iHMxNDhIxZI3LVmSI5/042A29YeNeD+rsIYvWTFzFOQV8+96+LlKUVPGWlouz3iK8hj
y6ZO9HmtDZ88MImV2MvaqAlskQx1BCFJwyzBX55j+oZUIfGX2Y7RnqzqXTW94hRZMIxKLd1PUivU
ZvHTRki9EpZALSsJ0unn19LEx+P+A2PaMCm4CryAf04F3ByLasWhO9H4jD8TTu9XGlQAxmkxigz3
Mecp5BEERuj4gLBQP+H+5vkHoZdswQ3AE6NDe6bv+hMAyvURSO8JCZbydeqM780L5Aqsw6z3T3aH
qoxb9fK+TfuapgTbGeJV1xDEx5i0Ogy9xJZxcpp5DpIw133FFUos85DxR2bq6nGQc3mzLDBMM/kn
OXC5wjmjknzJPnrNBOQNHjfYDR9KOGVIFHZPRlRrHDpB/8OGF5orMAVRhpc8k76E201qBxd9kuCX
o7FsuSsTDFKrjCHUTQAY+BGFPwcLqcAd5v1TGJpey8tM5B2lArPn/Fx7mmzWcG8uNf9pc+gnaBzT
KNscT8/nukOiJfP1yrQSzyvw7icqok7aA9tArKBZi6UfLDEYI95q0MCApverg4VX8M09CdpOIwlz
l20JiLyQ8aOdFHm82rD6Zyps93evsbgrkt4VtbfE9v8Otf5g4obPlgeshgPiD4Tzn9n/WT97jcEu
Du16H4TX8DzELZxCWMycU6yuH7GCjZnpQLRyvZ4KEVt0cKTLVJvS/bX4vgf26axDhJXdKVr4+5OZ
z3cccbhG1I+8JNKkNmWrdEaRgmtwNYWPJiM1nEdZez79v7iFEyOnZYh1k+pDr2PY/F4ti/z6MCcy
JQMgoFRyzc+31p0XCAHPxFFH/WldWk3eGMBA5PFAXBepD1KxzKtKlT6uyA5niMedbnCbpg1oDR7t
A7TWbqqE+UabSZfKlbR0sWHeQ8m3zfBotE2KvgKCljK1lefLI6/Tao7o1hyqsHZ40wnDzTUOdC1+
ET82RKcxuhj8560YPeKCcZ5YN57LYy2/cRgmCD0qFxOVUl7rzZrFeS+A6awL9Oke2mpRUtPyLLEF
BDeFzRV7c92yO4VxMJ7eKsOchUL5M4tskF7qkT6vruOiKOzssVZI7RNyKrZJOpWNfrvYz9L5MztP
miY3wzsZPXUtX+ZjkGA3a2tAnRdcrOOtJMB+xCswWC6JRRSa28E32wSuiH4b2/vU2CqITIEEXCh1
A401k/3b67AWdeCcBoU6pWhHsNtzNq1yL8vFWwxUeWM6lu/W6B2tbeGDp4F7bR0Ii4Y/ZZEROXOX
CWf0KVLjq9/p08WCkakRJHDjtHSBfnRLuTlwleWpW59hoDGGg/33RXqY7+1jqwdu5Htm91D7LoHn
EwiFwGXuzgcSMg4fr+CZCj1SwPHVg5oqgdPi3E+4WrKIDRzkM3GX0qVLxjTFFenEyF7sJQdZ/L03
wfrJFNi5PbXL4eqnx4B3V3uUIRLGm3OThpO0dZ+P1aSeLPF+r7NLAQdRLU7sh4TxutzqZiAlwtyE
zT995IHVSG6NWQUyE3qmGeZK77GiHswJKsyc663Fc3uxvzym4wH076rkhR4ehcAEjC7mB+4N3g2e
QRDOAq8b9FiI/mpXoioETrMfjj4KRLd+1XBqnj3P22aVjSjyipOFyECipJvufhafPZFMMY7f6jpJ
mDhzz0aNpbIe3+xywYXj/w3zq33wk5mqXga77iYgprGZuHRmvEGJrJ2r94RqQP3bFNhBQoT7swIQ
AedLfMeFhbB9zETbFO2MnMfHrmzmVLiCHeB0P8/0oo43QNSGcbpAxaDDOQ6qhvJgNitZs07oDSH9
LFw0N7Ac1o/fy5Fs8vpSM62dapzu4QMz/l2zTT4nJjNQEn4ynzfVghUss6f0mCIe8CU/QAO0AoD9
+Zha93UCr9ZWy01BlCNFU9WM4Vp4aMH9iISgHNv6i4KZ3SXS9dZWWFpoW0y745yrgTgUXYnfubDS
8mgjJ7KpvNtALwZ7PTLQrzLZPWIWgQU4Kj6vdVZrYvNXObWJQX1LFaTBdUqqJS9Jk432zVvC8yUH
a3phzJDsh0hdJAZ4L+s3YWUWist0thLBoTKHweAE4Ca3PxDROJxCA6BciGbXRZlpmq6emHSch+dQ
aXHbWLzEexNXEfxW3gHYoXQJBBYjLZWDt3zjqNhw3b9aWqx9x+JsCbutwhVHNQBNKBPZJ6f5SV7E
+CPRHyJNMQpMZha7dA0LOMoLHIWHi7wpZTYvB6RuvNpHbayjuqZn+g2Qz0zsPNzUWz+NSeG9j2Wr
ajebXq4dXZsfXrWsLuF/KyYYRIVJvLDiTScP4WBwybU3JXF66lx1z39LbX8ZTEPKsHpg2mdMdsHt
uoes0Ixj8Y4VdWsTEGoXfNz2LgsoLZMniMiZJGT//U4mKQLO5S0IoiYi+lT1b2c0uL1itFH53AJC
K9kJts4ZZslnBjLRcMj7aOGqTnuRvUITKYNe3rKSUFxXF9bxDVa/wdrECTEaxRKh8MLa65Qy7rEo
3Ty+NIO2lv9pKTFbka2tCCxd+QlLzUNfPomfGITbhrv77ISiykZ+P3MTbtOvDP9F/IWJvMNp3YeR
G7KEKgvfboGWBrGn/8ILBU8akKccC+8qURRc10A8VumpM/GeEl0QKAsDMbUfI53JM2Bv8mnh6KXo
P7nqTK9L+t2g/KxSA2ml3caQ4xdvBOEZOuJ0en0EI87DonuL2jipmlrQi6dpkAz7zeBUq+T9yohw
ik1EvikHHj47clcq3RfTVhOSjPnCZTUy/PEtlw+tJ+LP5TAdikTmo8K6BGH/9Ryp0RiegxpWXAG6
B6PmB5Rv/znBWXclnMNecIRRTAGbwO0k3ZGkfAdkSuIljqlJJcXyVGvhqBnB3AutAU03yUW3OlkZ
u6YuT3RIzf9Q00/9YSPyJE7dVnmsGFQUxVHNqlHuE7Xod3CQwcZ85dk1gj9GBPr0Y6h+9EVP+Elr
DSWlEtPS0pcFGgCssDVWwsEm8+Yrv2LscHV/kw/DCUrXq0N3xSfiJVshLyII1fJlHorW8YzVpRC+
Vt00devXduHuFj7okfbKQy00aRXutpU7yiI0Wc+hgbzhw+mOa347PJ4YsPTjvXPUXx8nUUR2ll+H
PHbI1g1r88diGaXKgN8aJ9p//jDXUfqxs2TfIgUAoA+6DxMTHIIzbO32jJSNILE9W5Q31GtXTUlG
DWtDuygMHtPQ/+ZwfGEwyCCoXH3PRvHo72iPIGa0b2moMaOmuCCa1oYtTcfbt0G27p1ut72yu/+l
JsqYiY3AlukJDtZK2438atSNTV2aZrkOT6fyjOeT4FSzD6coS2IpuyHJpWlkzFmgwRhypUrWtvj5
cK06Smo4N5iok7x8UUQvGPxWh6eWozT3G+jg3nCIv1knDxO05OX9kNeB8Fy9kYCkx5pZ2mZjMgtt
IvohLXR3Hysg2TSyQSSBwZujMKRmPUCSzywRSmUrVLwpU/5lAwyFG5UPMLZFvpbW13KN6zHxvcvO
OR0GhEddgqY2tcqaUX4wwBKgVWdmqBmob/Xlw5N0zaWWMSybUwPKKHiFRayB5R1rBbXjL4LCGnWx
22IlvGM7rOXv5EgZZrIDM2lC5503X31LR6x3F4yxzvEVOJI+VkzYHO4QJqauqY1Zf6Ib/RGZTfLm
2GTrIPhXtWLoKqZy+8VQh8Ma8L6M8qBGhDYMoARE9mEzhO3G9FZjRlvZMVoo6nQTrxGON5Oi9mzt
QS8t//0+X5QV4cfcKM9fWUNf+/jBEbxF4dIjejRxRAPWIGPKhUdp/EVUDiDHyVloWoic5WA7bBFZ
7pbudd01XJlYAMaroZhutJumoCgULfTAWTrxAtF9b6SLq0FVFZkAcqaX1GxMDZvQvErrXZWMAoRq
PuKNpAI0lmZFSYRDbTVbR24vHTiaRLILKlejZP0nCh+3muLuuSgoMuJ81Q2y0ohE+1/PZkkx4q3j
bUWB34U3Xd0uEuebz7eCOrXvtL/AWib/pNWjqX6FjrBwf+yq9G6C/mp2HuXxBAJGYg6bGUHf8S8E
bXyUeZgb1cKkxaUghvWpLRB1cGISGUD7+7t618X13rT6X0PCoxfZVNj4IJvRMDd81cN5ip3XoN3G
bZa4Qw+w/HVXgCNdZ8XjBF4pZjLemfsgi5L0haMtObWWInuqV4dkV6PUnus5IuwAoEpx5JXVAYiK
lNMoCV530Bhu9IAlGNRCeYQW+aZTeu8n68wRXpNnwXISHhehdJ+9GkhG9gulZUeJEUVSJdXtbeRm
QOBpfm4S75nfiTjiLd+B+oEJQALfl0YVeRgUyuCNwexKbLfUTwQin9pZFcGbXYpTbXZF9GW3ZgZD
0EY29S/s+ehCvNmUeStphMDTycg6VahikX7vkjS7rSjCGoW7lzLpgdihDTgZRKH9wcQPCco3eVSH
4NMn6pfcrP5kaPBUlyzhcK7+FZlAf7cYfSoox73jxgEq0jp2iqu7L2vEomwdnOHV14dAex0AuAlf
Kx4CSu7gLun8CKRNKwX53Ee6vVnEV8B3O4nzevSu9+P/olRMLlZGGa8kmf2fWOMqJRsM6Y7JXOUm
R43UjMyTAlIwRgjhWG6vyxk3GNEYlswWsOqysDzJ0zw4F/ryhj1UklTCxTBfqu+a4IWXxoiH21v3
7f2VaMJ3dwc3bA1hXaEo7OXMXFEk4bQPrjnGyw8CwwICgRn5cGv/uC31x9Xo3DYptC1L5le+kSbw
gNet2cPVee/JUWlyQ/eaw67Vn0jzLyDq5njoyWfYO792DdIFdDU/UGLVIi7PJ1l0rFDxid9GZG93
EiqpDNOR42TnfYA8Gy91F7OcFyITpc1EkjyiBv9BdhKPzdLk7L0Z6NJWHXHblO6+raDg2HF3ZZCW
Bmp3hMkSgvcwLP/x+0heo81iuyMOoNr+sTO0UrximLLwjt2DJB4FIejJloU0Jd4RNem6Xc82bLvO
6SRjBo85EihL9YEqeE9D1c/cw+kvphpN0sHF2Q2ky6/SbY2nZmuMYzFlEZRUl49krZk/LpklFy6C
4za4rfr27Zg3jBjeNthIQzkJ6P6x426NiC9uut42p2/75pshVJdP6WHXq1t5a4faZ6WjJwB70uHQ
By1MASaA5nUCltNgWt71+bpg3AX2U7L9Tc0dXezrujTHt/ZueLpHKULPuAQgmOX6dON9mctkN6Qj
CQZfnehKyqMvk8R2SyIKidGTTh+ARbexSl7E/3kiSKhJoNjLlckc49bbLHnklkvvTzOa4fa5sy6l
F678J+FqzS5ik0RkuS3vfCsT+kTx0zg4sL54SosN2YOQLV9Fn7Pf+SOZbRXSrMfihCqaxDIPof6y
eMPzHOkqQaOz6DPvRlu6x50lKpFiv55FBUbeUWK4xU9ilflNoQl+6VYjIUQESRK1FblppzRR1KqO
N/xkdI+gi57PqS2qj1Excwd5ZqbvpJaA+V1kqpW3Fi6SSO5YXo5tIia1k9wOtrMbWQXaNzv+3f1+
99Zr44AKsBwP1BN4XrwTIepuNCfwvkIUBEwasNMBgfw3p3AdjRRpR7G15Fmb79/9zDLdALBGlPpC
lyQfUJdZoCabOxF4v1y/uOgp2P4+sds2afe/nKqFNOPqsj4iZdBatoeDAcTDtqx52a14u1euRnNp
LzHalJ04gi1VaMD7rqa5G0GYKz2UBfmFWH0tNXT9sR+1Ld4ZfYfRAmeeJPW8L40f9YM1Hdz0icMd
Yk3jG/1DS6CHkwuFNtRaCsXnNU5eKcpl86TOExJMeSF1BKRK7AHGCfZffM4LloV+l7ri2arsyCEd
z4EhY/jAg8h/x2HxM4tCT3PrzxV59FTXiFJGKon1gbj9PW/rZE5zTnqgDY8Mwf9093z+nagj5HI9
/lAwGtzSJlfe15sfdPl5WMnu4Lj8BKFbeOW0l7Wq34iymprNL46oWwMm0IrBG977lJX20IO0lCz0
vwvPjsCb4Mat0OAd7H0VIsQ1LRymfLO5ms85VYo7d8ZAQSqr8Hf0xknADYyIetkbLbMGEHtxgq49
s11tCB5Rg+cRrfPdHM+uI/7/xoh9ugzwXiUFr9+gdPGTdBBPYg+UnRxL7qdKXf9AIorcJMCio/NE
Yyi4fkKrVH4HRFeDyvukcgDkvF2rzMGvOdrPxiTLawDitF3MZkyXx6EBGupAfa8xApv5Xm1+oh1Z
yPkcIPVuQX6hyopds9v3yO3rxWQeGHCoZQyZq8Og7CCWAku85u4X34SxUKZQi88ENpY5iRR1iKSF
LbljS4g4205XG2BCYT3+hnW3V4hN+2wE/hYHun2Ja8GpV7qaCNuRZSDNd5LrUUlY40lxZI6U1raQ
lMVHdWC+CNYya2LyQsKhr/BuugtDI4ajNGYWsQD1sH5UrO1Xtz4KP92p/LKb9ItuYT84JKQqIxuo
kIToOwdpHsiPo6/ulNMcqSxod+erIWNiTHBBkMfrJv5Aef5jq/lB3a55uu/1FjlUQniTKIr8g1X5
UFENon7Vl9PwE/+PAMIkBwJMXH6aLx1V0PfFDoRRqlt+lq9m5FrmBbS1DkgvMXD5wpxAzDt90kxA
DOGQWWCHQMh+K/eHq4rv5IXL8qfdgqJ5ypiHAdlyojlkT3J5HloKqwmH8mxhFSQOqgaxAlk/CXaX
6afqO8wWKd0ORhf3EH3bG9FSEtJ20I0AsXk4QhqjSlb5CUX/Sn2yUhgP849KXnEt5v5SzlbCaJpI
gD/F+RexgZwKKNrmvK/IY34ja8mSpDKB2FT+HMRyRec0NH+kccf14CD2/ppZQnJXfcPaKP1zJrQv
Uo/xeRlSGEbi7T4BLrjqF66GXI0jMdlQbA9beI1x8T6YXH4yo4Nr8IbKT1OnshypDeOddzI1YM8a
dy6xi+H546heWnok/MdBQWyHPrShPsfR2Ablz4hxLYfNMmV/j4MobYlD9ROdzMjAZahnLFjQTicD
lDZ4E9Z4qKPxIE75pqwHqGqc0CjVlza+Oh4YFumx8t6dGYjvC/vMez9mK0y8g9l47bH9sS7r6RfX
05sIas6A8jtpIQcgBhTBznoOdzyJ+S4oAA6O6QAg8rDe+ixp6Dx5NN1olK1frlyJMHL6jsjdRW87
TN6dD7Op6tFjwuVtTPCBw6taiuBdCzK5f6EDiXMpvCJu1o1h7tyjJX2lz9GgP1qcxqvpPr6YdNDM
y6R9QhT/JLqpCSmLGumhrHlKFj18q+WPnJQYlTPOmPTEtqqcccuQF10Ya1FVqGrTbox0/pBKncOS
3pJ8e3u2R0U/75a71d2QhYs3/rvoEJqlLypzlmwX+ktuWOEBgsZ5NLIrDztiGhGUlUVM0B+hSzCk
MwlcoeYcpc7fpJDRS+/m0SlahqwjsPh2MDUUPiBm0uDpoWtiLHwiAALtZLTr4PeMyDk1arIUzVqa
3I3aUREhEImE6FjG3hpRcDqXxl3T5nA3b6LtvKTFgnf+KtTaOck24Skmb8GPagzMgyMnbf5lHW+E
9Pvim3nNvvUtbQPTdDGDbpHM6ruW7WoNh69dJybWcv25BHr1B7OENDdO4WKsecgHhzVf/u1qxsDM
RhmfCMrSk8g9O2yfDs2wv2jPRXfp/9tZV57iR/kT5iFFmoM+Ria5pvcMcs6MELxMt6iC0g3Ox0ky
gPba37lh7ccEmxwjWQM6spnhGZs/lU5skrkkC10AoNgbxiAaL52hsQkhI7U2UVa9GmvlG7tC6+yz
vOBMLAvVnlVyfMDlwdmPC8Az3u+vEttbvzhCnyWzq+YZarmTw2WRnwc+od4RdAUG8veiqE/im+bS
ueehxAY2getefy78gyi8DdWt6xhZOlso5d42P1w8xsodm9r25ZKm/d4iz7SMENbvQOsY8BeEyQN/
mxRBVMcAHQlfRiQccON5RkHALi1GTlX+sncrFhQ+2/djoMuJWF+c/0LXEHP2DVfZPeFp4sSMSdMV
lii3JD8umNe2JSXvWxx7zbq2P9T1z+lVhO+8ExuSWFi4JI5cbfYUZBZFLt9uohXv2QN7UJZFmCTw
XXTH8IdgEnlClj2q8XC1P4w8+Fc9VallwGoWaNYP1mtxQc36pqWCClrx1iAHAvTTuBNxr4VAhkGl
CHOiJ52tplWBXLUjlnf5rj4XBc7uydYRmMiQH0uU01CdIDcL9m6nVZX3qiSubWZM2TkyCauxU2NF
SCebwONiLAYGipZahCG5CR7+OY2poLs9X1F0y9jIDaXwU3sZmx7spgyMphvLMbNLGbGoWTgQOl8r
DYkmA/Iv835TWykTquW0ehF56u+3zXqSDpK3dHL7HsTwv9ce+dENV8gq6smgYFyfFHTbUlEQnvaV
3iNNfgzJxB5x1Ae5vIYM+cpUr1oX5AIM6qO2belib2BEv6c2rlRfv/6ScG8xeTWtduPy6xj8bqLu
uGIZtYO/XorFgP/A0h4C21LxAbGvTpyvBphi/jLD4S9w378XXq8dzSFIyxvjxxAxvMvgGdXbCD1R
WR/b9Aik0/qViwYhcWJhkzmXQDUs8/Bi9d0/HUsRleW5PQfDasEnPx/p/ZJC/0oscdV9pPUEGYvn
3QEb0TAYRSh62me4IZNieSwkcIevvShFj2p2hcZl9TWENJWR325s5kdpsC/XqSMWcPlJkR17qr6P
mp+xzk/l6o3j4j7psMDUIAanZ5Ofh74mwy8Tn1m+7lvrcp9ofQuOXbhf1+UKM+uHTw1tAeXptr2W
OpkogN0d+zONN2rt0gijefFGsZmCYlOQOH96uBLN2S8ALNFAIV1enTgKQwjdzrhvrpbI1cnSHiog
f1dxkCJqR3szMjQ4YOD0Kin7j8fXuAkYO2jdg41qB+swo1Bqs4/BLNYxPlJ0MePGTlo5nAyFEHHH
U3BmpnE3Flxy7e/A7qCDirKTvGy9xuVuaU7yBdO8gqn8rEv9AU6vIm7oLq4Fq31WSDoYLcbuENJ6
8jsSYfF5l+dJgW/rTm2OynIH4satN/8e1WOND4q4Uztrv7xzGsoJCMRdLai81IxLVubydY3ZjaK5
hMj2sEHvJMwx7AQAwP7NM+QYc+GJIcYIEEqtgmNxn+rXB67T/gtZ6igm/6jxtEJ8xNlHoVFIFBM/
GUC2sMyGjLNZlv7paOPsmlUvBRA0RfJvX37f1nCi2+AzVGH228jEGWk6i0rkzmL4/W64O/max8CG
EIIY+vfS1Mvps7SVVTrDmS/DluEiY4xWfQvF93hT0C6xW8E1O9Evv9dtQiumscO/NGrMO8ZERwRs
xVIvxMS63fi6EmWtvlRxGpQwlqMG9FJQ8ax6KDoox1Q/roJlP3xpz4mdGI6rceNCkv5c0mzqm4lN
0acFGi4oR5hWDcQ10sSqmFY9w7t3qRqAwpeVTcIxx1svUzS/zW7cK5THzAwouo/Y2ahNJDOA7WAe
rvKyR1JAFoRBIUmtWPR9BlyKbEaJH+WsY9x4cot7h07Qh3/3C4tjRdKpZrrY2U0rbFCtU2nuy8Cg
ld1UPKZF/aeEHS+w/ZjdPTrTPC6UBhpgPno+MSaxuoj4Crxv3Khn5Zi4G8ryxLIx7f7MjWhA4nMT
J2lMXI3HKx2CGaWGojXeCW+G9nrGVTxR0i+QupKV3GTOUxGQEP3+jvLVKsatubY3tkykSHuDCgZS
Y5EVHJwx5/TFLK6Wn56nK5n+p/48cVs8f66bork1upV5w7kYtzwrnuOPl8c5g7BgVDGTEHcahlgh
NYOrtT/cbBYnhNbL44/xVAFyB3fKhmMpo2D0wsGXM77lS0jqfrQfe+Ui6UjnA1UAsZmosXIUIZKd
STQ+Us7UIH/+vfHSxPIzigY/bS9fMy3+lEA8DBL8o+eLS8V1S41cVNnQBugDC3SNAlKxc+91063/
gAskeRkvc7Zuvk3heerLV+LDJB8gI2x7cHqeczCh3vt7+wx9rUpaz3wWME88tW/uwp39D7VQs4k3
jq6D3DmSN4vIPh7LoYX+ieJ2yJsasBim1D+qrs/gAbLZNcZ+rClrGtZt5tZudrm2i3pzcSfJNuJr
UmLPFxvmJsZjRjnV2NZa3QoHZNLfCgJ+pnJv3bPDhL27dkXLlUmF3JBzcgPa+onFRZOw2y41z2DX
fXlFjpt/GYeEP3Qjff+1KGJh5dkas4olbi6Gl2qS4bkCOrPtfbfQlHA5F00fA8DUEg86yVh73ITN
9cDoelQuGPDN3p5q6BF3R50Hvg4k94+DpsnCOLzQU6EpLtcVefN+LGSdDnbRSXRo0vo/MIYre9WQ
mYEXkHHP9FSuIAGZ/QQfoBn4fJDXzWnR373NiwUevzjE+MZm+O/rXaCMRAYs3bv6w6wGHF1u+iBy
8HWbCfo3nsbeOpcgLDYNYHtk+yiuqRc5/coc/YzwRe9RhoELHrABZ7hiO1qwZgYlvM/Hw5g7jBTW
Dy4Olrq1tjoSm494WtFWaSyWyTsIYZk8jyFrBv85/3awwTP5m3JmeB/M51lYwvpR+NcUyFHERLJ/
6KOr5ft16RGqsFLNrnMNgIlz6WiYhJe8d2TlOTUamwREh/Tv8Oy6HLTYUj63Y7w8MLCsw5biwV7b
WtTJWO5lkjj88lBGGyTzj/XDl3W6PF5ka0veO5lpg5Q4o2gi5U4JrNW3xRKyRZM3DjJh9fQVuLEJ
TY6CJTGVjAQ7tskgCro1/VxLRTBWDkWTOV97ptecrcdZiq2tf4wz/8W7RaYxblpMRwwJAGM6HDsP
bx1T5O4OtEkFHkoNunI+yAG456M/4P5jFyGwUGFQBGjY0jd6dqeEsWb2fGi95Kbk218RJVD9OzTt
LOKx6/smv2TDGjfuFS5K4ez+ktWCJ7vyMmUDyGh/zwg8Wu61UA20kulvNB5QLrs66iinGJlkOJfe
0Vr3luy8Qg/F8ds4VImPPjjfCaibcTG6rPzvX/Q/xxHfn9BX3F8gLV3hotnbrdXa2zqikHH7ohJF
Tnt4hnv+u209nnzuxQorPBtlz6Iy3J2OPKKGb6LkbYG/u8Z+1OwSyn811kPv/Le8upKUixuzOT17
BcVFNhXswNOwOAGdHIV0Wi6Hx4OWJMHCgVKBDHJao3U7RtU9226kBGKfZH4Y9+sI0wHzHheJQJdN
PhUhcM20JpCGte50zwBhf5oRxgFKtbLRs3HatFFr7xaoH7dhxTSfdUanW00MnJwKflXNg1y1DFLp
G5vq0XE7inGWIKVmxjVXYj/njc2h0lEeY4Vpm7j4CKoFqGhOKXEx8MgVuAMuGdN96GzSGJRkFGD1
EAjxhRT1RuzO5Qp3yYTTwxZt+bk79s94JwpuvFWm9C9moCMq/TwOtnBEnEB6pPTgtQY+hry+hexh
hdGrZAdU/2tBluWWWHd1Rk/z2K0BBc3nhKUr2XBvhYNkFbM2+mY48Jz++2ro314Jbary5nSI6eSl
skArDUu8l85zoSzDWkFwxGSNMbneJBsE1OpeM1bZ7bF65I/7g4gkY8bbclNickgdTrxDVyBqkjZu
EBLatT2oVTjP2JxCDLyVrf0zdEuoGoWTrf6Q6TvrJRBnPYOGRCj1WhTTxIZVdlqzI+aGmQ2ULI+u
oNjHJZ9ikjFZu9f2iSi/ga+MaKP4qrti8iksX7uuQ6rYesG66aG0AOq/grLNCfhFyPvqQejQNSp/
A6HOAaiczWI1hGcADzNqOsEIR6hKU3Q0FScmP3lOZ8fVtl74esXeFl2CViTk8Oi/Goid5BgcDF4U
XK0GyjJYIi12HpzLJmB+EMpizxAYSF6pqvh1bQ3jTUCVjWhrQsr6GhRIu/e5VcFq2NSw02aHEMLB
YHti3b3xDVmDU5W+IPMdi7tTSP84miDQg+16UjNCcSniBj1rMM7zDYPqjPrpCx06w4wOh5ugYgbP
kgq0BLhLX/47rpIXRa/Ew25sbf+KjFSpwUxnAzwChPyeNdZ5DwHLHS7GIGtwONN0cdIrFa5UBDeg
tUChG78dp+objQvV8Zqpu1X7zpcgWY19yEAQKDKa/m9UhqOQqU0ddmAf50Fs5zBlqj7ae06GuHwp
khF1yPLFDQ39tRe+i/VNF8yLJZjiqLvyHi0O46bDAZgA6O0J2P+1YRrKKdvvP3gHN1cgBQqBLHCa
+dFUO+dYxzw793Ln2t9/ZiCN8+lDOdehUktordWMiAn8yVOXrI5MgF/VtJNqFX9VUJzWJ0rwZvl1
2sKEBFrTzxt7dtWm+9uLA1RM2vFAnsbuBtxmwkfJukZ+4IO/4y/bdttbQ+SLzFQzwGZrZ7Z7/0mN
K+Oepo6fM05kQD7mDil3oXSpePJWXtrHWqSDizC/u8v2CG2SNi2pmPcW6Z1x8gGdkLZXAcuPj2Dp
Xgk9j4aVSyEp24DQgQBhZG5eTgY1q7oCjKuI+MafyYgGLvpre3cf6TSwhTU/50wacGXz3ZwXE6sW
xRi21DA/1odBCUn4VN2Cv4DPC8HJHQBoRkDwC/QYRf9oHEiFk9QICWgewWnp+fjRNpc2bxkZh/YO
2Bewfn4waR6RpU302H/txjQtT2uMeCaZaY87doVEC2cwUE/cxaHymp0CHgmI/KxGgO6s0GlwjDIR
iTgSEO+njHrVNN6sgNgpKJWaKKJ1uRP3QLASN/Xc272aKUzUrSZqZkwBwixzznmHstQGO+xzGk2/
iI5nOt1nHPEuz7s2hJtZimdwURNG5TGSyzZwfZSVOk1/x4UKDl7nhM5lXv9DHczRAktf5HmWMmJw
65TQfI9I6T/6D/q3bXFwmoUqEiuGwrKFDwSAr04QRMMpIGAX3knZShqUL0hkRtjcWiRKx6k1zzxP
c4PqMkLDxlg1wcy/p8xbiZMvUeE8pIzHYzzCBfFEQ2KF/ixr0Sp/k3CTkqtfuKSCk3adnX85vEz0
j534KaYEFHgc+q2XpSRoaMgcKdW7fCjQ5iJnhg6pSmP7VPnbA90uzk+Ky5oCWPLcxKZT54J3hLfJ
wxv8YWOr5ERflm+VR/3id0R8KOaI4ewKa61/pQw4VNs97gS8MEarSCmD25s1f1gvCyf9kYPQIsb+
KzsR5voxC/FvM4TzZnbGhFmeXqGNDLwCbw4m5PWfQ3D8fs4JWv5WZfooSd8DkeV2u24izL+2LSDG
fgtJIjQ3CTjnW+Tqt4jTwQVVmIW19udoHVXDad317yGyd+HakdM/MheITp8qaIe9gK26s5MJweog
d9K57goiP0Q0o7g1FI93Ib3IiaGeQsngQv7h5LOpfUMn4ZBrxMYIizNwFNGOLr6yfFBI9pgdHk/g
fQS6jmqQnD3/fFjpnCuggCOva0eV/lm9p9EP1DLrYLv6FA7ZSyScsl3Ey7x5JbzIuTmCSrH+/q2e
i8RMfiQW+m1P1k/iNVlCbMsvKJQ24XMUEIB/dNuF21AZxxjI1myGKjv7jHvGHSMtl6rg5Z9gx23U
Adq/72i1jR8ue9o6rdtPbnl1X44Ok/EJ+DVsDDkk4L+ruxS4AShfpMqu0QzuaXG17dNdbeTOnbmp
VfoCtQV1qJDW1A/pcL18FcJpacTi0hP3wimazzni75oF4NjyzcfqwU8CkJFRvuu96UGaAHzhRp74
hH0dxI9Qhufe5Iz+abmH+EObcC26U2zSKV3M+4GLCEvlN8JNEKIT0mgZYkIO+rgEGtqRUjLa2dXk
HTlNBhjmx+fI9Is78laWcG97pqwdZtqj/0FL2Y4RSxfalhW/QGrf7bmYPj5o07mYZVTDY49jUHSV
thEY3sPurDC9ep9KKtBHTvjE36BmABvO8N0OIsNfjcFcAnN5jKHzDO3vGOT1/Pc4FMmbWT7lz3BE
KD/dor1nsR/yEbAuBORW4nf4XjSNPpRtP0zr0eKHb6r+aqUefnr+KspzfhmoBFtnIppjZy1FJEP6
/urk+6Uayuc8PcBBOkSPkGkNZDE13omv/0sTSVkHD8qJv19zyMmc0FCqtWRJj3SBPp1w329NG+PQ
OhWPsJgEnU/n/wfXm9Zi44jMIZp0nbwSrtml+LcYcd+fMGxfzf+bGzBcBYf0ynGn4p2hlZMaYeDk
U0CTS44zoo9SPhglEynbliH4AUWW3W6+CiBIbXkVt2eqMFSOgNRKJUvA8xUNxBdpaqEoatdwWIbB
NiuGJlerqyygHcF1ieX1RFB7xm6St8IAxK6DCHShOH762xTF+aR3DrfT1w6zW79YHUEBTMmMkLo+
pctaGjLblW0G86iZNj4GT5hWw0hDk8WHST1ZjxAG+Xh7cwQ3bvO8wu+VCHNRfTS0DLMJe2/IgrZe
Yqq0XMP7YqI9U3Crr1FsECJ/VFkF0amKeV6qOABYkzQ41cb9nuuef2YK06ZMwGqcZgw0FlXSvkc4
X9vHEPk85vcM//VS2WBigAYIBEKkkzc7bpyiKkYs+kuj9j+gmO9gL0h156CO6vuG8WRFeC2W+hMk
ravjpub+0jp/Kx21hQlcz2Qwc1Ec8SOONW4/NUufZzkRCwxQWLk3gt8IyBjBVfPIh5p34ogi/43X
9Ta+i+cHNlK7bkEdwM3gysjd2XNWAayOfEj/ZzwHaEXGME8SipYOCbma5c7yo7zY1c/6lYUEtC/F
7zyfMHA02MxXKNXFk9K06E71Fsy9wtk4cE1P/IKE3EqcG25s3dF/HdzrHkV2Hjnefx8uDkrXNmYN
oJIYXvKEvXCWT6Si15JrmxjRs7G8XTs7n8Ugm5QrKTPNp7UoXsh1U7MIOG2GG9uwPJTp5heF4mi2
F53uU9GpwYEiXPCnp/37XzKmXI7irnU+7c1wvoCx/b1HXv6AbnEjISeNBFeWDzyMMyqmI9Rcd2i0
6OjvD18yWrXZ5v5TlD9mtOIHZOC8sZcc6UtjZ6MP7Gz6FLq6pdZXESB6cSEuGdzHHA//nwyCCn8O
oENTUS0cQt7GqGBj2x+aeeHLIdomex6kvcKrGaEhbJj1eN2vNcsapzkeZc9z0D/W89JWYmV4JPjh
Yyj5iTATIfArF9jg4IGmLkbjoyUzhL5aDu1uxIsCgoWFeiRqS7pUgU9i0RIc2potO/t+m8t9gf1i
7/wVUGSoVTSP5TJW3NFakghSmr5JAcN5maeggj4Fk5i1nzfp78uErxazAkkNUOsEiRYDIlSQoff0
xc/4tPABnTP4ygupuIOWepSpcu6HCfUPggBXEX52u4y6psxVq6/X6klVzBDnfzW4y5rOpUOXU7wu
JTyUtSFQDf5rZRt/zItGlStA+HkrVXk7SzdhmCiKg8r7wBrIWJEHzVaMAIqpT5uZilv5oLkCvHks
D17iB3sZPaZjLyHvUL3BUcGQcTY7SDqouqqGyxtbi36yeR8RY90W+rEFnlT/Kh4sp/XS4u64HhC7
UWDiIq/3wR++NscWMDjHdK4i2IhjFOL9xZmBw0zuONhPoNQ7reYY49o34xZhgX3btn5kdDTf+P1N
VhRp1gjPwyLQQHN4Q4P7syKTfNU5YM0Nxrqn7p0ij1+bun/rKhKOYg3MfLEZg3ias+9BzrCEcdJC
xQ4OwbpS/Xaccpu/fWqF2ANVO+WA0Jk8bj2w3sG1xgWajjzY+SSkHnLE7tjKz2cf+/qLJSj9oEIE
QPA6t5BH83yXL8UE1RZ46rQxxAIc6Gk6jfh76xl4Wlyh3v47+Dws4j3S0p4P0XE8ac5z6YnR4l2x
ubWD7e2mN+MZWl7PoGzNcEKHF7rDn7Ng6WJ5VkBzcuL3HhL0O6IpSyxEke4ErGrOVcrWkkRDLBwG
8WiU3YOxjJYKQvApN+30JOZ5B+Kjbq6RYpyJsRQQLAsooR3EaD68vwneL3uNDKIR6YPgIUDNkesN
6yVtPFuL3nDJYKgDXSEw4pHgzclF4iT+Iz+uPBt1G1seW6LVEgaZrq6pBW7RPngqBYDjxqCLP1r/
oZ/WGTzwynA5zj+syDGUOScPGXnl5WMGpV8WlnWuh/UfMOBgVzFRAdy3J2ns0Kl1Wk1UG9s6pcqV
AZt6w4GROfZ67Y6lGltrfJ7FEKpq6B3PjzGxNthyyvu4ycCJSiF/yglaggT1Th/Vt0XNVYL/Witv
QMi9X8f5Ir6bwS/5kNGl4pkI/WIjDx3pF0W/Jp8lb37vQr9IbExATGyxXoDCwPwkFqD5Zlqj0DXD
B2rT6en90qm47zDP+oFlRfcdV6+CGsexvNvd/Qotp5jcK6PSxjS1PYmhoNuZJVRR696xCDMMF7H5
MI70j+ixeE/D+2IB5K90iD6VHQ/6V1XkplpewegChv7+znA1tyTn6PKCA+RwQt958dtKgqfmSlov
T7v3gAI9Zti45r0+O5+UvOGA1ntDkidhhSixyEF9rR+lYRv8CBjRNrlRUVpXEH/NJqWrvOOIJ/dg
qmlGfx7OjOGqfYIRsmnEOaJvMza5xjURV8CzBHp8VVcoY9FlkPUIfgjiOAaM9ROUm31LEFTEnID1
beUgFoqA3puSD9+MMVr+JhkeHAeFjK8M5dW5ZDm5e3Ir+W0SmGeH+HqYsE2/sb+cTSkiWw/z8/jz
IeoMNx49pGzmTR6we6JPj0FllHAm5mvOGZSoEBbFpqWD3+985AfDPsYo9uKSfZ1rtjwCzUDbebvv
mJ28S4z99jY8b+DfgNIjI5rC58POUuqCdtQ4YT5USJUu4hm1DMFuK2FLlzgHssQovCeQ587TMSbJ
QGn53saOPHsQaoMHg8YlVD0RtThwhLp4GD4XXYxyQMErc8UOtaNyNk46KfQwplwqe1TZWFFCEe9t
u9qy/Y9WpQ6kaWnTKsbnF9Nfw1KrFYRhNuxBGC9F0QiiGV+ltDabkNptAHUDzRAq131IQnXnZBt1
5K0G4YjDjFGK6cAENYuabXFqIYxIqmQD8ddKq3OZqnsmGgJ/Ompbb4E3wu+hz+pvvnswZC1WxvfX
73skkByKU8xcL/JtZo87SEjg1OTxs62ZhSyMNQETVBm4LZOiQMbspUg5AiT83gW+w6Yl6J0GpNgU
81OyePXYz51BglVIURNhhs5aERGi/IUAtTgpov4EvnmCJBmtIwV/W0r7OFm5fTWCPdG6YvFLeQu1
HDFdhUiHsBMu0PsyXtilEws7STpidcKfY97rz2QGIMXDdj8zPBWdaWQYkLoZDxpangrZ6z0+MHDA
iwTMCmRV99Ds2rXqRk9QNPiCp5uRgXhWxcgDMIw8ylHxCbMiUSx6cz3R1NdEj9QD7WqGZlMRlGB7
QBnok2BnjHU/NIbl2gEfceB8TrdACHSFtO/u5beM7GbIxjwXCpykCUVN5vmqmAVqni4tPVtZL9fG
rblaBb3O/G32lJ8iBrktkR3pDFt3VBsE++NRG2jIGEhnfHPnzMjNDMNwoEcoZVVuIAf/6QRccMnS
EGc7ndqGtCmEYvKeTVozVenqJSN9ufdqMk/frZqqG1ilKu0eIkRYEd1D/xBK7nzKlmNGQEAPLYqm
2F5ULU2Cb7WqYoiRCOv6U0lVwWRHY22vR+pKextifwGv0ui95LRwPxrVZXbP9y6zAbxvwLEhTN2F
278XfmEIQ2EQxts1dTvI6/UbulUBrQ2WmU4ChywSltS2vdddZE40ReykKoLr8wjb12HLxzniz3r1
V3Idv+2whlWrMlAa7+yhAg1c4RHsvdfQZBATMyXgNAf/VPVtZp6xUHuzh8BRdMnlaRAH9oD1Zcbg
IG7uDS6HSNgTP+jzrp0ZsjOLRncm59m1b6innd3zun8FaLQD1wCKlz1YxyyWrKvSYZq4HiRQVplQ
yxK4D0gjBA8wbGZOs6EG3pDXYCia5mwG/8QpN3PSvUnGImj3PFv3GtAYDQvLhx0LSthQSH4Jxbqz
CeJGr05FBAURBri8/d0zzXwkHMuhXwN20irGd/eC/sAj4xkeyuqvqEKT4PIEP/3MR5339pjSsHfn
wCzkJlEMBxao4PHvqvaJsFsg/fP8wBdac7lFjBGa3G3zwMsYHbG0B58Z5l2Yv9xVAz00PXtimrKi
w2qnuGrpnaY3EBy3auF7sQeylSx+4jauyXE4cyHVps+IPlZgRdkuahQz5oMdnTC/fnr3eWB1J1lr
CYJqcWBkerKlqUV8RDo1mkfmWu/sMAR3MGli2GqLxXUt+p4V13tdgITsvQ55ljEBG2yDC/3064wO
BAxjGPWKBUvZFBAz7sVJ5WeV+LSV6sSb3KXjmLQimNWIfJuch8wgaQecKWpiSzzddBi9ZD9Pq/Fa
jPvJTkLxWgR+dWbD/DMdI4jfNoxYgHj9JAi9N+n4Bu3qQhNOAII6Ak3B1lssFy8zxoGtdRuPjjr7
xZiGY4Wya/AIbBcfbqcmhN8/Ik8VWIrILwXCIMz330AXvOE5D5Q7BGNy3vP6hvtd0Z4BQ2+LbXKG
826oQDY0UZRVqOxTg8QaxjBeOimgtIcfvkdSD1NhBAjajW5dtnT5IIUEwEUj1tCcQ60cbCcrqeF8
FuGKVSfZ/x+OlgG6L5w6hsRDYsIircDsfY/FW+C9NyPMSRpjoLGpR8vxAwplMTXlpTgOv/4FyaFn
MZyus6jZLhvWnj1wLJBAkPhXgdgp2SEnAZWOBV0fuUv79r04PZC2D07yPjzMtoZu/5q6nOsCV7Vo
7ieJoCW8HPpYoxcZP5qiyXNlSUTyGq6in+63UM01xXayasHBFTJJFwQtNegyAcUtZkRVZywSPJVf
zWddCpLoMBVgKWsK6fzIh7wvFq2voHIRjQLaOxJ0yuAf3Qk9KTqIw0RzBEh60lg8XpZyjaxsoZ9x
GHds86CRE2mBHc/JSLdn2PvEihAJ6CDgnzoYL0W/OfFUbgXrhECwsn2EsrpK90BnQIguWdyU/zvH
D0hJBpAp1S5L3Q9zP6jOgHvHrVzVg2cS1YKCL2bqZcBt0n7XtoM7GcLwc9LQtGYg6ceQ5IIs5IeU
1ibi9qKGXgSjbKf76ALZ0OOKo8OFBwf8EWKtE5xcGLFAYAUctlVHWuKLd8sKOjFlaEPtWly9B7Xr
fhbhzSmLwa4nfP165PQCjyxw2HuPv5TboTP7ZqIKoKu7oR7DQQyeS/puEMoE4D1QaY7e1OknK1Jo
k9TuYdDd09VDNkkB+zX/AmHWXnTI0iGBggDTVgkBzw1+yoTgV6Ly2GpxMa0Rhs8u0Jhtl05kGtlR
Edu089VEupY6u/BzL2gc4VmxUM7Us/sYvG/BGbJy9CeHCaEfvH4UNDNWpRhq7fgSs43p8F6Jy5FJ
N+RcIzztIELmb5Rn0npg0O5I+tAEyedpjZM1k9utkbZfHUwVNt4PWiOUbHAZ52g80Wkb3+54ZtI5
V29lQKqSd5cfpQCC+ttFizq6ltdX7RruqwcWeV+AXtIVpHHNvA9kdIQwsnpNwhVq/3dMsa6FXh9p
ncuqZ9nc7ppdQZVJpvYTiU6NepnhginFhUjyJDEgwpoWY8xxvo2Qpp+fl/8p0tCMiio1QCYrIBWu
fcAPbb1kno1QAo/qSKGpe3TOyGJi85p4RVhk8opeJoITOSsoqjrFvAT6FfzTMZyjZWVjDvapXp1f
i0bYF3aBNerg/0aD8GORzA6x9g/qJILlJOLLzqrfQ20QYW2J88OxZ0zzigdJ56l+lyzJsIEa6fob
MlXIubnUAQFRhp2iTYOXD0CmLjVLsq0i+QkeBxw3b661qglerrjU7Grunli4q2ni3e7ngVd6JafV
tm66eGdRHAJNqYzBlLrKW8FHB5p2ZSGy30mjR9gVS/2MhrvVBjMwRXsvl22kzVwu6dONE8iTxmlZ
zbjb8FgoDiDZ1P3Wm3j4KwG96ErLJZvFBCyLvclfxHOxa4mRoih4oAsKm4C8ALHqpHioZxVe02j+
WyuEhVLxWunfQtSqmIEUUd9Ko5fuUeyJo9Iap80lJSvYCU7wbAXRi5iEaPZ6dvK2K3JyLiSBHZrv
XhE//SG/V4TsUCC925/OeEW0cP6lap8tr93ROnqBo4qfN1fTDmqjhKqT2mbIoK3rTirMQLVE4azC
oMIYDbnUMdSe2RdflBfWyfTuPArt1iq8Iqs/4JzArMycZau5HuF1yMHeb0/6qHsp6hdPrlxlMRZ5
++szQ2bsdaTvFxgh3Q71nPJse4O+CTtSHZ0HHuhUNpLj1elap8t5L1hRwv6eMJFyU84V1yKB7QyO
7WUYSsH6bXvsHmgN4tXe+wpcEEcgj00CR7ZrTC0mfcUXveRYok/sYjaN4eo1KH98pxnd/1XeeoiM
3QMHkqlyFGGIp3TihJFSkhcZUpbxvcqyXtXSG2lMK/tSc1ykslGNxext+BA3FxSFB5pEOcq7eqko
IeEd81WzC/b/0EgeEJTSvq/y+6DK9qmclaF6reGe8J6NtTChxRbq/CtJo/edrRvCixniEEHRV9zU
WU/HrEdaw5613G/wBIJJIVqyP2xFxLcG19y6d5T1gWNMlDS9GrJzranL/T+oj4QiknneiEbKKUqr
QK8/1Zj/9kMt9XnrieTCn4U0hIWF/JmaXL8+CAQpzm+RFrAuTC1jEMRI1bBqnGVcyAEZkpAJYs2c
G3XbcL+CWScqbHWOTNUjWcXmZJOT+GbhjrFSmb/sKGZa3FxbSSvdqJPjV5fz+YE7GFxoxcCwTU31
GNFQ0iUyxgMAqHxp9JToB+So4dC38agBt3Ggv3UnwZEoC2zb860sRTYxNvMxR5/Zv7p3K4sf/LCh
6evYVwzIE6Iee73cFdBtCqqT4n27EwUIfvrJ8SwUTGWVUBFVOTeVQUuGj8+VbSsmkJKQZQ7aQcuh
JjpQFJe3gAxiEltNXFXKbnMljQk18TQLSDi5fzlJr0CAZo85a6ICj0nwQdS6JfPKKE5++E7FzrEs
iIr4xsIHCtyXmYVL2B2AsXl0WphEuxbAmIy5sFVdtg2GbvBBhl7Bgo7bLBGGuWAy+OGPXCBzonuL
ZH7F5PJZDCFM2Bx7N3NBaNyq+eL3P0/ze8evjpz6TaoxW6TTKuhr62lCcSn+m3czk29t3Mv46EIX
/P6Wjzfl+SAoB/giqJNRp1w7cSbjpQVtDBnSQQSGCNVfxPPNiHFirvAAnNW4AIkE20dKaCeZIXGy
cwF9llMS4EXFY1qoZZ7ov9+0J2w/qlNy14Wk2fbybjeaxwK8+mdpBt6s6mbi/MhXSzUVC76b8tlQ
DFqVtpjSsXcneear17EYJv0dYFtW5BjloKQ4aoBkzS8jbY798fd4WLoddWdjSXHvjVkS26AK4Bwd
lViNaS6+XXcg/eaOaXktlRX7NN97KPLVUlpyJkcQuks1wJNi4yOkv7gtOPzvZ8YUwOwGRBoYyS0O
bf18bJ20Ce5ub4C9yBvap7JGD3mvlU5x6onDVXhB2UK9th4urTjQZcLA6ViF1SWUpqSoDr2YF23g
gTzP57SUl4IsemnyNimcFED1EPftZ2ePUbaUTeKmWbvoYV3jb6JBQ7mo17Ugw5aNN2rvb+QRAIal
WUfedCxUe2061fUsM/0mpbcu0WGx9FiNfMgbj2esARf6vWDr+QsRS6lAno5+p9SRDbJzSBh6IewO
Jrg6NMKyVfdHa/QH9Rp6bXUr+1h7VNQx6A6YUSH7Ya+4cM0HmeMivRrzt7DfSHsNmMrgMaUpIGFg
sXEAOB9tUo6LuA1tSbZSExBqjxYElMJMwrT9ET0XmiCeVL5qPVQu4Ony2XKusg+DIXHjveigCfY+
RRTFFov3ItrjsZ3KkIglo+5BlxJ3g0T3LdDyiEL7iRscfBIGGV0voiS1MqG8Oi2WaKmv8W2tu/3H
FFXnusKzSzM6kyYbNtzIXQVEFbLB/1mqy+gui5TZL01y6JML2bBizMt5nWfsMptOuJrIk/VhsIm1
k5V3grNxzS3bwfK1WFbCo6HCc/SErz4Rqbx1/zed4yVhuYh3l3m0bHRloZtA+W0QtcRkc7Bd18YZ
V7qUkWzExsWdnniJ/lHXrcN2HSG1H1bhhIDS+jI7P8Aorf7AUoTzsmOiBzRlWvsM0pO23TBnLZC2
pgG0dTKbzecUAS7Jbd9NRrlspu6angyaFTk7r3Zi9INopZ38+nZIP3b2vUyHpMkeAGVobcCXw80E
td0mnMInttqktUXOViZWC3qB+/P8xhsYmqpkrUvxm7hnRtasGhURH7w/78nh+qwldk+YZz+RwcXL
IIJsfM3LYRHKZTuL2TZueOBFFOS+ISr1gnHxUvi7zL+xqfqC6T4+GSkKkE8qGrwZpRhJiiVZiK9B
AHcHYG498DqCO3OyhC5ra6pGCuSXH4wdP2d3/o13/T9DIJ0PgPkFb2XQukj/NEcZMS4zybf9AY8c
Wy4w8cllEXGu9w8HRN/OWKqeIqHkNyEsNEccRP0sCywiRhQZp8BMTsBufQr8vth24CQ+GkIMjVXY
0QQrtXMurj1HVQ43W0Ghjh78SpY6QcJRyNB8pOfpTit/8Cm1XYRgIGs95AmZ3BP/H/AxtIo/dU1Q
ZAsbFuRhpzsa8qSo1e8tx9G/0T9sNP4Lh/vn6UBtyJlWsXAB8VJSaHjEUijgvFCH7w9YyAYRVYyZ
Dcg/n4YDjTXBBBjg3+8NfgBE9lcsPwzJry+rqQW5C5Gv5j5qenKT2Df4NXQ4KCk6fE+WHhz76noE
FPjHOsVOLSN7wHD8DI8eHtAzwoO5oWC4263Re4BwGERpWH+1RkH0Y3PllQtd8yReqAI666fOfSj2
Qikz8ZEwZ8mUBpvj71trMgGvz60x9ZzP2SbtKhtJN2JCYL9a5nCuXKFB4S69tX/z/gGTEQuQWjxA
CWF6hAzdpmni/9p0OcXMUUSmF24PCyzz80/+XDIDXZ/YfuNMysPalmQk3VGt6w07UuA9rFnVFfN/
sLaq7G8o6+MIn1kcvAotA3+3LxWdcaC3K+0FArNGA+gFI85VLEqsDCyHxEL0kXXxf1hH/XRz31jq
hGtZnY1Smv0XNh/Tznrg+HDtRVOOidFp1SjJgOTYxSudBi8i6+4NOYC8XeI7wmNRgDYztfC+Kx3V
nStzEIQn+i8hsxKx7JG23yOl0Invjt7UcZwYVVtd9cuiJJFKylIr4seQh/W6uYnZR4JfBd12evZW
nPZXb6uhRFYVuMifsawsuLerakkUSMzMFQ4pb9Mp2kn2wwNiDzptp1+9oF9opnEB37YKR3lEenED
JQGAd4S3oqjUKSOQ5hrIWMejUo1BaUsrZavkXX+BqSsjo1N/KDq/VE09KMbxkGQr+Z191O6+5PVC
gJdLFIVgF4vISQFJwUJnWOq8y9JZ/S9vHUfyzjDLddb8P0MYcyBr2qmsEseeFxP/MTWREcIJAGPa
CWQ7UlwWqOauyI8B4FrjBmS1jTKrze+UalaYCNuIrXSDNz2ugruYbZhnM5slei+wecEfw8f3VwLP
kR7qs91fw4r0fiLYQg5hLYfZnodHs5U2btRfQ+wx2e/uEABQS4xETjKzOxMn2tdip2ZJfs0YwWwu
T34AveTdq8kGjKcfbxKoQK2yp/cYjKgNgycAeN/dLfeObu9bkx7Kon1HVbVxMKKpj80u15FIla8o
H4WDNiuFMefzNnZo2OzdQrtKhiHvcYCvVAbASSzZr+rY8eG74r3Q8HOoKznay5xxQtntqRpBbRoN
Wd3nuJtmp2E3mZ0pjubXqLkzYfMFrGoL5yYXM5gG6RVDkggVqQWSpah4EcqbWmhbut+9xPBrOUhH
05Fw5PldHczt0BBk1WLrTEJd1jY0CkdJjtpJ7UuAUS63piqs5ES720IOOrlV7ifbwqUnZSsZpwnM
nGco7WvhjWEhJ5IqICK3hdQasnMhSoIQnCQ40Yj4/8VsCIfG9c/2BEifQV/wOquxWov3vtDOGu76
1w2vENKRFmzbXM/m4sJ1GqEqtOQatBk2+puYuMWaIVRL86T6QMrOH+rfioOVNfrD2+LzUExZCnF1
jvmSwSestb2PCDHB/7bM3+eijkE1lTYUuxES/xXs8qWXLWgSjN53cq3zoekuPySxli7TbAjkYEw3
j5T2ldchR9hlapHrTd5HpjPkOLprXI3nhENIkPwPLIFHkvjRRGcltFbLnOwWx8lKpdidAezsr1AQ
rxEenXOW5GNwLizpsg0Q8ixMMcMEfxqRBlpLVFUBa6tmlqkHbsABkDdiGu5zfpr/fmwDy1TQD/wS
U0cQqPYaLS4Trh8Q0EJ+fC2zs22TPDokfhE7nx1dwoHnph4Udq8tmIyYMJBG9E/tcCBz6k6PaUlS
upRoT28Mh2a1drd2jcxyi5coeIPNZdxpypVc+O50fJl712inq7/ZGRFOo13Ypwo/PW05t4aeqSjQ
O/MAfSyfVb4BYP+eViLhxUmvwJLA+CwEsrAi+xFgIBBHwRzTysO4MqRsAV/ecHRMYRK6tlTat/OF
NyfISYtBeAXQhES/3SIEyFS3Pe53BxOKOltLe+CXE33/GAi/wmmy1wsekYM2B1c0BdSb21tdc8pN
pR32q+fmo9xt63182aD9n0Isx5aUakdJpJDqrs7Ghu2kWyYfNBDWZjYYqsjBKxZrd8V331L3E1Xr
H/bE13mFtYtgJx0SFAq4l1ugzmirRRTI1ycXC7UlLbBbrYQrgOYLl5FvZNfURMPAJo3KuCgG/wIC
+hiPegOsLLA24oC3xbO7SrSR7yEHebVeoNKdverAZtn2GJhHFlCDvXMivYq28GEEYmvBY+fkj73T
3opNJMt1HBuCzgnyEYeC2ee5VqVjQNMAFYRcWyVXYsJ12jiqK6qsIRSBfm/rNjhMie4zOJhAS0Di
Sx2MKbhpzLZ2GtSZR6XGEz3IFHr71LjYExJ0JGn57qc8F0IRsHjHJg/ow7rl4iU/okZKKodWpOEW
uP/0W/51QefrAqG565kOWdpdp6/vCubP2vnE2M1Xb8nw5a85AqX2UPsZvW0e18JtQfL1BZHK4FZq
O6350npO3bwqrFt5dlshVt8t/W34AGwta807E55IDZId8/2SmcSV3DEwNwevpUgwPnz8ud7X3y/k
KEuEA5vdBfKUTbGRyDYtz2bje+e907a9gX9ar6rifJGLlD/WCf23OCI14jpjDHEOE/yUVH2gAxPS
sEDA7l1rPrQq8uv79AAQMr3UilHIq9zcCRnHT9Rn89BbNACuT142mYA0oF4wQKnBKXf1uUrFbZdu
NzKJNrLAQipZUh8CQhasYPOwmKrgX90VUhx044WVSpl3ROxW2k3OUhMleeyKC9bd8lIqoCVKn5FY
D+hz14xu3uCEWsRnFKapxw6SOkBmsRjOkq5mFZSDZgdPbNQiVSnF8e9gDM0MORY/iKosn/qu7ASS
DHc45iTH0EhlV1DXmtgP9aAqSL1WLzVPCYiSR650lk34Eglzl0o5oAetiZJImY/aUDVqdFYhECND
SXesv5ojVCPjZPDXBs2LomFbzZIbvJ7osSwl2M+0Zy6S3shiAz7FxgCNbJjjyVHY0uUPifDxbent
A/xAU1VcTwy4/Ta6HQPsoMu6f3IthaxuCsWUoVRwwzhbN4fWRnLKwtiOGucFi09oDDPHjF4FkWH4
u/JZuvUzPwsFZy69q6t/OZlEcQZU57lM6oJpsAu/y1NDevH1UCZ/AThX9OlFlRRIGA2clnSP+0MZ
15z9H9XFOBN53jsseCX3oDsMVcn0QrjH0YqvAJAwsYwkUT1LkV9es0nUajVzBQ46p04cc4BFK1W9
aIxAE0Gim0+xRkis7nU5iMkQNWTiSnsCLRIG3b2N1vp8ZrZob3R/tWeB7FQGGNlIyg0+ziSSHWcq
GGYEUj7NQRRWrfgOQCMFYO/L2ZmP0shBKXAleBrDxqdkLua6q2VbdnanjYFzFnO6H7WiV7Gar891
pKm8oCtz1Ya262TZ4p9vdVpZ9VUpMlCVwrWdP7dD5TjmXE7XIXmjBAnyW3EpGBvXivzqV1W7q8hn
9nqqg6uOCyJL0K6ppcE71rgELBlZptmn11diGLDBHRG/+kMbcS2RjMticfHZYoNktHNdZcAXg2CN
XPuHEHHiiKrKm6UHA1r+C0jzfLnDhIuzeKjxE+W/UVlYA6jdKpR/ZFeL4Q6n7Vnn5owZld8rQAeP
HFIQAaqg8UJ6nX96VkMXoujwGz/tS5VQf7wtz/8VfBuG1DQ7BeRSfAr58LKrkMXyuO/nGwfnAOZ5
fYWLwDOqmM2aCAsYN8bXNoQ/+ANx0aC7bV/vGcXI1gMslQKJIfJM4BNbIRqz4PxNlok5WMVzHauQ
b81ImpeW0FWLFIfOPoigvZPEIedQOvAPXqRu2PDoVuli9UApifJqYVTA3m+qXkINDrcIGrjLsyfO
eDw+l7ZeLCKbN9n+ADRIaUV1ZW7oDM9f67pbKuZmTGgnk7lXz00zvVm5WgZVAwLA3CY2cjGyV+g0
qSfOZuHU3+ykwC+Ce+Ba4/YHp1XNkn9xokht+DoUDY2amg+Ewq7hNGZNxk3O99IM2TQEMXxvhvuS
XBi9JuBYcKRhGWaZTIw6LnGVhXa9rXyJz1mnt9E3j7EpN4b4hzM8znsIKyS6NOXbhzyNxTujqji2
Tjk15QOviaoM1VYdHPsxiyGmHyNVstBPz7dkc4K0WatB40Wa14vG9b/BgfVG9MTbAoKnIHY52LsF
IPOWEavLAAJpUjUsuqIlciNxbu6/F4fmT+Xl13zCM/sqeNHdX1TcgHW539c3p52FlRNwKR+AGCpD
TglmT7He3H+R14H8GAtIiwy3QCyGScGPhGOhdeEOAB9T894QqoqzbodzcE2/RQJnlr9K9+3DFXD6
nFO/FYX1G5Ztf5g6PvMOkeXiFtSOe3hR63keATnvJcFvevqLKrHQ3KUu1kzmeUG93Dcjtz3rwpFe
ZlOgxfFvarwYNbtYfzK2g4FXaTBrX3NlFHeICqYn1ZzAWMmhTmIqGyzXtUy7uVehyvzAOyqB+Fct
r5SkhygB1tRdt6NalrXatzYuMjubTVga2VwFKlr6qjcM3zE7bMhdxGLnZ5hR5pGbcMBJB310TY6l
NpBHSkRoSXoVItqsBAkWViAbtK0oHiz20vRM5z0/g7lg5VRmGm5ysiH2ElD18ISLMda43dbVgnBB
kYsYD+8iNlUAkOQ4Uio5DxuGNYgWyOUWoGzcD64s0LkZ7dTnBeNqkDShQDtzjmgMxMq5C90BKvAc
ML9U5t5ea60rm/RxTtG+AVd6rWF1n2pXE7VNKm0HkoU8HwXt3f2FHXjTRseKb4MxOPxcqlMpct6D
xivMGn8S/Ra1gcKz9iSaaBCEy1+Ig95FDAXERh/OSXxjUmQ/IRGi9/sZ3NfppsjTF1YWh7VgLgJS
w5w1GDHqkWS6W0hMS/rd3hS7H1JLnT4XHpq9dk9q/vaQ069s86kBF3awhjV86mPdDksGxIcDNHRq
z2Oc54fRhSeODq8ZlbebZvA/zPz62dyDTzlkX0a3aApdIY4J179euNSHOOjwPW2r7/ItLeDYfAPr
9mnL9/XPjuoeRKcPek9vKkSX/TYbVGKH08zdMEHyAhhOAahYN2Zzrz6E9DXHBgcJCbT799gREtfM
MnbrpS/TJGDkLxYkVdAn7ysOacuvCY+j82wY461V6Sr42iOi/r5sbKeEeez66yfVyXq7uLXiqYxc
/3cTba8oKQ5+qE6F/DieuRXrZBfkRjuwWoBRUvIU6DbGveN774OIGu4t2BnQm1oJQ3Xi1B11TruY
W2B4hbVmXiWGxvPpg+MXUPQrGPTHliV4StbJvTx3WgyXK2vN9eE31uX3CioCSxksVmbNezERhLxi
6GNnB/9rlJZD21BJdMgOE/6VB96j7jElTmSo+t7KfH6CWoNm6hnpI9KRpkUY9dRBX/OZX/Kis8Ih
oUROBp6AiwncMZXz94GOuuqQSarPKwq80rn2fve2kayOPN99n06uP72SDUXte0o2qxffLGVdPirQ
cUs4rDGtvzg5wkWgiBPzlPPwIlYR/56jsXON41ZGAKh0tMgyQl7TZmRakra43KotOT6EjUU3DiaT
LGBdDWqGZ0Z78BYeLwioHn6oikZyRm1RG70zf9Ft1Qk1ITcO0TWycIP66m2tyvihrwOg+zwIuQRM
jooKR+AJJEH3OOD6qUK+uOl6GrzLa/n1yrtExcU5lub43/86tr+6mR9RKjiSrd46Y9EEVdvDElZy
3pYaiJyQ1F6sfdKWzzktRh3UYEQnRYxxjt1t2N1+VeUXf3eL7RlKlV0HY04SJGgK3xvp0yk/rQqk
2wGd2MzvqD9HDH0dbl1yeS1mTGddLPEufOQbzHLus9ZtE1BTaf1202Z+A4Nxyxg6xOmjVeh/kRLn
X+Tzd4VOHYzQmzATNXLLQ/x2DvY5WIbDZroYqSS6NP5TLd24iMGDgHz5mm6aayO1HQyFG+TcgH/j
8C3RCJNssyrioONiWyV+Xckh/ft7gKW7rk2RCrqWysy3LwPYt3Rs2ugKXMzYffsgko9RP7cEoKbt
BQU2ZEmpE7pvj0bMJm9TAhxbok1DoRckM7xW4du5vpr64pHzd9QQgMFK0SM4hFx8xE+2ji4yt8iN
BBFnQG2e2Hw6QU1nsJnKpogmDpUBuu2uuIydhiqDqHzd1QJ/MnfrwBaUSLqGk9QHoCmQ5e9Atbqt
pkamaM12NwnG2cpFRSSt/Q7+NvONsJ+HF9exCDHDMBvJZCwMELDEUFBZn7Fxbb4Ywwso8LJae9yw
tb8HVHKbOURm5qkTrjqaGxDc2nGua/VhASwdpoHTSUQ1ghUgkY2pmtzKNRsK6H8VNBHgWzELrwg8
p8HffKfms6Q0TyICCQn1+oitvyhItwkzz9/i0QaveG5Daoitg3bete2nlywiS5lPdgaMyVUnQoh1
zmbuaEDaD2K+CrdLF5Chag+68rjAXUbqvilUkwZGmveX8sUhbE0ASLXcYp23L9oJmJVeIPupUPMH
ICyZf9W3rNQkb0v0qr9Qu5FiWcqjzfJF4WcwsA/F1U+DM39FUhTtJWoQXgrGmDiWJuqUHdyr7Z91
9TAMR6i58jQik231GBWORVFyjE/8nRqRQRIpLb+qUrU48lQlZF8NUd+skZ5budKrpObfjeK/lNYf
nE/vqMtfUyb8KJNQUwmMXqt0xxqWF/K8hnDCGa72lMG9T4/t7ez3yoj5Uut+knSMPArRq12JiTN4
xRPoWvzXXlQT1sy3GIKCMzuENNjzW8l09BHn2MlMwQK5sxNm0Tawc4d0TWwegmrU/BNnaF1eg7Kc
57arF8qYcrCMUs2Y8BIP0agCZXiqsCBNHA24Docol39gSRpyHHFTxZNNvCUS63xgZfIAiliw76YN
HHhwpyxtqfwTX2k+YbSXUL7OkUNGzo2m3EmCmxLF2YdAbFqPe3E8SLFTk7GP/aZst/wJhjxhOk1C
K3NpkXUm8YylNqQFVd6c2XqdXuGPahNToPU/Rf0j0skesctNJL0hwLyT0VGO8UwnLudzGqkxOzTJ
bjOHrQ8CBVdfbve3ZHcW1Eso7GS/YpFc3neokx4ozRPP/vh5LnucoufyBKbzmAsTQy4lgZEvEhvx
Xlop3ahkx38jeBufkoPEFGF5aYg0SZG+wp8j5AY3Ohxlr+NcJoeibdrP7T5yn1Yl3V9eqlgfzeDN
f6jGgPG4xpMI8K5J0UEscWJc1KjsgJKEd2HfFY2T2Vmgz+K6aCiZ3rJMKLCjmJlYtp0hGHby8Zvq
FCoIJuYoQzg9XxtovgpF5NFWSwXfeOjTgHHIa5p/RZv2WerqymcS7sx5XXs1VhC+xFxMBwuRfnrD
2hcL9iWl7eYAg5XqsJA5FUKcVQGASkS6DZ01oRc6rcO6HQBGLwAuWQJQpZUNxKf3Q5uhAQP09o2f
Tsz+574Jwu7De1EkVhSFrRIIqxzbg4zLrNyjSKpKduNxO+NfmBvcjQ8J4dpOvgghNSixP7xhF3J0
x+9utJcOwtqvWvVolqbfH7jdYHUcr8AT5p/jgxMJgo53R3/pcRaPn4OsVluCo4lOaWFCcIL0oYfn
e9Kx4/3dNQscC3Hg0cvha24GaMAXljm86VJx3EnRu8F7o/IL4D6XFdwbxs7djrZDFiK9yExfUxQh
8CaJr3jguVmyAH9Eyh2we3obRJ9Nnv659aaw+S8RW8qCk7pXyJVi02Yx/Opx+W2eigz0V3OXEySa
eKhXlouw9alUF3OP0r+D/zr8V0JFl0am4NWQgxz/ERHv+Vk6eMzDlFtme0dfVo/VJvJjAa1Vb5wQ
n3tOXmCzthQSrdHlh1mo1WaD2sHWCIsU5zar7tBo1/OsEoa+ZWX6ziwOIj+LdhLMGaRlDpOxD7xI
Wwf7HRGWRP8LDbFpWPhescFIXvEPMiGSpfPzuMtKLenrg2u73Mv/O38giqwo1zbGbmzKtoqDX/7k
gtyEKedGcA2rfJaWrk9zFBXxpgjBWgHGgdaAKpgqpRC+79dgUr+pUgVC2jW/GHYcWYeg4FEsW5f7
OsSxAhIRBgPbBi0T6Rj+uVPoXTVGP0O0K1lj/KrwNpn4BH9FbXbukBgz5fF4enk+et/Qn6Jkb3Ro
yvxoHgos+NMID2IgYrGh0J9rstYp2xn4GpGHx+010l5gj1aM2gLs1I3rsC7murssOPdbSPuyvnaM
x5zvqBA+bBNHUTq3smc2DpJpEWwutdahJioqQGMWwJyPxQZEX6sxK7/bSJauFZbUovHFLV4sKx76
93c8qpxiLpO+o7IgFjY3UdbVossycqGOVFzSaD58J/Cg4MA3Oh4Ir80ApgveBD8SCzDB95NcLZkD
X7Q3A1XOPBfzoSf6yqugfgK1xSlTcIGx3W51Bl7tSqOj8NlOA6kdHkTMkxmj9+RTEad3j/Y3RG1r
k8YY/nlZgATRtj1yfRV0I45Fni+QvCRz6+5YVmvf2uk8AWSYA0cA6Md5JCNXnprF+jFMeGaYqSFw
sMjUPwhUumH89DCwjovuAv+mDJtJLJXsZli9rl5nFfnAk8gn8aXxMQdOK597+5Nygl+gB2lnO4gE
k5/M81MfxnIkQKadr0w4sbUlN7nQOU4zT4cx32qw4r/775o0N4OD1BpouV/zfayXDMgu7sanNXyd
QX+HkftHntmFkJuN2wK06ZsRjkSv1nMwZ+J0PEkOY37FESecPpNVnwefMB52D73xZm8nn6D7NEz8
O6eEIAtdAmv91s8ewZXb3yqDxMrIwpgRpwtWbcZC/y+fVAHc4LCQBMWowftvgGOx7fKxKzdglZ8r
uIeaxyLVCPE2RFRz8uGmfqSf7HbrGbtbF9/8HKWsK/7iTIx8gsG0T0eeME/h1qaUhGF32XOSUfCo
aBnLe4n0PYKPrnEljFZ8HOWQC1g387yfF11TBiQ80TNVOrIaFUi0vauuP7H5nuwKyDwjujWgsetH
Skf2miCKiIPi8NdQgWupdI2Ka1i2hzRO905ujZInW5UJm1NYukqf76wfp4JmTQmQMI8Irb9q1zHf
HRzIPOXhbLqst0znqYlfu2sh1Wf66vuOU4eXUxxTQhD9heR95oF/EBuK0fzqLlQFKt8CQlRhkvt7
6XiYtwIin1BOj5BJwiVnxlzO90WQE+QuWZfk1ROf5mAu9VRUU4w8on0688T+vhBCeFXXcaND5opr
5L2+LOGQd8A/zVtiRdCCyB/ui2V2ykG8OA0SNsjus2SiPdVH1IE1c2mLrluFpHxsJydWgw+b976d
HaOYsX1j0IWnnpC2LvYQAdZaoXPCGNNiYG/W/XVY1V0eBYBAqls0pCMUWWgnsH0w8UqB3X2THx9f
iKBPGj9T0olrSzZbek48TA068QkA2qt5UuKmwmjXwf8DguF8Y+BtMkuVRWlqh7KslsUspL9a8mQj
dWy/RdfP+tnClRC7l2Tfx8w8Xb/7ng65Vt6zrfrdNbO4muyYV7i4OLd2fPE4ECiW2dzAELRQoB8J
8RbujFKQQcQQQHLZ+DSHVpiB+yRmuaFBUjXHTCmBZGM8tMlmJ3X0E5JbCQsFHKcWlwp+/aITUNIA
6b/xUuO1ZB47jPQWZlavRvqjyR7xCOIZ7kFeE86sJ6Opi+9cCmFuQIv4dbm/WhBYolM5p4aBLuAD
mm+Jus+veOcrtIa6QiwxnARPCtNbIa1mIW5tKYPqgVVlssGaTaLRbtC5to+UiVvasCUtbglZEByX
jPa69hpIcbgqnlimepwMo5bIIS+ZanGqpL+P72ngALxGd7IEq+RsYGAbqT95vChgMa1AfgDm5+E3
CuuPz3cxUKJeNkMkH8ASEY0jwKzLlS1kYMH+yBMdU09pByzRXSGDZPU8iELv+fI24dbWeDI8GDxr
BM0SjXo69VuKYIZ+jY0Z/EniXyYQ2GOp7jB2OdZBGLn978MytoquQsnSoKoXPvA67f5ILl7Wn3Qj
1UjztvkCZZISSCO+mpZVMGpOItQ9R2eK1WbucCKDGitHXiL51P0DakosI6X8bkT7IIZs1Xc9XJlI
7Cz9tTtahqYDWSbwuQlY0KOJRoj3rilzSu9K1YHeFfRtfefrMqkypOxXmROVICcHHzXfDCk0fnu5
Tqcda7djwA/lmYaamdeYZRevo8XrVh4LIOqNVRIH6ol1AfUSoyEbKV6Pz26LU34EuWjGf5cdRftt
HM4IPjN4G4lAu5GbRqH4lMfVD8kqJYVf0X1tl7TlfJMh+lcD5anUlYfpGWTrpy3ieKmUmcOE1grK
tS8vDU0zVIsiq8FsG2lq40Ik7LLFdbAwdIX0FsuuJCCyOkTK0OP+RccBMFKKFoTE6KQZGwDAEMvL
at/CK2BxEAzdiDxUqhTwKZsTSmoxbYyW21JIJTbZ9z5OEzTqxHXeU4p4dZBoYQdPSulCB8RxEu1c
On09AZ9Pa7GT9EWswgXKtw3Xp4LBLBg3U40zEQaiMM7ogog1D6AhyZs34/4gVxT8hcpqu3ykp7qC
tjDInyKHvRy6JJjGhcS5YtVbBmEW3XSkl5r8VhsFX1XYvAUxG0ZcMj1cVGLhhAN1z6mskS0zqUOx
Oviha5SbO/Lqc1s2N8TCeTrWmQmvR3JCNH27iz+2uaoSzRojolTGdcmMVzEAzStOKLoHkqEksrum
pLMcOXEqY9GtmwffVDYS6vktUg8bOgMn8tbfWlywDiVyIOlpFZmcb1nOjXtPN4gxVkjaFhfQf9vL
FvoeYddfQUDgc5mYHK46yMO5miW130SE2W/wzFDUG4GlpLzqHqHWHfmCrET/MD0t/I8VDW23NXYT
Klq7u6QpdOgk3pmKZyGphXdwL9Tbr2l69y50wVc36feU2a1hGMLyqfq2giGln8prX4qkCfNr2Gtp
Y4Um8p9Mtq2KT9XPsDQ5M1B57i0IlX+Oh81bzx1RuOpZaL7kAxWTJCmI/VvUddTUKKLOxHCNnE6c
cYPApSOXitJ8uYiqCuZe1ACN71YSFZ8tOFTZgo6/fnQHEczaORW0gMZrflyk/6t7MFAqvg28m20S
uu8/oohUqDjv7DuDxDL9T5lh8nt76IOdzwrI20ZhszrCsbu99zQ2atb8uBj4iu5k47r7Tyr20jxn
Fjijz8eD9Kaohit5llPkm5PaBjEm+wJ4Cx9Vv68JnyEG7XrTdQ+LniPTN8E9TbuNYP9k/gey3FcY
SAiywAaBAyxE7xFNZF83/cEZXCy8UXPaqV6kS2nyU8kB8bGld63WAokG6feDe5qFAtBpjgdh2zU1
WxqTVNmImx89aoELjTBPHpeNRWKgHie8W6dA8OnIzd//3pD4ydXyb23BZrYcK9sHuqWbMPcrG4FJ
XgRJHiN51P+5hQmku1cCsk1UNLTLomeigr+cZtlYDcZXsyvr/3HNUOit60a9q823XG2Of744UQNk
ZFerGabfcfVWEjWXzDlE34wopfpjAkQfvSRpM1Wp0Lqvl2/446aJjDEIdBKMhSXomyqo8J48fQEz
1MZqZKqFl41IskUioy3HcSoDqERqbjFIEuuUHHPdsq71kgMAlKlBCLjt3VCo4ZMAF0ezWhZBQFJd
lfsDpb1HpBWig/nhT5kol+QMDb02glaQ5Vyj1WoIfYyzWlFTtmGdam3Av62Aq8PS354vjbiUrIMc
IQJ962F2RuSPywb48ydJv80rotM7H73U3gIIZnGJTLUlBLkgw293iO2ObHEAhrBW3Zi+qPCwwESu
dYLqEd5VifLlIsnio2rFwCvCmew76z91qFLXoUga9m7tNv3+wLtk6eJCWiwEThtonrpKDDyM1yie
VRP4NT+Inz9mXT0NK85xSfjti2kGgyhA9ZK9JnsZrLtR3/dOfkOBPqvT9MyM5NfUcvyxObpTD7xb
uzKhht1sw0pI2v6AvAoojnm2zSbeHjofGGyCssC9obr3d+p8pDtEbTZoalE4W0LKJxHiBQ/lOUfP
dzDklsmw6WCqbHy5b5KNm2BWj/U7B6UVVlk4BShJwcgl3e/m8EWg2AcXmcphPX8KugCeS6f/uRcq
b/tn6tdWGeyjbG1+82d+IQ+KY1hXBQuCJtQ3+IoPnc2EHuQ3HTj/m0Ny0gRGarG4EKTTdnbQKHbw
6J78x4Vuof1a7ckBh7sV2VcqatL2EtJgYdDDoUcS95OoBmUx9JeKhGkjoY9wOrPglckArT8VIZb4
DySIJ+sq9o4ysOxnHyXZhn7NiKzvXU5nI8txeiwmydK6IFRlYofhEymqVthbuvAJVth/zfgHGcu8
Ke5BOwAr37blzn5HuQwqRke/Weo9dGwLJRIoMrsv/SuKxpEczeEHLeRheJaGWQ4rMOReQTisCPrg
TlLd3GiqZbeY4vBeDQPXJnI6vvdvBsseZ3sGq2ORShxyN2sPMSbB4upPH2tNJ9qJZgncxGD72xX6
vOwlR/4tpUA4xE4qsefJSRr1FecdDIZnNwyDFqWU0e4feSfO9tcj6RRbpBow0e4psi+Mwq0rcOq5
y7PcKCLx3d+kbnACTRelGD/S1mjvJq65+gV5BM3zmpN2M74WQy+zBah/s4TL28/JEp8ov7g8E2UC
dQv+2dEEtxkpkfLvMFoZI07Ylo2maCbPEyzM4vdTuukdNmCBNXqWt41S8/TA6ZdHSRLVMMZzF0Ac
2klJhkPf8B2tqi51OMeJURXa1AmWteMZEYAp/PszjO+S2OPgJpyQKhjvGVFfD7b4xHAwjtY0Pn/k
7QWC6wNjBEhzNaKxAFIQUpOTb9tbeq+anI77lvgJvPUF95REvjOKdFFuMiBLfg4mEDFhQ8+fk8XP
04CiLPGKrrp0nU0uvavA6wMQ3GDmklun8+7b+A/Mxfrl8eK8KKa5TtntVebo7ObEIqcC8k0jkpRb
qE7nix0EvRPkrTUkKb9TJLBmkyfF2oN8UxbhbFr8T83jK+NG2YNjzDckksVKqIIIpQ+TY0OkjECs
pGaz7ym5OYr0mYDDogXt4JsHUjKo8uvbThgM1O91M/k6zjodVzYNAwRgxM2hIkXLd7szffs5jYrA
xBWNuSPw7yaPeAY/sCs9RB4KO4LlL6aQrq2EX+jPBN2vO5fHDA2rC29NVgaU6MOOtu6BNdCj7fHY
CRz15AIV/rherHL6SN5t/iXHdpaDwRywL364PtVpKdblzy2Y7NGFu/ozaToGuiYMZGgttY1sugxz
JXX6xzGYKKTvS0zhijhzgOFiNOMYL7KDtKynmaFO70m39s6tuOAO+hidJ2Rbj0NDGMIBwUv9Rxkj
JFwsa5SVBjNmhCH6JUuuBSWTFoHoYBnSHHAZnKcNJw0X9X1ELaFSyF1a7O8OrqlvsZbl4VORziWV
gQL2KBAdQXzajRsD+sIuUAzcKjDnP6I4i9XYfeoz/iZhYfjkIQU1WIx+vRWtYJplieGgxy9ZpgCD
JtU098FRDDFDzevefLU49fibaZD+8pwVgptuB/nqfVZv4eHIfYUoGJnwhc2Z8gSUN3UMf0ugObvi
IAD9jR4Cfyql+ti6qYMV42VjJJbqCNndaNW2kJ4PHVbYPe0i4xMP9DVVEetjKEHtXAhEoTMswwOX
W5Qm1VTeEmVMFcx3g83E8xpkimwJ2kPs+m7gfwKexETZRwlVFW2XBvfiU2umGIFLr/tVre7iJ36K
sN7TVon1omggcGgs6scGgj4hTnhkNB1+ZpyI5kSYacctLEURgeCSj0suA7V3FqBOWMZBhCCgpyh2
300yd0lxavTivNDUSKvavAwDQqOvAnwOHAgz7p96ud6jWvtVd45Kmx3XFqTDfRk4NyxrDAPuU7Xq
T0tp6milYAZrabgb/zl+HSExga4/wRh9ztXZFaTLnpBAG1GV6/IiQgD/1gGBdi4sYVi0/8WCX5Qa
kNrRGvHcRorXL3cc8yCqGw4cWmIjleGBovjmc4PwyJjazsxrLcK1ZmCcsxIc8yodyKMX1GvgR7aV
VV1TSUmksyPY2FqxRa++Xdf6V4yE5G3qPfzQ2frj/GwOhKhnwESAh8ygzTsbLEWVMly6GAaST7Wi
NZ72cymTOXOb7VEW+WTaimRIBeOrNL6L66+0kJZ/bc+UWYsHLNi+FXNyhPFcj8WaqlaT2qrBDDEq
8hGmerDV6I68YMg1qh2sGJzuIy67dEgNzwe0oROevDQFaHliumXWCBCjArgfJV1rYNwF8PIeA8PH
7m8k233vCXgFSXUyWuwwVyOecXK9VwTsuy2GZ1iS/9XmEc9rzMXqYXgV8db2iGBtiMbCG7EISWQw
QOigAKdzRNMj7DBz4d2dJtDRUqJ8dNYy3mU63YGlRzsuYtkMPzx3z7XtXmzmnHcoV+WMc8YaerVA
CGpqi8FFKmealMVmkZxrsieOJX7mgAtSakFUnuP3UzK/reI+pbOQKRXwXGEIOj6OellrmZEsxZLS
zvI4OH5L0CvLB7baG4AqQQT1QJMjIaN01s98TZmGyzVccji1TqMDkNP2LnxQKcaF0sm/Ss/i6fbz
38DGT3mv+RuRpUf2fcyQbxUA9xfYaSEiEA13kAz2R3Di0MKFZ8IWmQL08uuirFij1y3bUovdeqFB
Yq7FzT6MdL1OnTdRIVinK0GjSqKn8HVcCwk7TShlBYeiWWrqTGaqeLVXazwdEsdY5jmF/BL54MuG
9wQ6l7zzAKhkCr7vEvJGRIrjw3sGqgb84T/RvKReeSZQWFP7ryCi4kst6h+Co7/uQzxkV9nvLho9
rpOJg9opvzw1BhDSA1UNXmxNUZQGM5MuY8OJil+rqoSthXbKMPd0CbzjT2MdAibXysct1FeJES4E
Fm5ROBPh8Caf0COAIh6BNTbaCpPLpXhtJTYj+iVhiwIhNMXb+Y8hP6M92RVQ481svaGJMcyB4WS4
XmEBNPl0fbGv9VQI29HB3S0na1BbR9Ivus2wvlGoiEt8fVwhTT1rbTVem9ZuSf9Bg6hzbtEx7Llw
J5TkyiwNK/bCIW9gqbnN+aW+glJ4MuV8ruZKFRkIIRdMBnPnFxhq7r1FwS93Qdmwovn82dS7444Q
0zvHaqee1MWqla4KM6WaeYNdr9MwNBJTfzTfrb3p/cOPM818QMVzuuFPuhVhJohqneQKSxQPpMYb
2N7uF5jK19ZeWdwBxLXYpZGW4ikIPlbwq6h1H326kRsAFNIQ5931OeJot8giDW4OGeTFxh5MBz0n
+8OcALXLpnL3r7yYj+y7/tTIwHxGDckI8Caeu5hPBEFjeGgxuwQALu6Wzoxq4cJeKuGhTxA0fAtL
Sf2thtSdfPF4E2ACUsHMZbfI1gbzabsh053lxJsig4eHQQymlQBE1r5gPPRn0Ky6xc5AIMfwI2og
vLlptAVvXpPb19s/HrLfF9A0Ec23UkgA031mgaZpXU0qhpF+dS/S0k+HoKMBFDZmyhbZHmm7FMI1
I4O9vahwVgdj08F8XPkBC6s7NLGzeakAiMWcTmG0kzXeKSkM3L6xTS3eO9XLv8ZQ8/uyOlmmfuDp
icu/gkakFfcViJYClU0cR/ogRpMLk/EqYG84U5YY6nkE70sqTbm7s1xkWY4SZNwrmXO2voT/cKYB
/xYtgwNIKFkUxUfLRFbDIzaC8/TWTGcaXo2kk0L2aJlhMKMhNESqCEmZtnsK8NohbTIgfOrz5AdX
CzMOxNe6MR/FIcS03LJLXSkr5xMW+PcdtGT1tXORjJ4apCmROB98VqWEQH9xcy8XB6AeN/t8Oc0Z
ICXON5GQT5kO/3VsE9o+zlk/xV1Y8sRybOfO7Hn0WdwFrd9kMgCadj55PZ76lSrz8D5TypKNUfUa
+ysVRRW5AD65TeJR+imfwK4RPIGebEElhKVfoNkOxCmcQiK6b4Ur7pXOvih6FUPfw5/qQtO/uV04
IOzGg1U5PMttaCPT1yIh9SBJFoE/FJUDd6Z3YaQYq9HgNC7Vzc3Py8BuDjDQ2W9A6uYavg8cb2eO
mrY6+nQGU0q8m4Ga6wKOEha1rWzaDV3TUXoT2cj7oBGBYuaqicyXdpMCQgd4x2TlTvt3axHzYihT
pW0LaHG4LqjByZabowFAZgKKQ/QQ0gDwE2LFtj7OtUEDKjKMbl6thbVFCm7udCadyDmwZrHr7JsG
9RRBLEyrCFfg4I1z7q3hV7iS0ITk+CywhIXyC+tvQ0pIpeR13hAlZj2HxbP7Djs3VXPGVenv2K6h
K+gTLglXBwpl5mSyiC1/sAwtx+WqCkbO2SKTly2TOvdZs59SeMktulv8c83MFHWV7G/44N5mt7mL
5kIEzlU5hctSLL15CLy6GqRzYeoxygMlm4JlV9B5j/MIlQR6vI/d4H+Op/p1NILjecQUGVrKWpJz
RDELTWmHAUwAfm6vVHwB9ZFsTT6GOAmBjpBjXJhKsh53bZnV+D8zVfGyQtOWhgYrq1tP6p5s7rQC
Usoj4IbLe58dWSQJFDP0LZaCK1z84v5OFF+ntcUMMh6bLnt6iUKLgfQlqpv7pROPrjhVhpBBin3H
YGZ9FCSBbWWpFJgJc9EJTvzwr6Mt1Wzjpe6qfENV3J3NEjiUjlOiqkMR1VUdZ0uUgociytGSyEUD
SNlAl4TCUu+GaaaAhr47m9aR0yuHgil89G6FRki14eHb0o5W3z/mWrEuEt7WqyvyvorGcBwMmfRT
++dejFUEMmqnrfwfrvO+/pmcSoOD0gRoQy/LhnPVkxwqWthm8w4DymrL1G+CCpj2WgKbjWt4OFGa
nzT2MbEFA9WR7xRvuwP7wBz2bFFerJ5mDHMBz1jiozmbwHEDAGt92pe12LEc08Egsl0/DnEZI3U4
KQPfkyxFCy4UnOxwf0sQ8HU7vkhivE5Q/pHK0Z+ThXteySnselbf1pw2OPrV1f7UUw6CWni3Mce8
+lPjtyF24K0DRhJIHd+4PwBe7tTYHtIXJiZC7HBD1fDUw8R8ACmAS4SA54C1iqCSBVz3ohwX8Y3Q
9MI9kkgCkCkYk4Zl+VqqrPwAiF8XiojpsKuR0xk3h7RsWG9nOc89xJqMrKx5glgQO2RLP+CCMRWb
Ybprn0q6rDCYNTV7Dsu2P7d+b5HYQPCmXG33J5N6bQkHQ5asLeOKWJRa5uEwN4soXZAEMZcweFkn
G7c8PAQdvX1sygf/Pg6z/G91ibXJX3fN2M0vvdALXlp+nsYIYK5tuNX1g4MQQbQ1WUwEHx8XwN+T
SqjPxvPSJj/51YGzdjtSGwtISH+T/BXvcb6OXSlAHYg1LknUlRfQ7BjMmeMTWtUueNlAp7iaGpr2
VYK4zecdbw5mK80Sijgw+7WBvjmsj2bLkEumSj9u5knmVdf3DQ0THzAUGDT34RWbY4sdmrCZKFzu
7FTOkmuooisQh+1dC2o93WyFLLz+AciRgZsyuiNWiQHNAVc0xNlfs1D8GJ6d5j32E604Fphjc+h5
hlEfGlQr6Cn2RJvVR6KzBZP76zBoIEtim0D2UXO/7893507zv9A77wg2YBmMElgKOqBeq5VI8Rt9
HwZqn3lnS/4+eaxzwIa1qZR4nVxMFb5HRW3toZq6m2YHUyy4ZjeP4RriNhvUMecSqfO3lTHy99s5
YyZF/lou+3bnCW82wa0BGCW4WT/9Kgv4b79B7nXzqIZIYvIiO6EELj0VOQw3OKGKtugDRrsha2wK
96lojr7iRXYSE7YoLyvA8WqamGxVxAJ6yoeyNyiry3374qvfXVBZtw1SbUyg6V7A9Vo1IYVzEP/H
lcEwhRoTPKM2E7qHHPz7v+cbWOiVak4cElhs30tCbBUUwGiHY7x9lCWI5b5WVH/v5T11QTYmbfLg
9lEdC/0D6cULnmlRn5/n9/gMf3ukJ1BpsU0fP39OY6gOCVJc0cke1v4phxD5XNcVHraUaRWg/4XK
gcVKDaTRfNgfhs2MB+77cEbz8ofIJos81cLNYGUhfIYxb+PtR3B1BfUL9Fo3IxhHuUPOnDZ5bnO7
sLU0gbAhRMOW/wiQxBvVsXArqmaSY4yTC0gY+ANr75C2fwotVWJYW/CtqB7aF1iy/XUBaxTIXKMb
P2hUaHR1bfErH9/zRzeNsOzRR6wKpODHBTPDst66Tx1lm18gNElrR/2X9kzlAKWI+SBlxv0CD+Tz
kQfU5nUCSn44ZRhCU2W2GCMrICZIFbTHGTYUWDQAoxDL8dFbBZp8pNnFLyabOgKVp3pgMbg/n5dq
181AjJ3s/MMAuEAivVp0jdTZMeCBP6TmHCK3TmHKaE5oY4mZy4FU9UqbGOj0qe8MO1yywQ8CYCVz
MjQlk9m8AthQ7NHkinsymhbUanX6baE3lW97ij07wz9a2uirVBCmJGqjZyRL9q8dLK1OwmpV3y34
StkwtOHsK5MtImRvaAMNKXl//F87n0N/69rILAEs//XTuSHmoewexRvPVRKVa0LPGbh/KAdutcDU
vN3SiIjGlxhpCYQDasjUw84kU7ouwOq0qQFkSevaF1ZYvPQ9Ru7i495gCA1iXeV6xNUDCKXmUbkO
Pi4DE8K1w0gx99xaSRjViE3ws1Ov0Lp8EyvBzm5iz8QHt3DNBCpx3wSJ2TqJkVaUdNJR7v0oLSGY
OMeer8CocAErmRjlManEUkY6RZ4QAVK3DFu9IgHVWzTpWcJ33u5l9A4DcAIS69J/fZQ8+QrspQkF
AbU00eRUXp29Z2dY7IBAtunmaJjyeRK+4AB/RZ+QPQ9Rs1EKeEnyMW4nrKD6UUozTG8yyeWUStGG
0Ve7uRYpBJopwJidinbyyibh7Ef5SNm4gLz6lMNQN62EI8FBEJnfiUmTK0pwLNCF9KDw2Z6stpbG
qwJix4t3INJ0FO0ExmtksXE0+Z8xYlEw6u4EsMXpkxEBXNjIxiGD4SFPfkGqn38Nvn5WEjdgFiBO
9BrdgdcLtjsDp2eFyyB1nXTmtWLYUvC62oKZYAZCztQOGTvoBCdPX04SGmVCt8gCxtjGwVnTOXTO
wIzZfy8gIAVbfFenXZr5qvXEiVku3lPEeHhDo0PAnre+HRfXa8laB2PxyZtjKK2EvC4CRDIRZ58N
tfnXc7gr7MMj0MT8WAMaiwPBniYLVE2CrpkxHjUQfuvZvxClfXsne3UbUi0uyBr0vJMo6BSSB2AT
RkV8MfdypckwzLd0XSjV5+TH0UNU8Jvi0NI9JOE8bLU1YV/HiV25/lrGWUBm2VoIBzTw49OHiWRx
ezbQ+n988+m6q12YSDwmtuo0ZYs5d159j3O1puOwew1j2aU9Q5Hlq56OVG2oWHaR1DEf3iqg+4Rv
KNE85lKL41HM8PpeRjG3p7tN9okV4xaK26fT4jbBxk/3Iy+4alSd6iKeiT1rW73WeU3O6DRqZfpE
sPaonCjIhFMBgPIeMK3TkbewsLjp/Fdnl86KoSnvwD2IOFYU54SJtYntDG4IqkV2KPfIfaMDni3S
PshnUfyDyvqwawxkTmHnP/jEY0UMjnkmac+w6XexhLytL/UFhfYXSN4gO+htdC5XYf71cmfiBNGm
yVa4goBSCnQKmI57fjxriQW3eaMC3g/c1YZ2GDFkJ44T/+v5cLMtNl6c7wTw4m+KC+mTiDoK76g9
nqMp6aachcKvG+ZndtmWQPxEvJF5/AgPAx47+HiwAFPmIAGTLhUHkOqkFvsovCjyLw+El9Ls0GD9
MtijT+knlVlTE5+fLVjySG6IHeOnFbJMyaN9EGgdaiDKHZm1kzWmLJZCi6QeixUBgFjWeod0u2zw
/S2jpwou4L4nGbjFuTHq+o1JhTWbAi7ZfwRe+rM3jbM8z30OUPIio9RV7L35GMBbNru/rZMUoKhc
H7RQE9PNp/Io4TwBLuR3jFMRwLsIl7xHifZiHUygeiN2CcQf6m4OF0LRcKLRdJkeQ8O/q92n2b+g
u/xBNwbamHVEYTaRgKm0eGuXbjAybpU/o7hYTugzc8qJ0FctYmutEqHJpmDE7J6gGV6+P9rkH+Aw
yDfDjcywXqZ9YACmB7apK8oPlPS57CAPdpOFRxlotIWKXiaqSKBi4iA16vqru0VB+Kb7H0nZJBgp
jejVFAsTThgsMspzOszeJxVaJR4iQwK/PR4jXae4N24XXBbnwr371EQJYdJOZojjWg15WloZ/kUM
UP52FWgWYiNhyuNXE++4t51Rbt6n4Qpe1ZFLgzsAdQIE/WJUDqbrWc1BcxRYGTT0qd3ZWfe6Pa+2
eD0EyInSH2AaxoXCKG5yXTVav7r8udYO9dS7DYMn5mry8bWgOmHfMuEyl8SEgIoVt7np5El9lG6x
OxRNpKojgCnmQCyd2ZpO3u+i27qc0BKlTdXwg8kql4/wu0NgJ7PNrwCGvCrM//mIBidh5361BtNw
c3E2skZ6T313qqFMwvLu55qlWoQnEn8Us3pT+pzzgDLA2IKeh9PZ4QNz1gPNwov+i/Bj4HdhJC4A
7wuP1vdjn67nO3nTA1ly5sWOo9bn786dJ9Fi9XA+zgH/4g9dpvosy9WHZvtBzSSDoCHmDAxT7Zlq
L29oNfKPfc4tvII5nVjv7jN7d0JJELPVSV9fAITLEz80drMRmzRXbZ21QUQ9UMIDwcx8r4DYD3Um
1/WPhdnv9ubNs3w+EUBILXUdVUuP7yWcUpzPcsi4eZ5wEE/QkEorImwUPCFZhp9Bf/lPVIDnqqPC
lbJduqI457TnGeF4mw54N/Zh8xTzYzRLlEsUPGcZKtQyY7rYxALOu1cRZOS0YkMbeh8z9anaQZ5G
kCbXsqRyUF8IbLXnzuBcHSjJQ/ZN4flchY9G359+UWn9adYsz9ZN+BLk7jEzKQzHPwJ3jevu5bpA
DCl3GY6cnwUwTRhGhmuvCwRzbcsoF4ywtGc3i8jjHDyyHKQal3y/G/zgCmtIGPDrdZKFhccQxA3X
H4r5AmZhg/htDaA2hRFxX0/7G/FfqHycNUo+02krDcxEk6Rs8TzkmE9jWSJ6H+YohYd2RkH0iTLi
aJS4w9wLA+eWClLfN6LbBgjcDVzNc/8eqkcxASye59OgjA20tVcLNNUq1Zs/jb3qUNjibTa8+4dZ
1co2n8EG/bE5JTknFE1jDA+tClTDv7+qoLJHrHMxWFY+1wZEyLd2xu00f11dpUv5mblu+gVYaaO8
y5S4pFbt8AxXFzoBwg8AquEO99Gr7nFhdZC7g9kQawW+DuOygpNWjm+JEWLTdZp94am8jQfWzAh8
ApimgkzGVKgNBmr0klYx68Irxj0RuaQy0Cn55CfE6OeqRMiIFIWim/Td1x9N399zjSzMBYU74W+x
PyWdvNnHGpscYMoIUhXxcGDm9o+2YE1q4VftTB83sujCa8bcjXcoz+IzkdYUCzjG9eSWvc80/csz
rQ1TAgiRz/ip6Xo66oh+MKZSpUJum3ULWGtwcE5Td34RReaA5npojWS5ESnoHPVUCkv9vcUu3tGX
uuOq4H9YWMUDZsmKlvsq5TdNThsJueSocAIcWKlc0T0yQLhVkZ8FE1y8fiVHZcaEu5XH4CQuVeao
j/0nvuAqObdUOwV1kq4p/ZTrZ9NmESNhBgIMBZe4/g6BKfYi5+Hzcytlq3V0ymXH43OZR3QL7c/M
g+r7667JjJ1fhdSGk3PsARAOlogrcH2TywJWp98zlWH8SbKZAditdBIMvTIFpgSJX7IpwV2GJM1Z
KPc8lV1M1wcpJE4PafGxu+SIgWJPoctZj6w+kfsNrsGSePeaiItjnbvqvLfkBclTIpyVFdJ5OvHa
MToECwRW1XKUWizNIEuudv9Qk3wbDTPq5pJPSA8Cd1ACStOiywW0ESBFLmHrxSxu+OX308/QG8Z/
WIqllAEpBTjLpr/bAJAlmReuJt4/DCBQD4hmsL1QcBoa5Zm/V9ezes617ovEAA7EVkR6zSjaxkHN
jy1DYhFOv4/vMcwY+05zJCK5ddW3TuOrs18b998O3LqemkKwYb2lvfjiufLUo2Qsv/oACLCfSCOP
7J92ty5J7vMaeAU/Y4l3wJgqP6fri1ub5IQ44t3geNY0/VAinB8dTTmYKRGyX4FYbb/Cp6twzFzi
Bkt1dnYzYkuT4G9e34/XX/7AleUiB+z+n8OUdcvIg93Iw8LUO/cpiEFhWSyDDtjB5tGTJXz93cXM
x633EaAfVNGITvUVoVENNATg+lwclFoFoBQ6ZapwzSj+VTAcsXcQiaU3OeKsz0Rj8RM9n/7DrrLF
jDTASQLvQw8nzRs5hO61T8/yY1TOhUw7+EluJ8Ns9MKwurUsgVx84DEFENG9+vSx2yGFj3SA/7nh
s3xmp2jpeG1jTi9w/o7TIGwvcSbbKdKruEBr2TqtQ0Ti+o+Y/s6qziFT5kVIkwAXtkfIOwBKFq8m
Xg7yACPqWDFuD02nY1pXkEs8Nj1RGLg2tNZA6m7k97ji7/24gZpa81hvey5F9effmAI7JsJCHb7C
ApkVrUwFZ1mbDbg9eqRBQRAG4NTprtZ7q2BBco39CRXVZpjrT6UWdfFVyaQex6YoEbaRLKXALSfS
kJOv9a1SZNRfzeJySUIpSckDUJZs9vDb2PhXIcugVjFY7gdJa0P0b1rYMZKyLWJfo3Q4fAHyGLCU
fQm7uuoTdAaW9iDGAe8502zCh3cPbwyEgr/1NivCnhl631HIjiXkboWmmXokTJrf6tJBBpQJQrkQ
INzg2hofV51RyKxfYfdk9nGGD7LwUKNxeiG1mwFEBex/60qpLE+n7jA6cQt3JI+jK1aMJo7stidu
+gETL8JL/wIWZWf/KPXQHn3+CABKKx4lccfyAebaDo9+MzlI6eBjmhf0GX5pfCdg2takXDeEOc2U
kfEbJsIt0nbPcaxKns60h1FY5DKWawxnmCxuEc9w6NmNYVqqM9FqWDyAHpm4coMUt2aSrA3hrgbE
7aKnRQ++o+qOFVyZb855aFHE0kPUQYU8/h8FQ9LCRrUdP2NidJM3N5/f43XAxkdgZWQw0J17ye3I
mxCb6x6uImsk/iWkIDjq4prFFxgtfPSBe2MnVaFPXgHlW15n909ZYoK2aYsP54TDM+s2DrHSZWUD
GS/4fZaSf5eSzFpHvtdqtekfcYnX1qCEQ/6O4tNKyD9AblZVoXCz9kUDdvBRSf5hX2v7PvrT+Mwf
WzKrq/9/Qitu84ldzVblqdgMptfybMLU2Skde6BUpZx98XKvlWAamJ6bvvCuFmzr4RSttL0h479X
c15qXKgJ3FqVvab/MhByVNfDUBD158Rc5WZfk0JO+RZpDWJvt+Xd3ThmiYdmo6qI+3hgTWpLKMlj
fn8sZcFFMqv1ru2ckbV3O2HfQ6RN98N846E1S1sKdLPxhR3BjlhJtcuCBJ9KB/LAFnInXOCP9RXd
CgyLpyIHzw99ATTnO4WKIP3WiI/I744dOGJRGt972E+ZPyW3MvVPriCes5tyQW/GFWR/ghsJX8OI
pK8n8PqprHZj2bPPRu1BjZepLZu/QylSWiA0B1Eo4C/fvSP1Ts1R8zhDugMEpi/kvRdJx8xpfnu+
wGIyMO2bP5L0KhnaCB8n1WWFJDFhbooqFPq5/qbhxMf/FDLO+X07Fu8DNNGhaNdq+Qu+x9T5aJk0
h9tj/3C1ORE0mLnibJ+gEzu76eKBSHhS9Qgv+oGkZpvGK+/TRiqpanoWVDzDntmfWEYOaIGzAlUe
IL+nIMl4Inueq6W52pFG/xUbR9ipePEpB/6uNnrHrpUxWbcZJNMbQQn7tWmSHbIZJrwPJjmBgYQI
O1SPEtLWpkW3rf296Dhrd8Ek8KnnH1LTah/fNsKw2Dse7d3SytXblw9vNiYd6xCh7T+yvaeQCJaO
dSl7bsvdSVrXLQS9oL3bss78Lw4LgFYI7rXfh3IQf3pZpEmKBYcLlUA+KM3qhXj2SrlJee/wE4S8
PoScQdJKsMypo8mNEHhtOvjjxAbi2YfdyHneHqobqHMwz9l2vFDCIFAyFKdoonPoJVWQtS8iruNd
1ITS2Y/5BMIhuOfwsmNU/qwcIElQG6qLacGvn06s+8+odX0DpTIKt7TwcTNE6P6t8oNSkLBC7Otf
4CY0Mj6/WTMvfNCjlKtMFCltwnT/ycN/jhfl67DdOkcnixg0VWgVZax0kB0vk9B6vDXo2Pu1VjBk
JzvSaWAOsdmqOo1N9DMtD5s0d9nfApMnV3Jc/tHtlCJgiFGSZj51cdpyo/kJEj6ulR7Ai0YV/t7x
XYMX60lKbxfS6rxyrDyc3pM2I2iedmeifyB3PS8zYjLQEyAfvzOH2ktVwM6cm1iF3fLqeCjYjfJl
Y2pi7mMr1fTEgaOk46xaPe9Px/uRA2fTwAFkHMy6pRzd6sFqU8QD7sws1V4t4qXdOfBGBf+J8jhU
CH7aThAnUsDJx4L9coT50XahVowWwbgtaA5z6ya2Ye8JurBeSHuAs4zjYb76uODcHfjBKxq5l1xk
QZyps0NiQ426WM2Ux7zkd69dy+ZqqWfsn+p8Vja9UyxU1SYjpJQ72pTImEi1gw2beZ5TBKc0rbPx
hk8rS2dDxNLv+y1uINP+05UinYBPhgnEkQAKhxZdSGpLUdlMrBwcBt9BjS4j4ItOrdxwHi5LIzIL
9wmKe5LtaK3fvQuvHq2z2LfM/Eo8XIYH1+yaK7xauf/QIn2DmRVhjkcZ7NP2Njeu4VQyknVIRVRG
A8QI2SHyDzrM6OXqcrPwHoAqgEHp/Z4p0hqJ04FYGdLYjkgr+uT4YR7PMcL7gp9dMEXAK4afZlts
kaTIqwHUH69qMP72nHaX1U3KTkDtqGzIXGboq0hKa4c3cKBD86gx+TNTmL+HHv3N5xwR2OtemlD4
a6pS/o5E1Pvk2MShx9g456k4CwQuoHEuNBmSbFE1p9LrI6aprJ7dV3ZIg1fxoaV2Svm4IrcH6OkO
qezw4nbP4wN49yri4Kjgho32Fnx3yRsr9VbLLFxuW14WKq3iFSwNofhMMVATzD+XViFHKjExbZrL
nzhUsqMu83mpPr69+5wb+omfgjC7nwqpef2aTxVbzkrvcGXlKNeDK0jte4+/6lVeyP4tDBBPgnom
/bc+4NVrbuEHfiLolBvr/BHtaEH1kwUqGhTvOOSTqI/M50sg+D5+YLL0AJDdKjIckYuSYf3kjwQk
rjIpPfLJJ0CvTys6vvAuALlvx1LjrvRzy+bi8zaYi5NOSUOgr1pG5ASq+oomnbIIc/np6+irMjmO
BaUCK2+rpuSUklPI1u5H4hGuvpwS3o4ZsfI3qm/YZPu0pMzinDXz2UaZw8x5qtb6hFbmCIBEAqHc
/MtPunXH/jRcCYN8yFY7+Pbt3iuomInwRyV48LoaFWSOzPzDbMO7SOnmGKFm5ocgp70g/deDX2Dk
RdcyYt20TepnQ0LFTWRAIdB93EwV1uIrP+XKw1uBJtOeCx885pLjNZVnd8yG9i/l5hBQln9EMf/V
1UiWYggZhLp64Lir0f2DW4nxoynM+uYw1JyuonUb6w8SypS135Umtdxeenq+86jr8okxVQrXNW7H
FTBLgl5Lahu1CMTv/54Tg51IeYE0BNnwuT+aK91MNl//NUOOfFKJ5Vr2A9bKkFlMK26Zzj0rbyYb
g9CgLpwwLtBxIFsfxpUJTfGm+71E4qqAW0Q853G7ztHz9Jb3I3Yi4U5Hjbb7IU4R1cA/HmhyZ+r1
ERjm3gyY9aq7/3pgTr3CzDHW4KF5+F+o5/xkzGGSgIYUODNEkByMWLAmcTyq1apC0K6mSIBi/ou3
T9TMyoXsy9WK7YmpSjNyn5tEs7hrxPKqvSbMIZHND7svthnmzufO9e101IVw77fijIf/nPYYOsI5
j1ho3Sb8rItgyBlsLpkrxc9/7GfhpyFa2TUl+mrQOH6TNG+l0n8NbyLaaFbAiWt273+6zzfgJBuT
h/Bolf9hsaDxohRfpnvMKKQRbj6Nzl/uddKCokA+G8DMVHjWo/DA+MfkBnQHJCuKOaCpJCw3FwkI
VgDsJGGG2/PRQLmcQcwoD/jpN36AXlT7jDPejosOAXu8uiWZrMx7g2QlmPLD1hKPCeArSrkkkEth
XnmCGlZp601/9deMQey2AQ6vkoa5InJS+W5Z1T2VBL3ko/ocmvqx+9n2X8V8CC/uvyMHlmv0QMmH
Lsz4D8xxFoN3MJtUxnflQwAlRyOTHuf483U8pM5w3hyH125SaM4EooxtWtuWPiKYovCOQZBgv8YN
y4M1VvLKFJfiQE6z5WybM+3SS7NiJbHQyhW0NzTTcfuyPslc6wl5sxTbR7CRBIZN3GAC5mS7Lz0i
mT0CbRqBEGsoc20mBd6QFB9jYkMxPqzD/J0Pcxn7xp/XYQLAmBrFelGnHATMMNniVa9kQ4yJ3R+m
dbPcgt0wm2Qh5dQCpsXxLWDeeqJsuvV8rBT9ZEH/bRUHyEpU5vskLTgkj9qqAvmkBsbkbMLvYpVD
aLDThCefyjrw361jLaV5FLZvbjs1Yy9woybRTrlil+7pdvo9iGZ5gyBujzH/9F4a369XmOLh2lE/
vjFgtERhbtTNHP51Cpk4KvsxI+G9Nj8Mijmal0mYs+faotVhqXqLQl2ieXMdLT/Qpq9HTqwRvBsy
GCrF8eE4SSjuDV/C9lGNEp2DTgV5Yi8UXoPOqHfQbpy0SHsxTbV5suiik0Xqkrj5nkMrKpAYa0hh
DBxvlSTXEydHDLZwkufILM1y+0d4Ph4NgZSo00/XKANa3yzEJEQxZcBLUmtaVisxqGt6NZl7/McY
xJuRiJg87jjpifuiYxYhtVN4WP0dqej0uekd9cIwmSgpHu+TjeWtrNNpkEPjYuPQ9Exa2VEZoke7
a0DugsBWb6ClX7j7Q/rqmlmgcJuPWb0Ov41hCemCu4SxVdpvRCHqAMUi1V0hkm//ZgbDy15WLkxg
YlqpEkObteZ2JxfdCJjg4tEQLmFA0ES+E31mAgycEkCn846q/CshGeC6L8KtZwEq1H6WvbYMM3E/
Rqv4AJjk6ob9ujVnyLj2JZ2InY555btEwVevHBSLR4BpmLkan7AEktpvW+Thqs+GPoazadcFPjy2
LWfM+3nSg4bTTRIVLE9s7+jsea/JLjQOImdVa51HCoOl4DRjDQueide7QzNVuqf9AXz9YMcyJ/4d
xvQpp+J9j2VCfLBpF9GiNX9wbi9SQgKYBNdGvCkY+HxgbAhgqLiy9xcZtM/qUnlzMcKPK8SHSJo3
8VpOumL0HzuVk+C9XWGwOxRWLOE2NH4COHEzUZdhEk6YxdosjusZBKC80Ar00LI6KP6zueVyUmWH
S4XbyLqz7kEnPvOrrxoBU789EqzjR1gwq+C5B/EJpf2mcbX94MIxt/+65mBhsKieXHdBhUuK93ER
zipRcj5kSvZVvsxAyPe5rDXfgpAZgooudOfiN3fzWE9gvL3u2O1x4kbheh6qy+KA/XDSXK6yzrbL
QyOB+m7C8TyvNd5m9wCKlM90LsxGC02wR6isvl+le/e4uyRInk40jcm27FKVsIh8JC5AOVAzH//w
OlyoCM2DbPsJREtflarm783vPmca5ElYkD5xmovFFrzCHUoyeECTrGbagKeZwG1tNEYloKijyxKA
NFwDrl+GbQ2ckOYWRdYLipEGZxL8N1VHe/TF2fDeo7uzLoO0CxPpxqyaD6dk192XGNrjqV6vmrc9
QP7/ZdqlyCh7YquG//B3a2oTBB5Uvsr8r3S/MD1hW49KXsXxlXpMI0MYimwKDjcPrmJOkQWKDh5f
pIsQAmQphH1Kq5249qYC1a4bJJQgPbShTu/KEYU6NUhc1Ey48jILyWq+fPak0gTYSl4Pj5USySMC
cbXV3xNu4/oZHUch3LnuI622/b6Ej+pyVGrqT0/JxTGK4IDH+CdKkefslYY2xiBd4pFle91KhZwK
fIBUejhQbNTdPy3rQUGgw3QSuS1AxMLkwg6sWEAU/sBIIngPcyNOczrNJ6r8SaMgzdTkjl1AOSHp
JuqYqtJ1SYnkcXMRdyoPdrXgqQS5Cjr104JKGXDNN1rXPofTD0df9c8Utfjubo1idlGSQqzaNL/H
WGGCEG3eDdjgC66/IQgRjRnX+QTcT4TKNmh0ZD4rQ/Q2KfXGXUCP2V4MGeXxT4hnIfivQXJEgo9D
vPoWed35oNSbgeEqPjBrIwTY2ch5yVrSTKLatwt4WZhgx8T2VfZ8JAQqBq9P9ASzdj6kyFDAbRwa
MfyAojHqtDzza5ch14O0pdWtSeqF0vMP9vpbsIDlgTQ+2Plw+04JtSLUeujXKn9fbJl+hc/3xGaW
x7lShi1H6CJEPT48K2GodnbAmpJTo4i4qlpGuSXueJGpfirBTnPNllNOyJOaCQP/Y8UoJRbj5XXq
eC8u626ZzpU09GCKFr+ouaSWS65Yb/t35xwz+WipD1qs6TExq3JfeewUX5bwntnX95QU8d1ivMSv
c94w/7xbfrIgvVX/aOenvoMQlkLcDfC/HVJeU7TNvoizlSgmIZPQe/FFpv8TSXLG/CgRwoBt8bLR
tzaq3UgY2jxsBRTDHVqKYU7s0nVYdyV7rCEXSZcRODUt3aoK29/9OOyXBkanU4ovIdg7fircE3XK
DbzWpbIwx56ENd0pD5jHbJJMQ6ehwAkgm/UhuyW/lmzU2lcXX/8qu0K99+YWmf2bRoTvYG101vmn
1tUP+Fdj1WS0Non0KWkppIO1lXyDiBp70uEDNCtLtl5PBuXO5huSzTpJo1EbaE47uIrPPU9TmbMy
g6ZpDh+debEofQJOOq4eYLlrCi7JiI1xTkxMWCa7nhbd+7bnxztiuijwzpCrwR25jJTcbMevb3aH
Dnb54Ey8tposwlfz4lnRI/3q7Tw6xk8Og49hUUHBH+dFGEFKT53dLN2j0arv/W6lk6OC5AVsEat8
/m/VPlQU0YZtVrLGNQsvE9U74hWUnVk1h72XqtATcP4vP0z46ES8GGGLVDrQ/YaugyCQwankF9D+
gCVVYqxPz+swGQg8aKY6bzWSXUXWPhOxg+9GM9IznCCnXgOD8c6u/RLaUpLrp1Is5zq9jSumpmz2
K7LmKf+ALVqOwuCj7Vm92q6rsqC/bsxVdth3+0gIrNjLkBcFfzLl7fufIjUvhXkzYwVnIhr4eefc
E0CwF32BbT6iVXzCmuxqWHg557f26P6pTnXV6PkJYgtgT1oLeEyMbr6Y/Vu6S2YijlZEcVjMvk44
AYRqu+rj9+HU0cyzZiiSyWTjfvlOScjh5vs4CS8O/D40kyuscnAWBe4RIwojkcUQS8LeHWq4yDew
si3+HyvHI/N40BAbZqohjQy+flUkmKj4J92uadPhF4Ka38NQgEXJyCksV7HpkQT7gxQFyxlbOtY5
TjsXpdxvvWDMAPj5ZOqooGy+caTKg3ZexkdJZhZhflU8nOFIma3f0zo8ngjxg2qPZ/1SvxKI7R2c
81zuT4QTLOqqLdrfT0bOg36gSCcj1xKZ/DjZjDZdq0vp0a+8+A4rrqcozo5le2svS2/F0HXDIr56
cjopwbuYSxQc99t5XFwY9GMl79cR7BFFyZhmG/pksS+/dnhbmXURE4oHVz11dRT1S2Yy8pma9lk0
loRD26KZPYRb7BrrLaQkFLrjR4J9ersjCZYdaBkL6B2DBf1L9OX0PnIyWgYGTsfhzmxqIEWvkmXa
I0f0nuJUz71Cq/2L0SmLqIyORxpg/ZYuZNSzP9uFTAO4rLU/dCReVZhzBbYhZ//UtVOVZZbVdNMg
ZeYqUKG6EAwUqnJXJp6il3uZ04YYNBo++g3R/JlWavHhFC0hDoMBfaHskw98UcSZIpWCkRFW9VY2
QPU1cpiBnNZNoLCM4tGDU7jvqLOzxl49M8vlRSIaZFqfB7AygZ0S5blWcHlgoohUqPMRb+n4HyXS
t5Q+scQIGQojE8MPe5fE/bzIWwD7eCdiU/RzL3yAq+3w+p2elOdZiyQY2/KDUzF8vStxFf/6ZGab
PnhdU+24ZzX526I67tr++rU+VI1cidwiD2QUQ7+5BMr6WRFVavTmmdax5CCRuua7/y6j1npymEiP
xs7qNh3zgwqm11qjqT31v6Qr5fVRCNLtWhsmKcyFNgr1mWRp2SKW2RwDGA2S1ONNXnPb3B1NVgJF
0IwgcYbTpMIO1LR073vFO9x661uTj+qxJuP9U78hTpf/fIvCpgz1SjEKsCe2D/Vb5wUkVi3E8tSN
kOyr/iIsGTDT4RPCtGNuRJtQ3dVssO1c/eGPLitoIj/MUdHQUukTknTnP+W1DWjCa7T3bOl6sjDN
tWlR1GT3ABJJjdhESBCryJHk8+cpo/RjL5J479sEPSZaA/gEvoAkhL6ai+5Ke0VXRUsWTLyNRacT
7YSNRL0aF5baeG14l5eoyBKZ/T+4N+07V8lnTlu+MEbBxL+Feia4+WOlUjtRfkZPDaoWAlFoTI0A
zuHhBjNuopCBxMz9sznAEMNXL5wR28ymq6hhm+XwQk1mVBdoBJ4LcRyyl+Oox6zR37SLG1JMD/iJ
i357iNe+1x8WozEFlBMoj65iP2nOsRNVQSeIGavgMh6ehyNCzfYDFa3QlEN9juQERx5rUq5W1ZAv
Dxl1Rs1FNIBRXdoNZRiOLnluGVa+jqgr/F0ORGlmHWJ44VNqImXV7bRRig+wtRbKFU3HUt6GAqWd
fKNCJC2UOURSotIANv22qFFbA4vvZsfpgW9vp3FhS87vrPqVN4YA1KST+76FPgSvST+dGdSTf1ay
eO7NtMbQVRz1F9JN5BMxUH2QU4cZRR7q5MWnZ4zkT0Jhx9fugptesGgxL/N6Ww3H8Oe2fFAREoqP
MRNTeeC4aidH54ZzLWu8jIdomzgHRt8tP/wqkQlNDQ5fvE+koEp9W/hOQ3zIMeCKLyGI17koUTiP
hmJJmEYK6MLERGRe6hvrwJTrD/5HFrbH+PoXUrpEa6SQQAMkT6aVBo5cp8BwC6LWklhZi/vaR2tZ
MOTLAiXh/PoEu5Wl3FWAKOKdlYzCDhKN72IMhwtCcr7kP7G72KbGwEWhdNiVenQsksDf0cbxiHSm
U6yalzm5MTURJivb9tLRcYi3gMIF2TR1/nDoHCAHjCFNtEe2CKYz5SS5O1VUIw3O5lIpVVCHAHiR
FykeQJ/R0g63PgCiAU8HeetQudzuHz83tkeVXUNOOv8T6HhQy5RnJbDKi8STsgGf2aZ+vegXRaZY
IOG7Rmsw4fJ/oHncJ5b+lhMHgpICGjdC2bAUuv/RdtrsX/+k8jCJsAZNEOS0CUs1BJCEkk8fnOX4
5JrPyzXb6Zp3eDEsN+2nqB4VNc7qCE5WAITDe3NkmXJPQlGP8KoZcACQZzNUlaHxxPO5GMBfIy6d
C854Stn62mOUR95I8uaq0HUKezNQP6dTIpQlgP2D6PvR+KHddBcySfzRRMNxH8T4B8r3pJixr+ZC
OEiyeLaMyq4x2jxX5+MFwtObSIEjTHXGs4AVRxp8Q/fcrLTSpRpqd4s6b0+E3RgblWf+qkPTwUtj
THO0U3jBEMcoEjKg/J5Twkg7CaD//tUxe4fB38NVYS/q0LUC/Mi2OX2pqINRwn2q8BRBUHrp9Oey
FF+3ZQkxt21pVpYPOAROA0iEVHrC7CWVsQ8lyXC4BsHc5PQBSLTr4hlu8nR7YK+W4Kjo4w/AqCq8
BUDmi+qnmndJSVUz6ShptRaki/KmNuHwnJkjtJxN+hcFqaIhXTsXQlETX90N+MBaCZBr7QrQhkQ0
Dqf3NceGW+YdERhaY9RdHvncS150zxdt5foQtftILAp1M4cj1odVFENVf97iuNdfgkZwtV1oUrM+
nYrt4/2fw1gxmSj4W07wjjRaEtNTR+GbzClSWO2TKmgdPRQnW8erPHACb9kYHa8s1yXBtRpPBmJm
iaqj0LwNgRe04Tpf1XtE5DWppo7YM12C/0ZsbOihHFzYbG+VKRHY0A28lKm5oRTANosTJrFFWN4g
3c+jFBO0yPJPHNfHPaPu/D2gSd+bmxeui9Wmi3ZAHXX/hpaGHlg2C0XfF1kw9/wfR8ZkbGj6pt38
KMLaPBrNgO9+okeOkAGUUfmm08ReLLIMDfdjovB9ZvG2ilL8dSj1MYVMPIqkAF+dDTYJbg66Oa8b
P8+eqBUK/6GIq9xIwnFPDuyBDRkr+xiHzq7sH/6a1bB5qPNnidPGIWiR1T7iWCAvlxTjXngfTRa2
L/LPwV9VrmHgL17M8wkvR9wPB5dbDwvvGLUBGEGmdK0+gIcVGcH7fIpMzs3Kxqql16Idmah0Vs01
Fp6gUB1/Yo2UJWD8oX2nne0Sr19xY0FD8bJtLmQM9CET8IBz4ZjdVfsSNdVgGrAESgH+FvjIYD/s
PVLRMns9DbI+SUABduJgRuGMzb5VJrOWigbJ90Yp2psFRWPZOhHkWYbYLPw2ALPB5fTObTZ/wCII
coLz0I/URfxL7j9btwP1dUi+vbphC908jUoV3UAvVdb1VbFajLr7vhO5MsNCOvfDIkpPSpWBGiii
rJyj/FXz/A6lBUXlVpLroM14EaugDLLb+iOVXCBRNW405jNcZ6vMSYljkz2cbUO+MrWGODPnhLkK
MJ56pT99qeGYfx0cxBA9dy4ujGareClrS/vcwgl04VWDZDwrnHUELeSOjnbRLZNwxLP+BQ7B3JoE
hooVql1DksMD8w0fvRmQKjx6c7Ri9J0PKIBEEfarGroaS7dAW5W+x1uXyhfp5oqSi1CrhTu1VVag
L9jmTwND2jMyTqUafB7Uf/yo0WzuRm2f4Gy3FF1/izKYUfBMbIuJI2W0xnIAhewafjkuZuSLRZ4a
PLINOi7ST3q6qCUfWY6hQHzfDGNa6Jo23fkeru+lCz9DHE+paQisOGS3jMIqXB7mBEvkyfhrG6+L
s+aGG7N20VfQCVQDgC1PpOrPXcdngtQ0JlWZGNKzHhUeYfUH+FOeGSFaxlt/qMW3wXDlm+2ppHSL
MrChajfkYAwA6VDUajUnbVU4NnT6F9eCOJVjpCQ/BURs8wjIpyNk9vmjSObV/QyuCSO4LVHRHZUa
7kmHABsOh1QM3Yrg9GxNzuWAAH1A77KhxqRdM2w3AuDmcogKCPtZIlgDFu5W1BrmNsbs0yfaM/9X
zmYeLFvDQqEJ8pq06hCWcUJ51TErwPYSzQOUukGERLdeWzLbmDmyor40mMKRKVTrZVntvBF4BEvy
mOItC5+zbJcD692QKVx6IUlmf8IT2+Mz1TBG+QPVxe/E67rRtis7tqNT7ulh7o6WKzP8RxJGifPz
OsKHzx0mTekG/4WXzAp34pq781SA/lBTbLMKmThzwhBSpX29HkEhS+EfyHdxNU9BMj9ht9M4R1od
V/426ZqTmrojadIvnJU9SuvclhAqOGU81SbaX780yXnRK9BQhqfjVKoN1jF4nWaD5xVdMdYOujpe
XMOU7kgjAHvv9y1ZpOkO/1v2hqnV2aVMXRljXysSbD7wHTCa1jKbIEZWq7lLrPpD674h6/6JcETB
A0f5JxkWue9HHQAYGfzkgp1Z81u4MOvVlRmhM9u8BhFqjosORP8xxtfkSqDm34wBu7A0tVcEuZXt
yZVXGIhD6TTa5WKXoGwaDo5tZ6oDqYdhe9ctgL5bLNSNMglPPDTKSuMclwZ2c5rfepEHeqOzgxiY
C/wCkrNFuQxb5g9FbeAXFUbbq/eTykRAJluSdEME3TUSQ3qAQuusgM++OarQiO2Dh3/C1OVjAZ6x
7j6SeVhrny3wXRrir8PYgyOThiYE5NrxnkioYq+wAfg3tG5DahLr7tgFPAKwvelSqwUxP/ijol25
8aRQ2OFXwLLQhqQaWAcJCXoz8Rm7TXOPSF3imdYsMCh+rYtIF0naPVxC8LtbRgjDBXbD4k68plO2
aheKGkQKs03jpVsFNlmF1KEyLV2jEkyduVcm59zxN2JPOvo8d4VSwde9vT3McebYBHpkj6PsS05j
WlVxn2UDQeDOJoaT7vl0LPu6qfVCwJ6ab+Zdd3BtCcMASZ295iUIR1lcsvnL+sKiSiOejCgnH/Dv
a/CVu+8Jua+y5d1sBTylQrcLT9Xr/R0BVI8sAArjmwLEU/skMzC9aFR1IKhg8Ya/oR9rT4qG3/qv
zXppDxcw/KYEhdmOgPZHB4jCvzyRMacrOFPRiUN98PyAzb72eMFRNNvLWECj+mUgxXvOLlC0fiUO
XW7vznWRNvEfzZGXBuVdjV+d5DansVeOQNLGaP//rbxwXRo6VR3PDrvC7Q4SqhNcqAVZzcqKP31M
j6C1ParuhwSWWXHzsPjERnQx5frY5txTNvkrmKMxo9NFbXZ9JPA9T8Tnqq4xsv1+VfQLrl8vsyIb
eQm5P76gxt8dxUbHvdsfkWsuYpefFZEQ+PWWpe2qxYyftwXJ9g5Smh6MpfOWuQXiC6g1ACUllqkp
1lE8linJfd9jIOWYnAN6ZRHWU7rxUhRPwJ8bLG2hADsepQhmE854ps05wR4nKtswyfM/UNPgVIra
69ywpveq3juLaxcl3aVwznqMjedFRh7JsGfAcMaNOCp37Z5pB5+vpYgSrYDNEKNWJesyCZdCJa8i
uXB2xe5uWFy7j/58joLMt/UbIrM9Qh1RNlqbgpiK9p4OgofLp6/6dnWUFpkzEbFZKEPQ8eOFki7S
MTaOxvT13TPJX9OJ4BTC48edvhtHmW0uLiHIPn4S2UTiX5SHJTxzm41gAdPQzlXrf95kah02MxIB
h9cKpjinXa+lH6cP3FsYk3BdvGcHczcuqL8mpv0uXzKU7fpKU75AveX9IPGzlhFDpWi1gw+DS2DB
lssdvuum47Exv2Kos/FaKgq+d5HvPfRceOdhNI59CtOXbs/JSxpbgFsmyGRIrvIPh/alditpUgwR
FuZm046azlBJ15svL6K7lETOamczxxOS1+J0eediCKbiRpOfrLUr6IiF1s+leZ5OC0/FPxPzkE7R
mw4dwCBdiFT3o6oqWtzAYOmzQjDbQMlWPnb2gRKp8r/39cTzd3l7EGNxPnoJUuz8DwjM7VKtspTv
3Q+TPeYuD2pyAbb+I7EpXovOdbKAd2kNZwnVuWeOYo0NMm2Gk9PdlP5qoKU4TUFllcwatL43eGYq
6NKpbF3+AfSXNtBUKm54YA4ZYOD2Hsp17UScsWHhuQwkPRc/4w8pj1t3hJQbo53PC15U9HADdTXK
4BW2RvUXzmLMDc7Hp+gDoY2kaLc94yRjALDoxhwelAPLLufqmceqEw4SNyT9BjVhYX+mgGUB3fEn
SZCgls3UNv58hBR3dIfCVH0Kt6cbbT1abiN5DuC2Rn9tfWgVJe/4eudrXHeq08bEtH63xph849MB
Q3O1TBMMzuyxpFljqTxOlyXO2EzC+aIDjrZk1BgQLiccgtMCH8RmLCo3pugTrHxnJf64wKzoFx3E
+IhVyzySfIcinU/bUuTM9s1er3tLuBNPxU299SdQul0uzyC6bMz4VnzUVLuX81YLAIxJTfu1w4dm
ZP1G/iWM6cJ/sZ0TWT0h6F4BqDPHg5oPn2gPsRumoHRDVnoYcXpiCU7e5Wop8H/W3ps/9zp98CBd
sR8oAknD152fxcsobafuCT0+vIK+aXa9D6Msetx2wfnS85rvPBFOuGPp8LObcp5U1+FvpAfoV4z9
5dVlPeyM2ANLjs9o498wo9GxJREEbl5pdQs1za/pt/WaBar9gGIxL66AZKQJyaq2v10GgkMF1W3Q
E7xhf9FnIzn7V/oUhKDvzpltpvKyr1j95R9pyWzSRPF/NnSF0BMnhlEOvAK3GK2v3EshcWBQN8zv
DfuRmoX5DAgOPv/pV7mtZP2dCLlAD/6NJrReS+yfRINEOrUUSeqSFmRuzkzEjOfbn8D7OqqGZIpD
VuGAkT3290nw0PX0Lu/h9T3RmMBLr6yCesNa3MGrpo2D0xpw5lgwQfTyLyRbFAX2sC/WWAN80VcI
ke9hILYp2fGy2x4S5Pn5NZACZvalbsgeHwAdH/sSjyTUBEfkS84wVJ4kIKMy8YjoVO1OCTfUet4P
ldRm6QGSdU36hpaUwWn7zEmZyBaRMMPh/J65BN1AIA+xEfTIdJTavec7LsFbK4yQDF1CIxAxtkjG
dWDahTBEsFo7rWiaBJupxlYBVIUm9HVI0wbFeFLwW15IwYSO1THH/+O09Xg54movRDBMZQ+3pBIK
Hip+9O4uWDfKwy/0hCXu7Om2Qz3EXZFWRlzpQcIXPy+gGKOdAuz+ZUV/A6u6Rktg17e1yEgyRMjt
mA9jOZzd01jDvEJ8LoFnxaMOkLfRUngp/YUVjDc9Rhr7QqGp/DZLBF0+FVC+VeGw947LwaMW6KUn
6xQPocKC/+NQStN60cknC3JYpVqFikQNITrHCAjyXZlpbECYTJ7K5KAnR2U9K2rp8ilI1sSP20YS
6eWlDKlnRxz3fuxKJe+vM97MYOHN0v0MPes/a482HAGWCSzyPHKDVfaBhLP12hb59TwhkFHg6d5y
DTDaGHptWmO6/ho4DxWXLtxZ/4HzlCn+nRhKX0skLldpmWU7Ezwn+6YLcy3TLXYk0UHIPTdUzBt5
wm2DBm8ZrkmDl1U5J95k4icHm6WgJd//rFi+IQG604CsQLFP5yi2lBtmMxLL3y301KLzN7wQnQog
Qtj+gToo7OAKl/rfO132itD2/gjs8F5SfUI/vkseDP/VtXU8QtrOu4jvva6xHw0xMEAYcRhKFo0w
1hn2BbCacZTVwjE+8LE0dyPKD9fRn3gYD7IzFw4El+KmlEZgXLd4RNf0U7HlRSrf1hxtG5OfwfVZ
J4UoP8IVlhZZk4mxBXnCXTpWCrslg++5aU89ZAvwOI4y6c3f6KKQKaFyrG81pyerI4IDAxZvfbtc
gOf5JvIJ0pMAue6f30wi0MGrmCfgjz6h2D9xolv5tnBdjEhWAkiVUkRCZtlKvYNtzx1ZQpEy3iX6
u+qwqtfx3H4CLENdwDhfWIo8P8lyq92gWN29wkPSupKdgOU8FctwrLZkL3+jnNE0qGSf9pO5eCNC
Lzs0mNm1eQxumBRC066GF8wKt/Mp+lsaltkAUr+jJw7A9A6cUeI/+sUQY+lgXNCnVsbvVqdTAaqA
uDvEBvXT+83lT7ZWn6MkEQs4TPOzSLqrPxkJ4OUAbpp8ncHJNCbt+yenUSrQpAnhecuBlH/uuyPO
MITvv3CO27ovHx6TgueQ+sa0eQouQsxa5E9+EXPIx4i85ZMkSyZ5yZdpbWfBTajiv2qSDktd1P80
0E40VHshKXXbxSwNPG2tRzB2u3MJ16Acrznv3jyFgBgbRPV9n12VWfbOu8/At6j4byeOeOtxDVVG
I78tTnYpXE1193WAc5vsTGrosJrsjrwSmy9RG2kGsM9RJGEbp2x0jON6/rYXn3QI6qAVFuDgUhYq
IAmtlXGw+M4w0f5wnRunPTuqZOIpKEfuwIBc13vTPjtjvimW+SkfkxBr4o67QziTsdZmJLB+lMxd
0PUIihTeP2q2AVhTsIA948pg5aOS6pgcojtbHok1jN/9oL8SREPu/yl9WCkXVtZh1pPK+BSyczhL
6awD1LEc/ladXhuHFeZiAGh5sMg3ro3/sGasDgKkmdbWFQqBPRYZ6PgzhZPY7XDJ4dMjorqjMxuC
EVSfoX20vBSZOkd6/T0g1TPmI1aa3vTF9VZCJ40rlNwZ5LbKZUAVEMFS6jCXr32CtwRC2druiGeV
6rUNQOmFYAa0gJSg+Pnq8yNnP7m9VkWvuxa9jYZ4e3RKwi/uzy64WGJa8Kf1FodSpII4ig1YT3pY
mJw9bkGzFUfwbTLQ34TRM6Ze9KWb/X+oR+zNYeWOvklst28uaXxj7usao4+y9F/IKDvz9JUA98k6
me+xSnUQhWqfAvtcOFof41XZ8FqAoivN6X09v6r8eeSuJLnaGuOPRW6dxe84lfzqEDjqYLzJOADn
7WIHLQoWKbR75Poi5hhtiajbIy5gCiETCYzHZqtA/+2wKQZbDGoechxOfVGPxzcdiBO8ywgytbfV
9QuNTIDLadZaxF1PueJcfvpXqUm29pecS7jTMi/P63ZpUTje7lFyLuF+JKg+SWiX3/nvKiEJoQbl
YlOFoNcZGc6GGd/Igu1+96/ajpsgyotPzOGTlXpy5w4XeJrmwb6KDpr0J3MI/349Fo/mfAvPP+Zx
fKy19IAFAPqRI52xPoJsPH8KagyRoAnu6pQEAhnoHiBgZp609jEWrjm5N8fA9aeqFiBQZ1paSbGF
CpCYVsvAeonqFgF2bIaAGUgBffcNXYe3T7Vg97zVsHDQlLqoBTGEM7xjIXl/29HBNwkJ9jV7C1e1
PT8+D3OUEZHUogtMakSutNKVawE24hJN3eEaqKKZ0jnTyw0wdJvrOG6viz76YqzbTBpWXqzi6KB8
97v7u2j8lVvtK7DWBwyv1dslv2lKmYv+ChMNwBG2XBtpHl2PND8J+takRB5i55oROZsB/nZXccQh
cY4pKiQ7+SKKIZanKPzUpW+UoACkcPQcwvxTp6H+OsOoD3WoBg0mauxXiL2FCBUpPlmunPtE+h39
f7HUTVrpx4TXhsK5PRRouZjwHK4liiPEztaGnXDsgxplOXem02e2wg3iPAjXXogDxu76HC54nHdX
kI1hjAT5bZCV15v/gyPsHUbDl07LmjkiivTw+roUY3WwyuKM7yMb/Cdqb1BP2UfGM3AMiTQVt+2d
oFUKIbQY5DjSYjJT7SWi7vtl1SlYg4vaY1cJafavPZrMlGyr4YnbqZH7dNREEhgBYs7C0cUi3NXV
4fGIrHlPz88nA74kpxrLIHIBblzkf75n4Q3btpbqON5icthjcIqPDmLw4Y+ZDWr0vRIx4oocOJBQ
7yBA9kcOoyrO/Wnz45DN0Q1DUbbwVnHxQmOY3TDrWPjeRx25kyTLuLRpykHpFWjy/B+N4su7cCRB
1RbO85Ns1Exqx07ixXxdID0HVZW2aNPrhvQ3xCSMrrjwDBFckn/umxBWr+BEeDj90X6LTz5shxsl
GWZW12FVUxBYoIgZwY83oW0pIPGcoH8gRooBJeh0ekIVp02jHu7c2kCEcp1X2sbYUW/kWabqVMDy
9k8DFvCBbdlVvLscqrsZWllUsTKOf1pRqQSL4p3XtEC5eJiI9bPdYvN7iW+rcouSi/8yveSJm4fL
bavOwB+VksivXTKXoEkwRC7+EsnjkEoKPo/sL6hD7UESQoMHvudnQUO43Zgr7UnowYhWyU0PB3wf
5Us89zpP1oyg7b782wY5//6pdNOzRkr+ghSKh4/X3DIGUuiAHwJ2INXvEbkf9N57lHRP01a5rbGQ
c44/zXg6Pgm+q5o5aXxb/8L2sErfSKslYKISBlB+4Qy/D2Gfmxh5LsiO9dr6UKQ+OdCB6ijJB3yD
Qzy135cKVqSIAOXNPIjt2UKdVwNG3f6rguYcGkguxXOfPrO8xwr7FINv8MOgXeEPluHNqyOkwJg+
YRGkZiIXoUSV10PSvowliP2DMrvY7R6pFa5nIjhey25QpcgJgJBe1XF2PXyX0kEo/LUwRmWt1E+3
qVd7ZBpKEEiOFOa4V9Vd2rBMq7l2ujaaJooZfEkcZoQJFqa0t7z9jaTu4GSTFBqwdKwWJhshCYku
MD6nDd0eGzQ0EaEYNr6Mx8rACA28kq+DyrzH+gz3uKhDHzZUk8bgLViiz71p6/xOVoW6ULFTMM/j
ysrcyqxEXhjfmcMIen/Qydaqsee2sXC0hMkIRAz++hw28eVo0U2+wwxzRqVfhbaJ9Kv/6tvYmv59
yQAo71pRyCHIVdAPB7XZ/1RMxm9DSA9rA/c3D6Lcd6MNlWkCH7cZ3mRtpJ8Xc6JnDL9THkv5cU5q
RRU0vTDKsgostDMPWFlEaLOHVSrpF7/wfqNh0G+cHiRIpn7y202C/evWlgX+55ApuVAlNBDMsGis
uvIie9pH4jVXRmH95IF+vPXnfQI+Oz5b+cHMx3lQXySwdjNkxgNCQj8aF9AlY+0c3QVCvXGXv1oD
3xDJxvBM5haXsqF95SzpEiR9rIblcGHfkspOQm/mpF363Aq0ZIHA5efpSjQKmQKib58HwADC3l2i
QY4165V7B/eLVQhjzoIYndYHncEowivgDacp1+wSm8AOA4g40GXF+KqMnrb3MWqUSg/X3LpOX2k0
GgTiR/ZRsKAtUtkzeP3S+cSaBdOfqAtyVM7Uu6lwBDGPQQPNjcO6kyG0e351HumjQhe9iMICsnJ3
dLTYnNlebXL8orSCRPfHWw+Abh8SuLBYA2MsiJzu8o/CwCNwae0+tCl9zFVB062MmPS16Htn5JPo
gdRToqwuu42R7AqrjjkF2t8ATUNsNYW0FPmmcV38u1DUuj13EuNmKBmDbaqgvRE18eM8mJr2oIgz
Klk0pCaYSEdJs2XlVztrpz7XqluBuBuCd+fVfEaCs6AH9GyHFp6iN9davGv1vQxx94CgIsF2pl8r
i/f0G4GRmC2W92oDjPNGorXsPksWUiffuCACZS5mNjyRmOnoPPM4gQ2UchV0RXc/dY/46R4IRiXm
5eKX0PXni36sEaBy7lvwJ0hBGG2/W815JWIyarFwhZgooVeadebJ4nZ60JF3JyIhRfvxAiQ0YHO5
LTlW/YJK+Jt295sjWR27jYnXF3HXsczBWTwqEyfV8ru5ea6ACXm+UeKDfbEbF4CoZWVdtea8FfNW
9Q/TNhScL9N//BkGPRNsAl7R9BDr9xjYpY7Gr158jjTEFRRGxFR1xdAnaEywBfkak9ML0p/+SkB8
5QiIf6vKNjYzQ/1mqreb8MxxrPZdO42cgYsd74JJAxv/hS6212erqyrNohUE1mg1L6QVEUEM1JyO
WxPAM88rNtGnJhYwSEI23vXR71E3KHKkudAnHRyzRJ8uzhFEGyUKBY58Bktf8FIiIZw4qMkB5uGx
WHM7/JpARD4POBiuwuLS4GumgzFyn+UdlNzSoeXp8jH2vPicXtbgT7d7voo3ZsQ/7KNCp4lf+6Pf
JYrz+vFIsavcEVNx2iV6b6Hkpn+hnGCGDTRgTXerRHbOOS1pEO56u1lbBFOFUgAnIInNAaoBqXP1
uH5L3Iasmuei/KVZ7Ssv+8hxRtr+cZ+ym/k7UvewEWcaSpJsQMDgLZaOWjyizO/Q/Gi1rQmqk/bU
DCIQ8+a0cqbLyABb1v/IEiacw2C9GCwBGZ6bbbmxXxWvQ4S/DBphcpnfZOndC3MI3IMrraBiU/Bi
lf9weU/TUrAA3c0p9kv3qXy15klwkAaeTUGBOTVBgeEdKuPV/gGMIHmOJiXw7y74BekW0nWooPzZ
koF6zJ4LiGXbA0lGLe9zfYMDERU0yBeJhjz6SM+ZfQNcHYfzQvbF3rQz3VZNfflsxQtii4Tneh1z
2pNZ9nUx9PJ8CPyOoO3p8OdcVhV+YmI/90HdoFpRlAwfi86KVOb5lu4CcMAe7Js/lSUDUFNY64GL
ZMkqIEkUs9zsdTPEqtEJllWzcxMZ/xSvp/eAtwEKWesb7O5+IH1mS0lZzGm+LRibS9QKrNq+LvoI
Av5kZsaSMWrGzGUna6Y5F2V7Zu/kEX81g9xli4pTHcgPQOCP0ZxQej2oMvQuuT0yjbKKeGCVvuPo
tzZnIdbh2dd0Zw5Pp2bJfKWzbwggMtajov4qIJkiK+hAk1DqUIEkVPBJrP1qNwhvEasrnpcLBKUT
Z0PILPrdlGdcW/Vy2qKafTXLuquQ5RaGVybDysaMsAmG4BKFod5sYmdlG9ga/DjVxsYW6O/WCHu1
E/aeEtrXbpUGc0srIa2MvuXAU1WyY5iG7x1vHYCm6lUJgWilEbgJV7uI1MkVJL0xYd3D91mHP7gK
1X7RlAIm1of5xmDwZqxZ4wdnjuP8BynUPGT/2OhnkxusOLPBQXnLrVeTt7T5HgfwVXLAj5LBP9GV
VhTS3j8auiB2pUcJ7yT/EciW39siu1jCLwq7eruLRgiKL4M8IaEgr0qJGQ2DsHdr1tX8JSKxxRov
GAgG8bFYg23af6sdlK046806GUUt9Zb6Ogws3dH+ZzX56nvfSGXA6MjIIvRiTVrlrNFbUVVTYD1q
BdzBueKERWNn/lfKJSxGPFCginI/w18l+yyVbsVxWWeFQuKHR69N0yw1ZCBeYST4Ltaqvb6YzP+k
H2sQ6KuyLkxa1aAoTRFivCqvVMUP0lRqn/BDbLGuStbexWeFzbuDMEWqAEe8aMIm68pHQNvqFD5+
awWpCkQE4o2UKiu6BWAPHb1YFXP7sKFFOZtk3G41hJBaKrE8Z1gt8cFD9aYX0WoP0qbpggn2s9ty
Ks9+3RWJtinoiuNoJfJbGuOVMyy753vpa5fmLC8Emc4iztKmhB6urqD2MaZNb5khUS82jsvaB0NN
X1aj864veAvdyP16PTC4tWZMlcNrPUBkSEH80mGLAg2jVyS35dVOjljk8bj+wdtFdpB3QwXSc1oI
wjt+cj3kZdJ21d7r530yP4zHewG4dprrS2Bp2qql8RX7b0zWA33YMRpOXpeNUZK1OD0zqHopjAgA
j0kHvPXZr/VQgcIAZbUzNtaneP3YSAYwZ9vrp5Il+Tmi/XWmWK4fCxVXBktniRdzz31KZDnYUwbT
JqsokRLyDPvtpQJOrdvHej+0yOuAA6Pdsp0JhLZeU1Sn0aQL+66+N6m/e5/gOiAaqt/S4DeH2y2z
s1HJq+9tFDOptBM2Mhrq6f/I1cekxDX4dbiF92J26bKtAMYdw0XBtCQ1sjrwcFWsy+Szq/Rw3AIN
KK+VYdKYlqY/l+Qillrpdu42NBe413TA15zqGMczZ+nhMJdfoFhlMw+mNyVD50pb4sHnD1Rs6eYt
+/KnWSrfwhIQ0bIemNlMH5GBhtVYyOKCNjb54Ss8YAnV69N9nc7iVo1D6KVGd3PQ+4KDjqNdoNpG
WHUlh63dt8kebaHy/MWsqKqhVk+Avf5nd5ckDtwb5kx5eO+oJYTm8dsJy3t2nI4hiXWQfEnzvJrj
AJ8/kCRsGwj/u+aaHfhIVm2n8D9uAWOfdUnjyb0uJUxRPM2qQYotOoH/ObxGPjb0uUvom35cGYnT
RrXZhIJ3abvgAJAFG9/8EjrtzhegbPRWllIab+Cg06ICyHjJ+ntMcCCrAaOv+1Kb7yjPIfrAFyuN
nl99+mr/QAMezFflZrOMrpmrJI2w3NRCn4RKdC5cHbF5Um7Prhk/OexGtdf5oNG4nqmDr688W0B1
kEF6gl6xSCpTIW/SZaDKqUCN1pACVyG/4oJaxWSEFHMyBcO2G8Id+PrZAzizvfzPM5qkwWNKHkoa
fuZdwJBr5X1hROLb8vLEZGCqkhtdFLOTBBRY5nEs/VhDBlVNYYcx3w2O85BmveNFXf/1nNsPVEGs
rFb8Vq0PsS29kLxLw+eFQiIXZDK3AYB8QHj+BNmEooZV8oRY0brffNzN3foXO/3iijZEMgQUTn7B
nVtLliLE+UhdqeuVMlljKGIbHCAYg4/XUec/quf1ccS6OUEgCbgW8Gbzm5qXPJlOlU7KflCnYoyX
r9HX7I8Y70gZgmoyzTTxpA4kU8T5pPt5hNuokXjKLzlSU/Ec9pIXFroQ+9rH7DGdbfdOG0coPvOQ
G3Fj5LyLUYgUy9ogy4+E1JB/pnX63aJ5JbLsUvp/7mKYnGQViPEK9x5ohs/9fpPPzYpgq5wKff8B
MEtzkeTeR1Tws50JdOQ2otKFkcVWM/OLMrP38AejFyoRsgQ9ujV5R86/DEtjr+D06AkvUW5D5lIb
TkBgZMhj8QAMMYcSQiPeY2jNs0t6hxcc1SR07s/HwfAjMNUPMvrxHZA533vLIW0XFLCPQfzrhWPi
svuImNueGv1V3xrd+rMlUqQXjn6olFBlA1T2Yg6dTvBgj23hF5023ttrr5R20umt5RtWvELY1zkz
xotrjZu2i3FO1rKlLbVbowNJyS+kON+Mif6AE7Q/Ds+c10oN0SnujcrlHWDQ/f4Yt0Ar4cYCOTjQ
mgJX9OKInVkbfncU4x6yzsrcoJlDPN0YcUZLZNjkkFbrDgvU/j5qQhsJIKpBKCR1e+Vo1rYUFi//
hLEIX2sLJfGB2UEtBi1GDgpqUKRjO1Xpxfi2K4Oepj6p9LXtgzNT3WVClPLSFMFf9ym6c6ILHxNd
Qkxib1XfehOSIl1bUlnjR8+Ml4GgZiq/p5iv3FY820Z4Rypkp0g7G1xBU5pPEWBt6r+B068EGoRM
0ZhyFenKWlFEnwgLWXGgBydIbOfT1VJZ+G54giB0ETtIC2T1rlAIwnoxazpER4OimfI2O0adom/8
+z8TP8uYHagiKkP0BCqrxsljjPYr78jzosXHCH5ESfh4tHoS1tEi/3zYSKm3EGSbK4Nfq/5k6aSv
i5zAb5inrjBgo/wFiTOxl7g5snjQAoK8+yUMKGjwNyn7AwWYTLTRz4PfBtLOdy5bZ5gdKIby2ydn
3PurTZT+JzEmZMaiNrXDTJnzMfT0vFdBlp2weP8cBZXU7PJgErbrxCFJNTCOmB8woIeiMeVpAB2Q
dLN0BjNN16e/NO/d/W5xswxwRuoyL7aVaGV1Ay6D7VFYCxC2VcdjFLl4jRvMmzFtrwfPk8wPYui0
RmyZk0pIH0e1imN1rZorQuHF0BTKeyWvRMF1QYpas+TpRl8zluwbbMQqAAFgdwBE9qzfL2Ax3rBH
l4JrIGQnysvlHy5X1qB3kPSnRCtpbils+uwxvpmhD3usLEFcnMroA9FQquG0ppUwJIRld8qudSks
+KCp85HW6gWP/7/wCxF2JhWh5SAjAtd6PawiaMH+ggNeGjA2AGpCvLraRypXzk7CAF1wpi5LHOot
sS93/XIGTWx5JqHbQL9K7kIxbxnVRCeGhnxsXDkaffnc5/e8Wo/tLbgsJNaieWuXg7fsnJIxEvsF
PO9Amv8j2PGG+xewTV/FV9FXHqwJp0Oz+hUwmx7AZ55z+xAGwp6yEAuZA4meJoIwGJYHBNi+/Q88
btmpp8owLk2l7GI3jtHtZ4nsWdqm2eafYtiY2AeMgStnLJE9h629FyiXiJ0PPrEVFHOBk+7rSvzf
vBD2pl6ZQ8ilUAcaPSiyMmeqineU8dUumMtGckhxtv+XIsmUM8ZxBE7j4nXpgA1uHzo+GC9ZVc4A
dzpN+bDS2BLkyfeFNr8mSuQqjU91wM57e34rED6CizXjWzc7eEDhuwCncs9OtjqAyI9iltZV8JhD
Teilq8IoMzRde5EVzCTG4lZ+dWFwdKQ3lBPzJdjFsH5kuEbmLxrus70NApG9pwMCJTsPucyyBIzY
iCWR+tLWEiks9V3azbZRXvsg3clqogmWkJ+SpWoLad05qr0sBX2mJ5TdMQwXEPEiHcyUc2vUZb76
iql0mN4BLLJi6uRSBd0Dk7KGxqiimE8rE3AmguAu0avsZXz/F4QDcOoH1OHDK06lWNsNevBKvcPV
unvs7Q33+AHwAZ81GVnd9PrgBArDwMoo61r2IP5b9IUGSpBsNnAHwzE6mfHjFIcWq8NrAh8qoBSu
21NdTWRIbZDfRI73qXkEGNRYckjRRSRpPPEt1Y5sz38Q2UNCjOb2XCUhnFMhpymhxTUX6S0UQDkx
G9c3arhPN9dcP84a0kuzwv1J+iankSJrQC5iNCYcwHlV5ZOgDx8w5aoYBzsd+Q6Xu/K0G6SCJn2B
SEoezykuUYhYoCvTTijSxQblcNkucL5TpfzeTmPJ1hIglPbQwx3dFjV3VZku2yZrKD2SSNhb571l
iIwd4WX/nAzpSO3ArwN47VDkzh1cpZEnaLnvzhE5o3rVnLNZk/v3afMZT0eN5u1Krqk+OGNk3RIl
55zBRl4bUP2c21l/GZPy4GdndF7RJE2QbhSNc6Vej8dQfYBKqAP7oAI47qM2Ys+PXtyDlR0OXiPN
kReZxeLKpbybG/bAMrZv/NwhdaU/gIsg/2fG4ON2nUb0Z4Iaxt2p5OW2ZWyCLtj7Rdk0gXGer3Yc
K3iDWHvFCjY5eOoxw8YmfSA01gLb6UAFvfwf8+FMn5LvdvQlDlPZ4+tvgleaqq6LoaFSiWLIpWjM
qDn1csdZsv4ZogeewUGPJ1ECCnBU/9l+3bovpb/wVGi5/wa2f791DzJjA1Xwlwg5j4VYNwcI1tGq
VnksYzZm2WCZv8r5URM0FiqxMrS3NjYltOO89j2PlGThZCU1UaU7/EtzjHilbzdI1c8At2PA9K+r
TgH9iUwPcTMxHvhSsCkllulTMJ7Juw8TQvZj92MV3DoQjNi8RwjjmwuYdmVR9zTUqvsAV9P1psZg
ByFBb/XBQKq7S/B7/Shz0r7hl4psF9/lOtuf2Ir0dWjRIHHGcc9cE6Jc8xv+cOC3p5VEmZiO8ACT
ZFB96dKNAUaB5KV7jOMO7HQNE8VeQ+SZLZfX6iuCozm6LJnVVGIMkbM51d3NPFJcNCrx87ReojNH
oU59JqJtz+gWSO/PG9syy3n/lQ4wSkF1ALUp1+BTga66Q2ICGaOaxdvQ6MHeXspYggKYCEFhDzXu
58VrdKsCH7Oxtucwty4vcKJRlYdWCymcbP7xqLU0GHVjRN6TS2OFKyebSAzxuJg7mSmMyQeYlciW
R5OLX7ml5d+KmAzPTj+2CagZfA2gJV0zR7Ttjb4qacSLKk8Idk8ALMnAREs+mmAY3MsgN+iy80rq
AvgE+Ktz1eZILZV7ZO8n/tq4j0aQE9ZSEA/jNcaFfMcBy61M3WOEN9R+5eZ7tEiVcMlM0wpBIA8k
zJX/j6SqVCcvNlkmznpeO9zCX1ciGj8/V5Igtacc3SBoc8pffadcBe2Og7sohnBqKEk8UVkYnOV3
GRFTNmgiin8wEZ1kFgAMv8xBvchqBVtGTqJo2yiKqiUzMNfioo1ohK/X9rQZ5Dd/lOASfS4xksUM
o64/ns983vJzXIeyHfFTRCMAyx3T/TdjFWJl+T4bHShbzHi4hjr1/ESjnCPLLokJlO9CVt0rKPUE
7gdIGrCdwmXSVMkVtOibrcUgePyI23HpSEZ1nYYc5A86NBEdiTgV8HUqjJM+vvmVwSx3skGFaany
e01XFjuEDyoWzljuf3nQtgh3AKjNsEbooLv/KMrzdHHoBAPIYmNVsU9XRlOBGFW0xINUEOu75n6U
Ay8oVHuhyoA8AcygH7PzVYgavGBaki+P7MbDpFKsjIxML5e8X/c+Lk+XoD2hwL0e15qCe1ndTDT0
3jvDVOldkJ7Ov0HEkAt7j/NfWqExeDh2eohZnSaSQa73HpHZMEEMj/gp5AwqauCLLoA0pYsvwp8M
EOJH7oKDEi0swVykUycfeUX3yF9IMsLli93u4mcy1/+JJYMMxcqwTOsJ9Bd9fXbrkgE3I74B0ON1
pVa+bLQpiad1Ny/CYHUzXGY3Cg0lxcoS7YSDKq3JkOetnBPsB8gd4LDbBCC5VfNv/5aCH8jg/MQV
U175z+V3ezLj/+QbFuZhvZYwAYVQXPAo2fo4bCWM6ppSOEyzMlDrGzelAQa2UTFSXcb+Hsvz9QZD
JkPzSnOIcGvQx65bDpxiDgHF1Y70dNwVj4KPm+AaXpPLrCSrwfx7uOHGwkp0QFGiPmwYvUNh1fNE
yQjVSBELICsVls1OCXjTzWpnlAxooEgibxsXAS7lUfB8of3eMFGed4Q3idfCI7vjMjZzmfuyb5tx
dDwkAJIsVKcMGq5jQa3DMC929Y+jMyR/cecubmoelIJvFtKZ1KnPutof8lM7h+L+gAXMUJI7p4YL
W8MDbY7mv+pmHWZA/9/suA3mF3txHR4lRjyfn1Rz5ug9dxXvpzo7uZfNiryD4NZNsrI2yvpjUv+Y
UxMZk32MvArtRlCl7jNy8FofAv/WI2gt/NUkmOuqvU8Gw7KWM5lHBCf3MSbzqUP4XwX/IZI1bX/x
smSv7ycYWGz4ghuS6+VfGtxfnS3BlEXNjZ+s+khSbibbIe63ad1umMUuCQc8fduDdaG4NQe7l+Z3
N1dkYX1Dj21U0exMzM7hwlfQIXg2Ms53Yh8nA2RtSYqHVXXgkwNkXkt6Cbv+b5JLNBfv1bPu58He
AIvsKrmNPUWSLXDkK46COTu1d1q8epth3zS28CjzjxmUYmlPcQzCwqKFNUZzwALZAuOyKlCw/1IB
dfsUYaxJe2JdVZO1zl3wir7a2Nl19+M/lnmpglz7W+oE8+dAZYTSfg1Dif7Bh9zg4lwQHDCplCI5
1AfwxNS4tPtWZeZrfBoFHYBJ6CJsvqNi0f3l6PJejo/BwOIbMLpUJns4sY/+Ut/Oy8itoFKjokP1
8242pU+6WrzANPROMm+SYUaNlEXqfWj1lVY1vpaoMWKwrNlU0k+csF1Yvm2FvZnfxXSb6zhKighH
E+wVlvytNupY9iPk9Oldnm/l65pN8b800V/8y9uqEuJtqqhwppR+wRnpWTBhHoHmNsz08LkuM4we
E5VUYpP0mgC/S8njwlEYE1pRkI25FUXbUQC5KfzPyolgYugr6LDNfsuTZR/XLtfbhrZs3FTmc68h
dvyCqwyii+2vxo2SfwlMKrUaubkBlF3SR1RuHN49pSYHSOZ5DbSIm6arJDTN+x07Jl4AHyHNCRKF
0+eQ71fT2WQg1BPPtZzqQmmFr6cLmnInHh9t1CBp1Za+aTb2dwLeHoCygI++p91w6P83z4JiASrp
QvHdu6fI5kLINN6rZt3gCS06DEFOmOcK1q7lqxRPNx4NWyzvQmkJBs3RgAFKaUxopwwthEcEFGTZ
/vRwDBmkmnvMUoeSR8EFLTj+gfUnYmAvHOboqj58QlJHElgwgz3rjjuFb93qCdqOp/FSViuy+vv7
G2Jc/XJ1P6i4K9FxQELt4c7YPIelcpTfGwSFSrHCU1jt2u4tNOKamKEUIPvmfWn2dZn3BXpkcZ6q
Q1a1OM23Bq4NZyHGkjPa2F7c2wQrpGvV9+yLjjZUb1qMl3R3chAUa3EH4DuF1mI7roj71JO7F+o3
PXM52qPnqaE3SL7YE7qKRWMbd3z/twVCr1O5vUkH4qZyyVNk+z4L1MYgSR8VNkim4KQab6ooe7GK
H2X/wgARQvApZMWPg4bFWV1AJWaT0L3Ef4fEm+ysA7Phy7r1HSKvd4RBNngIqpy7mBL1BD57fQJc
BiijakuaSftvW30nbjNu+FTe2G3kLkEcaT+/ilVk1de5NJbB9fm8SNilFikRMzrkarTqfYpX7vIJ
RPhVFqNUnH1QSKu8OHeSnZ43oHgkLkemLj50kZ70lYleqdMfwtWTMekfGIaMJj406yvyzCaE6sPT
uk6PNasNZFtkh7Wh3Isue96AZ6LOPMP5ZoKUgVKAiVdX0lxcg1SJLZ451JDowUMnaNsfrNmrx8GI
6xk0ESZNB40B9d/R93f1rOF06IGjE/kmbBwj2JzmQQ9RfyzDDJBTw+D3GRUGljpEmei2QjfcfB/y
gnt8xw299OWqNrQuZxeEyRR/0UkBtnNuCCa5Xn9Vi88T0dN7QU+yg05EDW3Mc2s/5Qu3QI6Vp8NN
yt77ZVrIRsRw/hjIcND8e8A1RGECfdYxRc+3FuhuW4wmwKP/x8Y/ktHQhCW9OcTsXNP/aLRQ3f1v
0RQcrkxJKr46+P6ZtS/n6pbX5Chhzz9SaQQkp/TRlblZ/8eUrAK70rwleKsjfwP9ceOiYcvbUii2
eAA+/QjE+O2emopV5rrjoXR6uIaxcHQNC4SERBwwGoapsi7wd2m6Z/fPmw+Gj1M1+wQtOzR0XAM4
0/TTc3DmQD0Ho+ytOLZGncZr5R4Hb1/FqSMZ5VAZA92ARhENq9T3Rd/E/TrPOfCa0O6kqjNrNvRP
59n8maPez43GCwgMtbCo+HbqPaS5YQR+ZSnGJaS7mwfLgE1Wm+V5/N/w4XWgv6CjhZx225uVUgKp
X5rNQrDqQBuy5lre/C8T+MFvdiD807m2tdxyBwp8ug+i7j38BRc0j7K2qaxr+rl6L+VqLI3iRP5V
8pcI3i6oFRI+VbPy6+S+kUHEjIXXNLv69tJ6guf+4jZHy0Ky2dlTq7wjxVTzejgzXjH5IIgqrzk7
+1g9dvGsinqp/Vvide5+ii2znCci9k+B4coc7AAx5aZZ+ws35OvXQ6ZKUDxqq/NbMUMZ2L23R7Co
PpjwtmkQ+RcEvW3zj+ws0JsTMrWqd77EWu81T4TRxo5guuZcFsjZxqUD4ElZhAcJEOVCYMpxxbTM
31NgqR7GHBfk1tWUzqkTFc4re50/CxaosOYzop4do5nsTdyqw1G5Bb7ZtZCq0g+8jMCCfp5yR1GA
H6iYoKP4pASmwiXSLCA/5tgL2MvVRPvWmjIlrUEN2Jvc5yOQAfCwdtCFgTsxwu/E0M7/6xvxGMjL
hFLOKaBccCoF/3q3LnllyUPdzHIs4EO9FPTjynO0PFM61nu1gJTGRgeZwPk41E4QPgclZt4VoKPI
w7xYtQOXyTlJ6MsHeZX6L6i0oF5pOWYBnXmh7xZq4cTKh2h/Pt4ga92lhtk65XDpQe3iXlZ+pb+a
kc9EoHKmQmKNbBfQvTz6Wiw84GnX2t9gTPXdAvibGuYkIGWMxROMsnaonarJQs7R7GwxLlkBnTjG
eUuVkDfXEAHYqX+F7Hdm0nO9pvVOlvqvgocOiproINiLh/hnoMfXgZWq4bOY3YhNCiU+CnztJ+dM
9Imbog1VJqXCO5uBBjoNrcuTUtdjHUiGHh/fqFsRuAxThvbod8Z+tOZxvEDwjI/3KOlLPC9zcVrP
IULLsolRkgx0quHzsEPYrRZxWffQWNf45NafmfQoh1mbBhtw+W/KA3n6xhUzXWhFw8hzkOfeIjp+
0rQE6xgGwCCE3GYoBX4hDNyXhlfcF7krLrW8jYhhfcvkKr/m9g3oFtRPOXi0q9knrveXBUivom46
L+LlvEgNLBO8rKqRGX/oPWVU3asRs+H5e65K/j4NOUFY0WEuVhNwLXComg/6r4KXdzzNXfdNnGhI
fcJ5OcIRYyRoLCZ1wrjkhVMYxKE4ZjGiio2PfZpJbfvW/oVXBijwW3JjRt2jK6T4X4aQVp16uU62
S9zyyigK1cfy3TuYCBDxDlTG3fYNPkMOrllyYLDcRR+0eDsSkfvpBmM+1gn8OqXuxQBKF1CMAlDW
IFL1gxKpXtrs/CCsAXZUhhQHrL4es15pimMZYL7SSzE+j3P8oaukjamwH2TKd31Xyba33ze37RuQ
qNLKPanUnDOaEQwd0MEGwKTo1LOyFTdy430gJTb8dfili2oHlVFtoxeufZO+dEoTGejOTwoRJ/0o
FI5+D1Xbwv7wvt7mlWKlTs57Ever9cWWR0cHLsLFfMGe8sHytoO8w4XobnIk4U+HW4CCu4d5xHGV
FAseos1W6s8et9pGSxEIRX/yAME7g7J7qes/tGrJJeUaqGH7PYCB7IdZiS1kTi/GGKBBf9Rl6H4J
UO8ggpIAA60MmxKWeOID3uq3B/MIRUNpBMCGCJYJK3tqDV6Zn9BDsn0xyFX9z7jOwbLe+B3W0m3H
uv6bDQ1aPKxkgIRf0JcFb8iY3daKlSHAtTlT2mUeTcnDWOnRvX2gZfu2zb+HedGVwY8RdNhXURaG
ATbUMbMFaXqIr7OmKX/US8vUr9Reyvu7pCAn/CSUYTOvw2PmoVaOpdp87UrZT3LlvZak58IDAIPP
SW3dESiC0g5AjgNM+zudYOfUO0hSrR7AOzWWNisVdvV2puxT5FkKV4r+bOh6TvxocL6ULqvu7ceo
/6yxcDzKcSgRbjQ4L/wUVQgQoyEYLTtb7RoWvQe44OQXxOMuSoOz0JWJb/aZAyH18AeC67O+QveD
1FZXu08BZfPd7vAEsZqm5HKDVGbUzXSvX9Pc0Cs10ELhJCNd/ZxheWULTl3uJl7hkeH8Yc0lBZx2
EfbKTYDB2xHWXHgp/kstOLmlNmummmPJJKg9ZSLxwb3lEjW9RwA2AlveB1spWCXZpkoLIO+yRE32
4a6IKbZeYebFjrMtbYh3sdhBdlZBtmjJ7AMIXyCOOIRsVjp8ho3pC3aviQvQ8IOZ20ps0Cvuqhiy
S0HYtoIow0EA2vAe8Pagz0jUKonn9/zDGPWrSGSRnD7TbjuLJKnJiVzT5IqLZkuWQJwybulec3fT
YKgObhMJikBuwsoo1NVWIJgutro/VIjdnE9gARpAVY3vf2qs2YI+1uOWppEWh6BWgkR2sfnqiXgr
qAJoRC+Ey4taa8gn7EnFpJ3zUwUoaZxti4ZbFSR4ueLW1qVlLhlcNy3IX+1YTmj1iiDyG7osFv3K
pMZcp11xY9pAsQNIdjf9JjbDlBD/TuiWyogQuL/Hqn//EF8pmoZ+Ts4OBk+UPOZYWbO9gbWO2lFe
WqIjjUL5fCP56L19UzHU5vvhVLuotsFiITNKj5lzrK0pNWjjSH9sWgF/3t+hCzEvoG7l3YDbAM/w
QFcgbOokBwyTodBc1CMp2QFce+WkgrEsiH6c4QGMxCHEY0ZDl0bAiDugIAZCEpza+8HKCnPblluo
jZPTzgH6gkJ9mgUj2Xxk2EKQyJ+dC0hDwnqFdjCgbuZyIGY0EAgvb3wuAXL68a+MxToVf6YQn/w7
4fr8d11Td+7qbLq3opqAkMYSiB6rOViB+EIUEwn9xDTtTdL+jFpLIx6Kq0BAbWfvIuN1l+BbZIH6
2nMM4eMNIagl0MkmLwciJTdTHIZnKeWv5AMY8xCFtZe0SrRIpW6d5NiEw4uOxz3FbO1ffA/t9jnE
RZ1WdeBn2njCn5SfPfNbcfHPeaPEEbxObayEc18rHZs5SK3FYIrLajB1UyOGLRXWUSIJR78b5yst
YFip30ywx3ZXa7N2BxuYXhWtwx+KdYNHsKOsyC62AU9z4Gk5T2sgubWwBmPnG5u1q+2sJFz7aerv
HatZSHsEWSiWi9HqYioOP2RR3oMX+Qy6JOnUU+qJfo8tLPBVMTCimGcXLK84Wxl54hHPp+ypC/KI
F0mL1zHe1CaAYNte6O72mHqsyaSbNEDXDX4qhA9tjrUeQ2qvPgvZ+mSuCfoD90tdotXvomw7ji5x
/m3zuFrP/FioWknmZXXorGnXy6Uah7IS4Z1yZZc1USbTolAAjHf+R0Lrg58cRJ2Mg6faJ6yn1JXQ
DokYsaumzKcUI898R3bEDVJ2rawLace3nUKSagTSHQOD4e5iqWDpAbhcpRu1R/WQaRctofnUijnM
NbiO0XwVisP8ikrVgd/6/bYsQnNTgWhXYD9YebsMqHp6HjvFc9keHJFXOzhfyrAPAMIo+Pt5Rqgp
shNRDS3Z/6HLR2CS9iWPDQIgPokGGvxuowPLGX2Pwnpt+PqcrgIDTJOUURZBNOpvyBuK1QA0cZTf
taRSnZ7BbSpm08dOdpJwpl5RbjpArmTsmJVqN1ASn9RpiB28LTdFYb+fW+dQk3l/WCbtdehebH8u
H1cbwOBTSzPuBe3I1xZtejGkt5PbbQVQA5YgDZQUyqCdnwEtMPwaLIcQJAdo3Dm3dcdtP7xZHNrh
WRZ0p4U8Vqwf0cMVjf2t6iEIgwWUl5zWxaWOoln7aUm0gEOpF/f9pEBAPp1jj1tZRo0fbwHnwAry
b/nTBs2f3RE1MyWzlknSTiAZW5w7EA2Jss2VVfptRtsG11smlKDQGpePzi8tuosNf/zC30p5m31f
YsL1dTIBSCtNisL2aoZ6xJ8Rq+0jbBq55AZnSw/90Y2NxivMF8ujs7uhFvUM2yTbxteQYE20K5DJ
crjmajpf1J9rtor2daHEpAMwf6QVPm6lqB7uxwJUEmJnZTo07xTR960plRJ8sDbxQF2HU8LuTmWj
oJ2zOGAiBhMhsT/bTr6Art0NaO2fXqfKMaKpXvbwK+bS8AE145ycgVFD9Brt3GL++F6tjIvFz3jy
zKAQNQ1bBwIy9snddX6rT+LjwFpVPM3fzG820+IDudCs4fuhDYDOjtZvPDx9+dUQbTLAFnjoH1dC
p0L+oMMEKzDYcehvIHAvz7e5NpAAM4/XUQTSFOZ+BvPO8WNpDnElwsfWtsneNeyq/towNGipb0Du
z68Irjwyq11duYGRcsS7ptdx/K6cx50ZOVQBn6jekfLEj5zYeYKTgfUqjvNE9PP2nw6fPPShM3mY
IDsvc7EL24yoZl9TB9Q14VFwEK3lYEpOHIjyzN6qvywj0Zh8m0k+70dhgPy3k/6JMjaLcoawFUTc
SOTgfmorx4IoRFr3/ffijQBS2+pIQzqAwjQ3mxMGDBTRvWASI20TbZ/BRPGK7i7etQSnCQNjE0G0
6LGnTMBYUnmM5f2KDTJ8aHAX7oMH9U28dFQi9EdU9ID3/q3C02JtTaoWQF+M83ObgreCXVpDQI7+
DoBBNtFLMdbuYGnrrRj0VTkl/wRoPiwaonyCfU7Y9YEpoZFy4Zv+8kSFuPqPU8PAx8BpTeeJ/c1a
Lz3e8UR4c0qNv3qa0NnNXq8t3fPsD3UBo5odptsfugAJVLoAV72gURypSghpFgnlYtgZ5dqlnqsn
mFh0BqdD6DtvyxE4HyRC7I6erlSyqhVAATJs8WD5tAV7TlttQlcw7QvAEL+V9SnXk+gZzGKiipmm
3+iWqgDVkGpFcBaF9qxuxqVhFjBNNU+wg88e+a+fspYD6YLEMv9sen25FL9fav6P9Sa50XRmhT2t
YdSPZMAwALkofWo6HHhUAMvDPQxszQjPbATodbq0EDp8W4JftkdHWapp7Owv3RpL4nWUcl88l5eB
l0dHopsh1eNIVZIhOZKO5/je0yw1Euo3p3S9NKm61btpqvLTsBZiPp7J6lUXwztNkShNe4zAeci+
Ku7MJt7G/B8Cp16lDpFLhEjM8vXkvzIScknMcSaq65tOJ1wspwIJjMxX0i1+ijG5cgW/bMQA2hwN
Z5xJ8vhKC5MngVqC6aYk2bQ2XTjyxB8E/REi3uvnBH8nZGZGVyWSQXZUJbA3d+MuZZm+jNbuxVbB
A8wi7OiAi3DuApRM03VQQ/J/4303xeDzxYmTeSTtl/cs/EDRkX1sbFtOIsBuwluAB6N2cAxtoSpw
eaujGPi4dmWPKczQc7NQ0So7JiT9ZqOVeMmCAMKucGTjqw/+caZJrI/rBT+Gn+4Ijj/Zf/SttdgV
SZuC0SeRAcIroY64VO8DtfnC7ppnv3aAKn3lqRa31g3rFiD73k1nxyMj/uJv0n81+0AZVEIEp+wx
Xir/V2yHfX2ZNW8FEgp0yI74JpxRMIA/kN0wtgjP1Acd1bVwdPxBH75TH33A7ce7wcBx3DW+DcBn
JhNSDy/rWe4JbfU0swgqPH+bAqOVnoF9JqxvFpiW7ZQXuf8B/won3CNuEq3GkhHJcbiMba65YkKO
TwS9gtPmIiLCB5ro9TOVjX32ZEaoMhDGa1ER9ajEdkLmPDvmIPQIsuVtFFpg7a8BwqfnKO0D3Nk/
x/BofOUwX+4nGRm7WznP2pDZ8q8+4qnuEyQjwev7EqOJQwS0G8TIuXyLR3dJm+GEOIX1yPJ6O/Kb
aQGgo7/xeYIweBpm7ujxeZPLxVySkkSIFcjNuDOZSbiFevfENY1Q/FRsOmQCvHq0A9t/ByzHAyxc
UGqtZgktlubmBqR6OVm3s/9o5BgE1FrNRcdYuSNz1P9Z8Xxgi07cnRcj9nxAtJKCGSHfqVGo85fW
/K5IkOfrZ6MbMIp+7tshoEyu9CwNnOVRouF1fMWN12DxQTTVu1XK14kR+qdxYNsYEqsfXswMXdle
rcWGpUpJYkzql0kxdKL9mMmmfPiamQiZhcM/90uPy+YxSl4G+jhSzcZDo+ULBccAnO8GwKrlmEMc
jOWRQ+oZbfdgc8xBnTQBYf7ohsQZJjVb5Y9DgSqgHCrvh9lafNpBTvJaNHt5Ff/8a3k2QC7//bPa
GjI1h/GY0WTQVNQud2fTHdukVbbxwRkGcYL3u8HqDZvRh4jZpNthErE9UaIWx/4+rw4EEGULBusz
f4iQhKsy1LJZPBzGBt3j77S5FENgk9JE9+1DDwW0FOqGDOtV6+2vn/n2Osh+5PbgtN3j/1Vex8EL
TzBhy/Yrsn6HBVEVVX/IbnrbTRGy7S61wcwupQQMf3dil3YB9oyinB+DKyREa1OTbiqnQOItbYhc
Xr0kQgwuiXBrKGl9T8BJHb5GEWMAqlFA7EYq+lhcfA0H7sR4ABMUptKaGZz4Kyqtoh1H/X/9jRp3
iQgPg0homZQY1MH1FEjV0TQou3Ez01eE1BU8I6lxFREUbz3PYcDERWUHqijh+2CQbYhnh91ZKi7S
3p9QTp+wRXX9BoyM38lX6laxfxZ1a2BlBLO6N7EcBtHQLD0yyLymtI7UglugsP/135FJm8OJg9GW
sPvKCdxHn/x01hKKqNJEEzf2b+cquZGVtsYZRVprKMibgO+ZErgP27HwINHS+5xOh6YhP9K13IG+
JD/tQtiM7jG6bO1EBvLsO47H2sVFTJKnD2qy33TqQ08nEZmLXcL+8551p4MU31xsqYedUKggz6Oi
YHrB4WyzBGC9cl5ovtt4xeiST6st6wXFA2hdgmTxPhOCB3i7gZOt/hjPDyNxg/X13aixNB8bQ9EF
8dfhqDvihQ34RY/ztakiJI43LtYGg3dvNn99OgzXKi/2QNHlPwzU3Bh2e4KOfp4PQfB7tCSpQtjb
g9EqWnl8lZGzqeWRrr4MiVzlWBJ7TVuBJAYyeRc2xMxbVDO67cY2TPDrWWzVKPo29CWyXLDwcLEQ
3Z15WEw7PsaBM8rM3+Z6IF5oKMpT9PoNmBr8FmYEYgHGEc+Q81pPhqDoG3GzS82YN8G/GgOGJg6L
iHqd+ME43iRezGmUOczpv1MKW2XdTf8qXvpZhbI+rMi5KIJVZjrdVFI1eU2ltXXxFHXgUGBcUSc2
qIv88LGCie6VfvfCS05PCGGLSg/XTjJ34VS1d/j3fukChDTYwxF+siLb7CT9nl3jw/UL9SxnFJ2X
ZbIDBVH6IP3owFcFICyukJPXDtOy2xsn75ZqQgG+WD2rAnih7BltuAtDc4PDkJmapTZkaYgdQgkR
SriLZi2VJRXBSZsErPBRGE09+5QCk6VVXLeTALOVypnbdVS5Ne3VKzNGmI9BzIR0LPdy+T+voOWv
mFq0kmRRsACSIxEklFo+ktMafscUhVL5ek6PLDbxXzv1he1xKt7D7S96hzlRDEhozG4UBEeQlCHH
dBa/Ap+EDbC+klYxQb3Y7zL3aUhTy8HGr2QAn4/ZpBPWXvw1/QubPcC4U0tzu8oyCMF8afA/8CJI
uTZVddV5UHlKCMPqfr8X8lubb2jB2Ax1OZgoV31fa6pkuzWJKgyzj2OickiUDE9wvO3jZ+sdoz4W
5VfafZOOHKsAu3mlQIp9ahdPJuZYNY0OgZXVKHC1CeOlh1mNA3zi5ChE6Z4pYjqmLPvVycVejWPv
P+YPdCMwge1OSef/chVfayKV0/OKFb1rZpUivcqkkHvxKUxcWc+YTP2tG56QjOB4VUkVI5DUkuaw
4c3CCxv9m7PUD0FqLD/gvzrhxWhZJXHzHSmWDdAzTt2iOtHP5j1a7pCgLBbo2damlwmh8Igl6maS
y5uzPwUDuic1pvrReV/pH165GxluwicfZN4LrDjVBHdZzdDBdkUST0M9wnT13ZkkF+eUlQfY4+Jp
jk9Aubo3ZFlyZtaxKapR3G9lDW+M5wq0XbS/S2VsIjMuadAaE83lDnlNYOf20RE0e7Bpqy1VsNEU
yE9HwR7zWsQmzZO497bYQnJ52Ok5auHpdYokcp3PmwIbdAgwPE53FB0Y9uAPUeJths/bj+swFm5g
v5vD9ca8tQT7mPD+cC/HRYdR4W0GKYdOt0sXKc0XiJkVEkyH4qCnmvkaK2eab864DKDRBIrashUW
oYhs05yJJF3sNXB3ZUmq6ruxLYlrSQctrmP7chxbqxYqxYAYQl4tqvGvtzj4+ac9Zph9wd3L1bxG
48mAvWuuqQmPY//8O5XQG1OUQJsvJj4MjrjE/YMAS9/RolkdWwAs9pBhHMCwxUuTHpJpgSfzoWTq
tyQ1M2NpRrtyPgu6l8k50G2oMIJmJA4h9XslgdufrZK2VaRzczvgz6z2Fcn8AqhMMkAZBNZBtPBv
pVNEbnPJYR6b8A3ai7LHTY3iRqx9AwgqGKKLMT8SzCqIO6EZmRx+6zA2QgdSqvSMvGGBh+Y0NXxs
ktSNNdRGuZpWGod81jrgU0bw2mnCzPkDEiOVB/fsR0stHLlfj0w/kzac5ga2e5zCDpAWGUyWH5+c
mRCeemaDqUonCoSoh2t2jcUTrDasFl6fxsFAkwVfPl6imDuxTxwvJz5bt4WVjaRAw3zTSPXg6f61
3PJH/F5mAniCa5AcQwX62Jqo2HVaAlMpJtI3SsBA/SskB/RVZwGMTFw1yJinskdckKAQU3iAYv9l
wu3sHSBLP7XF0n3bHdoIQV09mFceHloCJUbiCopfg3eWLMZ5AjUb3T1JBqzUnZhpXm4QhPAIcXyI
GRSaYNam4tCQvIrkkctDsT4zAjxOsr8UNMYHCRS7HK+LQllL07nehgeFAYf61aRXVDnkhp/YKWuV
j+IVbTkO57KviWLtil/zN+nwEVPQj4qhYcOPT/EjTwuIWOsx9LjIdq/zRDXgzrploy2kF/iIIf2/
Mj5kA59Kp3dcOL2uUHXT3GnNTT8OZf05RJ1MYKscU8fG4/i0c8D3psBhyzRuii2Hx+OlSCbz+3DI
8O13V39+2nBJxeM1CjJ0lZE+zuUqec07HiH+rGpYzAlxSXm2qyQZyF3Yq1dTZWPmxO2qQ8UbdjUN
pCwig2bi8grfNGi5b3v9mZetZ9cR9bqXcUfYZ09Ta9vHMHus6NtEE5FNjxgaa7yFh6vlIvW3+AD7
SAGD4abwZPHh08sqrjXORLKAB+Jstboi9sHR/3zM4Dhs/gFb8Mu3oeS/g3rVCJjDAas606DDyXj2
TBeapP4scR4SvMgLE3IFUmscEJjrOCWlorwWZ3i6aqPjuNPYcrek1zfEGVskPL448nXt5qPUjHsB
InqtIQ0FwKQrwUhd3J5O7S7hcdN7pdoJ7ferp4TLUoevCLvfJtceL7q05Ty7BfgsFLltFmt55L3m
O7TAFG1rqonlC04o3hAk4V2yoqVGTaXEegkxJhW1tHXvI28d/reA10v0fKTpsqE6zL1wtOcM6Ta/
pEzRZuLAb+we3qfYZVYlfsdOzfdwIm+/ezRoZ+dJFLAZ9ntpJZPRM3OlNu87WcI6cttlxknZD6pJ
JDDCm6wCpj/6EUUcTR8wRx7RiTyZfLquE/pGHsbdS/wXSt1iSkZnirR1JMEzIc1x7FijVkp+XxI/
cjoS9haLMIhhzQmq3mPyk387JtGplFzg8DC9yNJgqVi2yN0qbJWaYe+Gk3prZVD4Qocws+h27wP9
F7mScrig1rIvSMdq+NvF9tYBV8XZmOs1oA4uwhFZ2SZ0GThjWx+KwGzQdq2S4gYVzt/mx3zoGmbi
6BvAXfg83bK5Hk5CrU7j9bGdNUKW/ZMTMa4zq6qvQeezz5UN7lMcXdP+SVT1MA3vaDLwtJ59XepO
jkTxUokcN3H/R2/GebveqUPQ7orCg8mzlaJ1fBKQxE6tBHwtnofsYzZyf3Gkt9CEva47Md5Cap3N
h8AmxoEnK57KzEhLgpJU5YXms95FcMBlApGNRLo+3CyNiRm+WHmFQYjYPA8nBJPcj17Du822ETx8
+wVePHxNHms8MNpxyi+vtSAeZbIqb0s2wjGPBjl2Y4i54b6P1+9IlcXZycSZBvZTLFb21OZFhMEV
iCxtY0brTHWK+HH+8zQpyRngoncNyA3+Y8TUAYa4HHJrGNfmtV10fTdhqaVgNj70R4FexVaKxPun
h94d1ICzoDjFd2WZuz6XIdyh8oUZllhNIhJEw6SNsoMzH+elVpeKKGVaMpHACU4iZpd9g9WET/iZ
Sg8qCs76KPu/2d+6pRen8LDCfawfkiRwQsEShDkjduqHU2mqDItTYLhzJTJXiRbt77YtcGIA8dHE
POktAaqbT1CqJeac5Tu3Tut3IIfri2pqMHR7o3nGKinA9TnMoe9inh3iei1ZkSZ1GYX7TvqeCR0C
wjYqLAXqUcfVRtBBvoocd8bak7/pbuOH/Envxc04peHF1mHZZEOYTe4TwqIlC5B1CLsUjeOd8sj4
2t8Q66UCyv5ubxulokazIALp2rtLMaj+Z9vZcEQuGYlsphC+hDz0txVtsMdOh2nAPzqif4CRTCyN
QEcaermdy67NMITlmpWxCJdpD+QV38glwPPeTrkmGpsIHuutiHHv7Bi+Y4vbgGRO9Y0GqCEUBLMu
qx54fW2gKRMYKg72q0Hu/J8uyCUbPdsuOJpSa5+5fQT2uVj3szMZxxnvn1BuTmwHIXpJgYCd1CpH
938fO3XibtoDJwHBi+6NvtUD53aVyHuBE3BG2SLFIJQujSZ9aJyTxtLiS9ZEJA1jhJNDbRSAdooV
t5sIo4ggz4YemmZojNEzja8PUYCsVz/jtRnHtMZCwdJEowFKotfGH91JCVN60CiTdeH6jaq2MHLT
WLlln9QUK7Ek6EaWayeUCXuxqQ4YfCklQ5rCXJ8D9xdINdcYX8esU3IP+Vzo4iHijVudl4FYpR1K
0NxIg+FHMrCaIzhFoPaay3D2hYYgczmJK/4itOBCC5iOrzVJvhYtOJUV+WCFocUo8mHUu8n/9G52
XvtGMVqqLxU+DfdNoaCA1gfJFJyeiLyKAACWR1D6NOFtws/OzBr24b2OF9Bft6Zf3t7meX0xAWz8
dupCr0X949qu4fkTE4UxgDGPb/mvGKTWRUMQmLW6QGB9iDOIXBZW5WJ1NZhTC4pcZZC9itMV/hFU
kipk/hVvu0IMlsA3H7jgCBUDflxjeazkyzCVWhe6rXyIZ+2kRysxJHW0I+eMeNg9nRsLsD6HZKKQ
dIHfPobyNpMnAFsT4Mz9YvnSAXXgKaON6b/cDELoR71QshGFn8gOEqXJpCqYoXcIvMT3/MZMOCMS
XM7ZRgk4Movz6t190kU/b1JuXsZFb2bjSV6DJbLYY/PqTwU/NyIksYpMEINEqxtVV25yQVvT0AEg
t8DGAGnoCKKc/p46ieU3S5cHqH2Qavaxow+NvxLGN2/OLvZysHjnlLkyV7M8lzVlJTFhECU9LZMe
d9/goe4ANevRAtoiuk24kNjKXgmM3+QhbCIAEWI/1yWORgV/PvYgXyoxBDS+6KxRkUxBX6+2jFdI
aNSS+mLYxnnK8OXLyKBROPv7va48D2mGqt3Fjd+uHwL65sOACO88Yy/A505Es96fhVcuPIEaCCpf
GbJIxgZyPHz+vlUIpsYj8NDsae4jjQjas00/xLnQH1olj/m5yPbiYRohw4b3nakrMSib6huLjASp
Rve/TdYyXFhMS1veg4Zl7Cd3g7lNxmU0Zv+c/iYlagSQxVQ4/NADuBebldFiiRZYmCYFYncGKwN6
yDVi4CtOKQyQuh2B37Z44QjttAWceyEqdv7UJGcQ9bstM3ah8+Vt7kBDnEeQEhxNNaGmiZQN9P5Y
Ao+rleEpGaZp0dq/63T55bB6YbgAVAn8E21mTLULlofMQkVTnueMwRVgKU6SACGvKaC1E2DCjOYo
UCILohYiC0z0pUHaKWqQsUxy7WWPodKQQZuCUo5Oow4vDogFViMWVIe41imWnzqpsPttXpU8Rpot
p0YTACk9iwGA9C9Jhe2R0TpOtNiAHCSzQl8MwggztSn5P7tTYY1EI32OimN+1PE85qYGO+xODENH
f7PKavnwsoNXUE/M564sMkA0SJAHFzQjulpvDElzANgu8+LImSwCIZKm8mkAD3ZBDypoGjreah2B
CX0oBfroUdyhFfeSEKtqV8RxjtoJOFitUeRct8W32K1QkWJm3tG8bpMEpVz1mc7CggwUrF1Og1bw
xHsmOGmMDsCJG0cCHfocEa4h3qMWqkYG9u6bEZrxZ17c4M7DQ8rSxeBYrLrC5zaBBJuwi/GQxdiR
lMSlYqZ9O+Pn3l/LhSXfdiuKLnaGwphoqjix5ze3Ap4lQe2U6z3xt+WU8y0qJF1/01XkjTBy5mA/
vfovkBd0MbKCMRA8r97oUCDM+95YHTp+P62SlYfTAc4zI3TRHo8G18RsxjkmzOItpMRigSycU6Jv
yrjNtZnqUD3zXopaw3EOhHKFGio7Al6Q9l9ZXcamh55VWRWCY9rW5/vijhE2pFP8sfFiKa42eWcy
a3+4POp24JXYiGRFWjg1wjJ99vr+CUTLT8FDhkJ5iZvIGdZg0BFeyiZeAqvYWrI4FbLNN3UJls44
oSTpCnohusEIKrVMWEekSKXf+N6feIOWSfBJM0fKd8zaA5oO/QLimz6kEU/txsZINwpuCmz5RkZV
g0PcGj55XNYGFo79mVrox/G8GPYax6aOFbPWlhL28RKvBUlbAGcPq0rFdFraTbSauYcRDuumEPs8
iGz2W28ut6Dv4ObGTV3eOe8fi++iytft7f5MZbdwPdpQGA68mx2rX43hikpiYwjbqeEJARyjkK+U
TTM53VRKf97i4Cp08gMUJX6n3HxXu/jYRJ2cSnG+6XRTrkvat7l5+0XS+2YS+BKGn84zfT5XJcZW
V9CYjRulqqgCktPpuhXGhfwqvGi8dqSic1cvHRCycAl7Gwc0NayvEfFGMMj03yg3/7N+i3QHdSKF
NCH5VWBaM9JOw8ltOyuRl/k9zB1KyBFmF81TmfkmOXvts0+lFU8ugJcj5T/nbeGzpn/nbNeB8Lhq
01D/26pGZk9ywNhs0WcaPJAAp2/vdHcPkW4GIdfWH6I4EQsMG2GA1eVGel/+YVDWwFDlpVpldjvU
Yp6YkgxjVmnQGR/YcuzPXceyYp08r9WrIN0LmOoYn2LHkXY2VFiimoZCnrWMqkgdZFB7oO7kC3bi
QiN7rLhg03ycqBEOKwkIuYKOEngnOwatzt7Z5fKecmuiWEnQTCO5s0TmV0Sdpp/4H88H0szfXNKg
ADkV6TXkzLw0lN1K6IPxYMHE5rb63Fds8gqXxZvkJD5BZgmxqiFhoWe9yYb9pDpIcLKHRGb/0+E/
p7bpR68Tc/QLPYhX7T522E3VgTsHg6TjusC0h6M00TQS+bOGffioYsj9kvzYwDwcsuNtlNzM2rDQ
IrToL6fNALqu1B1Vu2ZuTgO6bReSC8tTVunRUe8gSXGNr0ZsjjFugGp9JY3zLoaA1rR7cfyAHnoH
s8IqYjn4aPe2WWRbTUn9LVAIjafuN85mhF2OCAa6HLQdQJO2NCQTGosw5TkL0VicVQMjrU/1Tvxt
HRY0CodD5C1IA1cXwjrtzrMdLVkc5By2KeQkSU8JaCaFmTHGJsrxTFyqOAsxOJin4LRgA/SZnGny
lFglMRCREeX6ueYoMzRaUYii4ZnlXjVcuIuRZeEKsIeweMJ+pz6djr/ZdWPm2gCnCaV5VnOrwEPP
KQ4AJg24iJI6FgpPFCqr1Fjo8nqDo8D5wexISIMvQVCXTbXC+yJQsT5LUnxFrobyIs9KCZXwW8RI
MM/xpYsWy5lJd5Hx3HptdYFWabwT6BBVYDAXWWB4FsFhEyUCwhL93sv2g5YOSmxcQuiV2Np1398N
W2Nx70yvixSnDU6F2rLmQX3wSFjRzrCFldjO82Sk89EqixjvE8OdD+4EFaNGT2KUwA0sGweQrGGL
/RFmbqFLJP57hrHATpWHJJKtXPAeu21AYfvR8Cvha9mNynV/JR7yJJQauGU0TSJjNRPUZVSI+ljB
29Dp6Uid19dlN4/1CZ0iRt8oYvou3xvecqI7SSNLA/uzazJkCpi2CENtgC3n9Hk0C8W/otoIWEM3
Og+pq+U8HYClSnpd+BU8tfSafj4Ky3iQzllKks3oUNRXr+5Lotu2Y7kiVv//2ZXp2Q0y5FklJUja
2aye8mEkEL7VDQrgNRqnC9JM59qUE3Uwrk8MAoWScrHYFr9ko2MI0OlK6cNlAsfOyzIgpPRUq7MA
CgNUMYaDrLpzj8t9yr/key90xL559iAauj3DY8apnHyEMKPaPfkuZ24ImIiovEvMtFMp8+6R7blL
nlNPMemnb1s1gi6a3mDSm7qfKpwfUhlcKTcIwfhS9pT6X/yAdSRB1dtBnMuXe6H3459YehxuKT2l
J0zKQgHsfLxU/LnWR5iFkcjYU+6pvUne0MfT3edZXrDhgQCLuMtdkrigZBCGTSKzzQpGHt6sqV+/
hPB826BFSoG520s/Gf3uORzk6qvzFSVgq8JI72nHbsnIOmhWkrxGfZkApMSaeMLADB/ojz0W2ozH
zGS7hK4FKo5rrxGSbcKwQkARY3ihyswq6U2L6Wpu1iOk9Ceh2m142eoZuLtxBjT9ruPn585cVckC
tjP/gXftWZK/wdmF91DeECB0tgdx9J2z39hKMR+GUN5oWmTdWZc/JIaB29sDCGSXf+ssZ93B2cgJ
zopltRYhiLuWaJ8OVDTT/9PefUOwAqfvjSUDKCP9cFowdagAq0cWgJYnTQCc0Cw6qros1/Gh+XiA
V4T8gGo+ldDP4s2s3AQw6UsH1FM0KxHVEctWsXEYl3QwAU8Cb3KRK1n9VgXcqpQ2Jjr66bKPQjPI
Vc4Xx9P0SgPDJr0hbo3ZfA3SmYiuzF6t0/gfDgPTY0S7IJjU2bLicXHoPRF01zX4sWojAsNqYsZR
XqDWgutEgP6f1g2e0L/bBVzkEuAL6yUhaoWXLib6kgb/NbHmVfcp+5Nw2ap+Q9J1H1iYozib++wj
Yt+dTryrES94se0AKk+WA/KfHeDPy/fTRsEzxGmH745oWAUz3wD42e8GmMtzWCs/LsuE8TTS92hV
m80DvKdFqVm4lbeYpYiwAoqRLpjNs/DYd3hbzRCsgZJMA9NkCaYZo2BMAgqpIXDrVSSnpdXaH/Ru
Dx9CJKan9OSvq1MewelY0dXv9v/HXesHiLxUsAZ69fR0ZVHWv38x5lDw4C1Z7c4KPHR4hWPluzlJ
QaJuibjXLc21lkgVU4VxC1KPwSJWKbwXh6sLlPZKYeJjeWVMP7sThA6hZVhxUUfb6HxinvizK4tv
iE/dZeho+bCD4P8ZOI3Vr/AEN9fFAvscHnAxhHemx1e4S8in0ro9m2XXnxvHS3FHtQIw/m08c3Jm
SMppNVCINVjwpOTvuVvjNPLMou32innCS9ZzlJO7bQBshXyS57YmDIPgMlNVBuVtG7TdB1sqyIGe
TfD7UeN7h1oGSI/oliwYUWjsGP/pcBDws+k4WVPBMMMh/pGpWiQ6Y9otNvuhkl3FMNp3On52hPHV
P/UlEEMz8B1tw8OKgwrBm095lc9S7gcg/xEdWiiq3NEWyz8jtfBWWfwd8AHzFfywA6aimNi3s2Ji
gjFeqK+dYVzuiE/dtgfmlGSGN8+n+wpk9Qvyixhj1D7WZlDzfsUAD2Cc8zpMU1ulC/Ix7F+LUWU/
i8V3X+0TxA66SPD8PcjI/MOQZCKZMPhEED4GOJxocPoqbj1lLVZYu/3EIpBtGYRBNYI/f6b2ZmJ2
0c/Pj7Xgjl62aIb4GS6yJuGWfMOV22tDG81PYORnAGT7IHYQ1UNSkuMFktt7gnwdLa1lsa7p/HzN
P74UX9MBzZe21B9T1IWJeOVNH2iuTKR7Z+nYs7QecnkIJcJ4iX8NfzPJHM1Qn7RZYZcCrWsEEx+N
qhEi9u3kgblZvVwAznruY8Was38RNDvaDqqLO7ixcEJr7AVX/dywrHvA3VL+CCSwI7TGFz6aJKvN
GlNSgI2mAIIcpV4zh1Bl8p56AHU4hPFwa+P+iJ/gGVaWPVAmNukmq0IJ6nrLSjPKeUv+OJuTMpE+
riASdLc/98gC4YNrdRHpvr8cdVHXrxfLxiDcAADXcsob6NE9eDDjnSR2Q/fTHpbTtsurpjMGszFD
EDxWRcJZxu4zmSm1Vomih0I9kAZ81kLyNEeRmt3DS/dB2ktnMDPVfsn8/bDkpMF55z3NooJSWn9D
5hHuSv0UlOtATJ+z9rqjiPg04jdyhq2Y9wPpBsp2ZXkVJPn4nEYDOndpA8XC4Ihu74z4rJUWw3uP
GQUaUxLuQUeAPIC6hzQJxvPb2vcaSL7i1T90iSgY+OMNY81Ov2ARIIqdXr2UlRzxdT2Gg3DPqsgj
T5yPHHR5mLp+l9dC7tUcTXDmjEtqG9A3fJ2MS27hgL7l10u18Noa6GOPyad/e+4C3UtRooXEjM0z
4IGFNWwPLfyqPRpO+TYuafDyI0OouCdi9T07wtS+NcV2Ja2DxoX/+UKDjMJU3+ObSVvEn5tFO2x4
4WJFj/rjcgd3V027O6iYHIfUQBxgvLbq/qWTg8+C4tvr3i25/s0TW354OkcTVkH2wsrfGwbIR9Qk
N2P8r5rDr5nKr4ISSypDdeLViChbJ4Sp7135s+X92M7shG3LYOBq/i3Htmt30m5zz0b2CvNm0a+R
wwEuiQ6YfKAZ88QHgbbNZ9YUy206ILrisPUiTa58hENS8hwYAZpJ1UO8wFL/jrt3xGJ8RrWZomi2
PQkL1wwD+asfKGHOnoAUskbDeKSdvW9bROqHl1JqdVJSO69v/HsSsNrKICSvDaiMGb3+5BtH87FA
/z/LvmSt4bBF40sBPdMrXyRa32adf+b04iRg2op8oTHiEIiHriwmRSSgpb5u4PG/vgtbKr61fID8
+Ve0CvZ22mDAVjE30R4RbzWLnB4aYK/Bsl/7+v0IuyZOxa5J7ciY7aSYsCk3JYdAuyD+2ciGFxa7
8CX2ByrQ2Z5gMwVNoJU4ZotGNN6f652lSy2LuV/BxAk/DA5UTUFDaGRl4lCYe4d9se/9jfbxB0JO
nVVbqPmAsgd7RwTiaaNNQ2vtx5XdIotFFeXGL5Z/6LwhgDaJxzgYr+kb/vA3xWJSHX2SXSrpHqyF
uZi8dDA21joijtx9pQKI6wB/uVq2gWQcwvG0WxSLv9XN943yatL0ZgwAkLI8AoKQuYbCsMjIO2eD
Q4XyaDOTRyvavKZVLd2YPUkOAIl8EnxpgkUU343GHchjL5AsuqDXD5OTvs1g20xW7zBNYX0RYc/c
AM5pQE3UKcVe/OqY3al552hSGV93/7bTPAVLRLXIbdKDjFLXAEwx9aE/5n6vVmkldFYvhghoZxhz
y7H7asoJcRDFsC7gmSYYqmrq7JeljLdQYgU1RRs/92yKHEEodRXoYgNZU+nxfBBje3Xs8hN6tWbh
ZNj9vKlxOZus5l9O3wiFvCuY9a74gOHH4oAuULs55k+RVggGf2B+Du1oZCsIBGqQfsyOX/PZfki4
AFZCLUIrd/cG4DahwXhQzH1UqWRFSMLlQPS7M71euFz5eF0H04UgD2pAD1bv9DXVARlZrYdROZlr
wCbFGwc8ggm+3veQQKV6jG5N6051SEDpTPzecMP/mX3+ul8jvK580nZoDFbDWh8YqF0DVZX9sEZk
ToJwHw/heax9XBWU0FOV0lVZdrW9g88gZ9yryWMFac/ugGqa8nPggvy5xWjlWyyI08S17WkR74/W
oLL+TI0MIj5d6ATR3VUbbSZtrX5Z333t4v6mKPhunaK6VwuoUVdOBGZUO4HReRn7JOJ1oT6gxyGd
asElxStVNfQgRNxcQ6/U8LTXH37RmKGgGlBGUQmX7xGLrdRSAwz1R19E/QeE/4r56/89SQPRHsOE
cny4d16m4x0vLCmlgT3mHc+1U7k6UyRbo0KbJhtKbnmhr67UB/hfEmlcCaRdh676ga9uYjohf2i/
uah9y+EblVojKyc265fsjKFZCCv2NT6cnE+/NNf0IWZsDX714CcN2rt5OQaNtfxErf12ttIwMjMC
FrPa5wsR7+Tf0WDawHMOGDEzvQ7ZCxrlSmIPAB5WXIqbUZ1SLpnowZfrJOYsgwq6cj807naB9hTW
Iv4887uPUfWSObBNItieAX2chVYd39G279baI28JncRwY2sqvDAaGYqRtFHEfK76lj/Eaufh+Kuu
kFZQcnKCM8Yz5rNWLYBJk7iXasJhgZLIfkrr/kjLRY5JaEDLKcUZ8OpZ2fRJFwW6B3sHOnedzTPj
gY4FPle5lQMJIJ3ll+L43SOVLBxrrKemd7V5HiIHwjd4Hx1Utmw/o6mM2ml83icLSmK5fGiOA/cK
a8Fa8KOe8fPA5RSiwrGWsvbsfLRuo90XCtRxdZAn05VHHBY/8m+1tHaSt1rRy/N4sDo8XpLyJlYk
kGnGSHjghat+HySC16xZGTACc0g581sRiEx7jxn2Vcx/ERFIh3ceAANN5gEwdyNVtq4PAQQEv7gI
jTWFHCaNTrZfq+WMVuQo5an1YPHsAVllqV+QHLzJunhOq8on7guYv9WLIGwiJKKFNrHPqdxNL/lX
Rs1wJGgayQXba9ZkExlGP0qw2BmYwXr5rzk9nzCBa63ewIw7dy++UtKazs6a9b828QQR/7ZeNaSM
Ed/TNcKKEWQdGVBIvQEffLWGZKV7T2RPztJc9+mx69RUgZGdv9extwSJXAGcFjfKiKVwvGmLgJxa
HjW3VA4w2nmyRDSBZF8UBNdX1sNdrdgxeRQ/Yn9p6xmw5I1XLeznEOoPp6rEsPEIlY0m87+Gie0y
aq/kPN/3DQOiSUdq+dNBRcvqaaLHPZyrTFs5Gvo04HmEjIb0ur1IR6k3w2GSxX0asvSr+q+zNqdO
YO5uKsjsL6L0mbH0UgYPKEiDCDBfNXJizONIhUg1mAqTfR+K1NnVCvlrcWH8D5qGnK8ajulLTeFj
aH58nFochcvQCuuFpdw1THvry27MhHEYUUrpxs4MflTnFcNXVX8qWxkirMoF17U4FloJ2fiZcOVE
xX72d9re0O8NCyXUDNszKtkDMwMCRSP9lvRrI9IG9KEJYqvsaa6GU0gZmZQHn5swgO0fBmKRQ3Bi
6cEjqlESDHUJTaWb20KRYaheyIXzQtth9Vvx/rYMHCFEAmP+u/g81q3ziKsIRgiFJ0WLZZ9nk5bq
rlIYDXjRDB8pdGrNFciCiiaLuPo4ZfRUTdYxR6lBkCe6CQhb1O665k+2fFi1sEHw9H0BxtF9U81y
g1JOGSeqszd2hKTVHF5BPQ5Zl5NFuOhEh8/PTzU0JDmKhvs321I4/nNHV7eWWku6X0vQbqYbHsvY
+dOCjPu6liWroL7oY4qflo2hrv6fn+m+jkWhLQvwDBhIXrrZpffE4CejXHWzGl5kA0K9MxMIqdSC
9EIiBfO5erxw9vk6WVSC4TvtyoCy3uduk4MSJ5Mv7s2S8Ng8ZvJtM+dMsaQCg+/80WIlh9C2MhVV
be97G+B4KIJ+6lrTe15oo/DADYdhKMlQWDK9D1oUkVE/VJXUTQdNpFzg2y3a96QKpMmSmQJt5Af0
Lm94+3/I/sRrxVHDQooN/sKSAt+5aD7wW62KBQFpAotrLqZ9bfOTUuAbzpPPsI1OP7VU1PdXy1Xx
t1TA0Vk5Pe+vhO/+9/wx61sTmUZTiVmHE7r7T4FzE7MQG9XeYtoIq1CJwAbA5mUBvhSkKDCGB37v
+QTu0rQuz8jUzNlDZVRkAALBFaK8tSut2DpxJni8JIYZenFkoqV7S0gifdA3T4ty5NJasoqhKA97
R/tcpeSUZZjzNzchLQqpbbKhTBGnhUU33QujJIoilY6MrlCTo9JQdX2hs87yx/vtQfI3TRU+U3i3
eb0lidk6NysqOFi6kXZfVv9GpWe/7T8SmpSnoFH+IL3N8J8/RWluMvla69mruoaBU25OF3rAfq+l
ISmVMGC5KPoTKBpPYlHP3OTSoe/yzNXR2Iwxp/qP7Zyhvau5OlciaaT7bXanGqVq0t/7wxqlrbLK
H7fbPJXn0hoGV1nHSyajQdscPVk2asiPuifSTkPEmscMd0lfpr1ah4Xs4sPeyQk/+sXMx855Zgbh
76cRiWfgFMKX1uyIioFuZJfPNNxcj1hZo9loniwXWUReDfKYaGDgZvdJdQ/mJQ7eNkV7fM42nbc7
6tFjIWiHiAvCOXi7OKiy0eL7Lq8u4PAqNJxxAD/SjGAboQsNcKHbmDOBU/8oyDKjK5eTmPL/iJx0
Z/TibzcC3V0HFZhXBwbzwTA+wqQS1vvoSlLq7hKp/fa0xSh9CUUsvtUqHa8gMcZH52Awoei4nZpn
mclV3q3eGRG/X6657RmLTwdJ+iC5cWvlkQs0XwJBFh4s0YwaKpeJsP6gZGG9fkBuoJ6/XtcqOwYG
bfrr3Ng+aaXKRlFDL0YW7tXvaBynPqht0BqVQbxM8IVkXy8s00ek/Uy2p8uudYcuEf1Yf2BKVKB3
kjCS0pjoQY8j6ehNYVO5WXHXuIPWuMA/9pBrftDWVbZh1a0uaGTogAhE/i7NzbPhsUlgqD331zEG
rRenJNnhoQ99slettM1WKgpgVvv21NyLzA27VtC77sSW+UdIkhC/WWKD2a3DSx6OERDW02Ot4z9b
PEl9oLgDbf4wTbO4ZZQeTybgVHk2n+GPMqnexFOTps24eZhintkpwqDFnca13kDkeMLssT9v3sSu
9hGcqe/7h4clxqebJKPOJLTv2uFCLbG3mPOk9vD8dg0PlLX6Qmi3lVDC/VfcporY33DnWOBZZ7Zh
9JKMIKzqPnCyByIBIHAoogEXHfIipxXTpziEw6dkZByDUApWfoIbuptOIBv8YaRw+mnrYo0W3z3Y
ILaHq268nMzQdq4fo7vrBwy6qefNtbzVTamv3GwCnGi10mOVD4kvQH3e17l0d3cdTRcVfhTRCwgH
WZLKdHbask2lAEcE6OZkUM7gXx5IslGWMQ/MQBghSOXSX245l9vsZLrsspmMDk7TgiM0oEQn1qQ4
ZruA2gUDkmT02+PGfIMuJZKIH+7tFWaCAOE2AKPHVH1LLsexmduiLzetpb+UURVJWFeBWq4JVInB
bXivf8Wm0DzoPhLTM20NznRqfOsRyNeuSPv8E0tvFIqyybDlMKcRGkd73cOwC2QbzMnsq6SUfPsW
BxJZtoxOgPmvFxhIxpfPa4BS+LVUCPMsH5n00jHcn88hFj5YBaCex1v2bSio8HulF0BgmWUtvqF1
iS5/FaoVndRaZVDHVlTdPi6+gCsWGU4Q9gxwbywf9b2n4gCPhHfWh7HgO2zj3+JeKEujlf84Nerd
C7G8BWvAsNQvIjWz+tur+07ORY4Ue4rmMP0OK4PE6yRXqqlHcUCRdTZ1nKZ+L29y87eg0us4RL9K
EO4GBsx9YDDAi/NaA+KHaxVn4JLAJPpPSNf+KcuKFPU681CrCITu8qsalghM24prHxjFVocpktc5
dOoHqQcPM1ZWhjiUAGscjN4elY/gQt0IP+XwVdoDsp0KCIU0vzfy90+LXLKCzHaRI6p4HgKSqhaB
bBk3vOStIEwqDtj8WUG4HF51fwqBI57b3ptP65phzHAqRKwq/s0tF71h1/wBmsKyPoAEJQdotfgi
dE7o7FR2DGQLxJb+nwPwHUe11GEB73D4tLMJvjgPsN3rlDZNv9mJeHfeQ4Y/yDmZc44gwsiQ+AT8
i3GPHJrlz1R4Vt4gGtiL58QirsBmYPFjkOGNmyLfzvJlEYUMQQaIkp+j1TA0QMQHVIyiYUHOdew8
hV9Z9htD7mFVMLNidNecWbnjpqOCjcNW66K8XTBb3W63G6AnMfISnzy9CJALgIoPNmChf68PWcoQ
4BMQ8bgqqIp9wUla/016aTgooShVWwfABaQYdCGsRaMe5sD1jbjdXQrrtqE6A/S5CsmpSZ+BOWA3
twXOJOHwGCuWML8QoAow+fDp5yjht5X2u29V8A187Gtc+mWTzl3Wo35vdrxGq1Ssn4H7PCbogKdp
Q7M9JCHuzyq2VL66VSdBUNfn3aMKRcnY2yp9WImTdIGBMZ9Oajb/Xsp4c050VIyw+q349gGdJvPQ
2aSKcKJpdMtBpwJAXU3UebT5iuHqkoGXPXr7d4Omy/cWrPTFxE0Cfp0hp7oTOFFNybb8r7T3GF3f
7zSGcl5k+1DtY5PawDXdXl1O5sLmlqihdomkUewkugno3M3HSDivMWKGMKkxuX6YZwZdLB3EzXco
rsxlvStTFzcf2x+RAs1DFKvaOjwhCr/j4gA7WjLV7W+QOF6QfGHDIp0Xpwtboff7UG4liy+SI1D7
M+Pp0ZVfA15vAt9PJ4R1fXkb7I/R0yhFdie/TcHw+fqKlNXDcobtGXnwXaxlvGv+uheujK2PTKxM
F4H+tMmpKwpCKeQIvlkLQZvoe50vIJs1I4umaw2WVuADezcbN3azEu83bjSXAQEvz7+1looHh9gQ
HG+M+78Ra35fLC8mgtNFdVcsRfbmWiyBCAotBdy/73BTnRpo2PG9ARiEodkVaGvrQq0dD/+2NUxv
g0E8S9wEa9joKh/rOAsFNl0nCRilgHrSk3mExZKwx40GtnsXrNSU23FxUX6qEzaRlkaj7Os+pTcu
SSe91vS99rHlHRG6wExmUqjpww3oHkMz3sdNKkSUtDWuv1QnSPwhox6dAVNujBecL5V5odEyEBfK
dQQ+ypQ7Z1CZXjBnlCUp1Z9rBENrx+KnZLV732mbmYqynl5d19X3euZK05SNMoK5IoC8zpLpFKvR
24BlLnqWe550Dn/BnMWF9DPjebrq3AM98bHchOmAgihnkJqQtou+vo2vr8hN3SV4Jo8klaU9BhFN
8wI5szWUJv/ThqymLlqhCwdtHr3WPy3v+ixNsITIWdTU9z1Zmf91+hPNSD+uvV+2Nu7/88UBLFxV
Eo4P82z04JDVyu4MVrWG1B3sJqtA06kTcpKQnjd4ropyguETjiPm/D/7+gdhoWW2vuRZc1SwzIUb
VbPvVlOO/+qrQhSkZemDOLAkDBTNSr4ZtUs31FaHA9CvzObSm1rvdLmQZ4Nebd7uiSxOFZTUeqcR
Qss8zyBqZk1kdZxB+INPFHjNqSNE4Oe+OlaDZu97Cn6t+bHN7DEAIs5/XM2l6WEOdQ5Nh8hHcPPy
595wd+4w43w915qyiVE0cToi6Bjlg8B9JYb+FPoAYJIZuo8/PDU1SBkP7IChuujrnAgdsVAFHQJe
LdJJOTc8oCbzK0mw91OMxbiVkqn2MfHKnBIaHAK/ywajjHQwGfpYoojzMrXPFAVs7HdyuwbbdaHR
gbArgj67P8BhzRkU2LeZrhvaoZi6jx6wZ5QOKfMt8+rXTcVmDMJX6ZXpgauCsIOi+TAQzVq9Lr/S
wD5DrtvPCWGAkq1G5cekwCRzE3AdTh4gwYiu3PDibltgUtNEl9+evDpGTCNNrWYifGh0WYxYviXc
tx10kj+o0BYfPNtSgpLHq5c7RXDIloimiWGbEiIlUbK1XqeeXK5GLmvJBBNXQygKi2mYEXZ9+Ijf
ywc+rVa5ia7HSUluy5MtrPYa2dWJdwqF8/xkK3h44IS98JOroPSznUvg217E+NQAa5NfkJ8UphTr
z0Ytl4IXIBumoI070e624ayF/t1MOTy6tkM7JZpBGSOcBZg2smrEzzQBgz+fXSxZBw4MyJAEl7FM
3xxcyI+jb4uER7XBgQ6BcPVvuF52hZAW0Drae7w/iU6PfreMwPf67F7kE98He/Iy3ze7DpoQW/LR
XZpV7AyyYJjwy6AaPxAV8iyKg4Sv4rDiIBf/M1UCNxJvEiDfFn6DW5KyyzDkvwJrxM9WBb9VfxQX
eqCQ06MhEH4R8UYxYY6fi3t1PHzWBT3uGbRCfIbl4GFQfwVSNP9aRA9c/7xPu2SmLCymGXjMlZsH
6fHeqYbb20imylRkpckX/E1TLJ95uoZ2vkyrASE0lW/qfGoxOKwB4MZHFgS9RdHAVHnr8nK1xg4R
D8pUdM6gmK69qoPSd4lCNNu0Crnn7KbWxq0+BlE/RxqglGLafKWH9dioH8wn0vDrZFSrk6SnYCSG
dEoINA6kQ1fpCdmdMrSAWel41+PFHartYOH2ooRgeWreVOX+QL0aegQGdUy7r/cbAVx8If2sIIe0
ceX0ALIk05rWzFzx1nhCRZ2/JAS0HSACkFKIquyQjwzXwkqnuitjyHDdPZYXAu95kZzXLoYi55Tr
a/Y8N4nm6FJRzeKUYNb9AV/mAXe2BYl4f8uX72rTKVDL1yvXsOMu5Az7Qzo8gADWDaRIPiw/si68
A7Q0je00WfwO/4GMArmTgNZyG65O1a5j36vUidwIMSoUHio0xVdIO5v+BzcB0/zzvF6QZWwPHKrO
CakXUo5KEyJglM4+AhuGb2C4qRhVzBxaHV4sr34+Doherm9TyTyP7tBLIiHER25O4XkxYtQ6iw6q
7yu+KSoLhW3N9pv/ezR5MasOZG9tEqe9j2HKF6AD0I1w0VGskkeqgVUowa7oexLlvbd5yCpLCsZR
0BgI8y6X5hkpjmuAJvhIJ8PzZxowA9XZXbrDufy86hXFR9zL/d0dio9NoJ2fN5tGve9nJzPB1h8c
SudbwY2IphHsZWqUaYOeVZIzPfZGpx5zTr4qdDsroTy7tnyl5vxCX76ZJEH7lWKPC2wQHQ3koDm2
/bF09JPsXIphG8NWbZPpyS5PDyo8ZxNaRBWM6gri6PJh+juOhzqXG4gNNIsru0c2J0vfydyDTdbY
d5ihypJ8IwVAk5IaMYEvw3YQ8VRV8Y86NwFYznuzbnjx9GqSxOnoZdx6Wige+GXKvCiJxGTFKWHN
QJqHgPF0xaWXzk2DzFCotBbZJtjZEAzjZ/fPmbYRbMuPZGySRoD3WKZ2Pk/cmEwWMrMdRfUW8vYU
f7+zvXVO5GkEMfpEx0K9ReDAC3Y4FCi7Qkot/575e1qz/79fkFQ/FXpAkVzAmH1e6YE5tVjLHZfj
DWABNF/6eFgzVOuJulN8pz1FTmDo3RXuAkh85rfDFZLJlFGnF72WSmRkFx4I1ypGvvSl1uRIaDai
7d+ReprDuG1RTT0Cfz5eJZZBHPPvxAowD6FdtCvIWgLUklbM0pmv3PSUBm2LOFw8r4EdlXGGoVOQ
7WhCe1DR9Rmh0wKP/oenh5uSIwhqf0jtZqEKOYvoVNHEvc8WAtMqcMFPaUqyRydGhR00LVuKWsGu
+IGaWRkeEUsdaJl5zneZlaBAU6DS+tZ1Cmo17ytxix5VWlzq3c6R5Oo5S5iJV2Wo8bIjLC+0W8wB
QWUUgiMqovSN0NO76UoanV758ge8ejmr56S4IJoAu/0UT5Lc7fZAQpKsCpSm/oGOIF2+7CNf4akE
Ub+zfT9muGPWSipk+pETj9dJ3q7FwUCj81bYxEVDXbQvLf0TsNWRK7ZDC4Ux6yPnhEGHbKUBm40U
/nDF8DCnWm2AvRq1TDgKujQv91nrd2Tsa+fJ42dJBOHpjiSbhh72OBP9Fgu7BZ8nIGf55lUqjZ3t
rGf2BbaqToC5hfpWA28XwQ/rMc4Jhbn0b+XVA7HzqontO4ZLVyrmK0iS8x4PTt/j9d5E3oZXQI/W
vm1bK9FcwZwdRvazd27YjXMVE0P2xSsJmXGQjc49zRBLGn5RnD1U0hf1k5kAPTN0CD77rVQa9HlZ
VrzYC+PvZ5SLzACr55rnPT2JVTN2jSlrpnfUTNjwGfrEz0MViJZNtR0iRIxVsMD0rb/mSLxR1nXx
KJSt0Lbw/mB806LNsvp6vi5KNzPIBcyjc693bf+iCInIr0g01JkwIirhKylrZ0K3MYRPDkvd17gb
I7XiIt/PqzRbK7eUoyJ8PI2x/8L1LHB2Y0moTfWZpEa16KGOPRq50Lhojq+g8F6WpUBm+R+ZX9e/
IQLIX0fPIr9MZECL9tUciTMk4lYFEDgxdNm1PjgjeOiMdUvAIy1sySJSz/08cqmMNLrTDasDqC/w
qoPshhXdmcgmazK5f1FxWFacYCxXfJEmIgYOXIXljQ/2amAWbP4tlVcJuuu9rTrQnCu4yYATQalg
I/dSHghzZXas7Hp+Eqxd/iaiPe4JXvKWPOcZky+sxE7iFKWeR8Wyrh5wGKJAyyFg60xYQoamp3IF
jzljKOoLw/G56qdMkWG/R3EMgeZD0iWz+3/hv112KQsJYZ4Z5iA5LmsdwJVX4GKwk10e7FCV8tz+
IhTG/QLL0EQ1hcKy8YShMlQ2sMtgd0nPiDHzyZcTBDupl7+du/dHGBBlQCNBZOdtcw/4vtXMw6Tb
tqn3Q0SLung5t/wq8HKaKD1vIqCNQVWmeyYXaUff6/4OOnGhHrg2BXnrvjc5VFSSu+HjXDCmHt5W
DL0uE6fe6dtVfmLamgkRJ84s0jE0kKpSvCZkZ3isfAClv/unAu6W2u6KduSH6FUG2QZbVxw4nAhC
ll8vwznKeKVN5zp+SRvrnxAUN/c45W6MkBH8m/kUQRwsdJs2jIG51FC2+cdFw7GaLr3sREbUYngb
qw3SZtZOOOcBgQzKfAtOwB1TczKQU70BF43/HDrGYOqOhSEe/fjoCC8x2aLjgRuQYK/ilr2YTn/I
Hk94GUGz4M96UbGtZ1j3YBMS7O3FqMjiDgfjpUquFGVwUJk+rjHzr6V3kzCo7pkMaK7PiRMXYvNm
6vl32eODqsHX3IiA5z1G4j93+MvQx7nG94xFSDiPbODpfjLfcyz7ILpzSV22NwUT3LuTpswFuy+b
ajSbYz5eQeSEA8PZu1h8MDdnQcsti2XFU2GETy4QRwH4DkDtTAoZgJGiyZvHYSGIRVLuQDV4SNxT
f+8SIf8p4j68S1iq9W5q68OMLKlWAof6BFdJFDPo7g7aN8KIzTZ+bkZ+Cmkys6mqcQ0Jvz6dzdXT
XWwR8lllkDX8UiJVpbsPRAPFGHjwh1DRl7p/ta/8fOXRC95547EVcnartXzUv9sXtZnN3QK3xvZW
42voUrxzG/EfqPvAqOvf/2FhrLe2O3EX6Y8ak5m2NSvohQkAuesXgdQ9VYAC83v5nCV5k6lM2/x0
YM3oXIaDf6h8plR2/UnUvCB9ZzJBRXfOYrnY/xaiGS4krZ5QuU8UQa1V9bcLBXKwXWQc6Hq52AWT
WLMW278rRmHQiA+figKonil4fXC5udl4JM8g/jU/Z7N3EA/BkhtGd4xbeG91P4L3/3p2FTpDHvJq
q1QyX4GglLCThodT86e1q68IJ8tF1Kj1gfrVTamnDR/OgCuWGoAXkhtmcx7ZeYRM7KcG3F1RJk6i
KHtfXlFnoAffZAemyyRbDlVd1aB4omePoEMchSCUHBmnlEDXEcgF03/qqvW5egWwQXIXAmQX9Fd+
2JUwsz60OWg/r9TqCXKPDnSusJ7ILeXcfuMUzJTy52+e5P3hpI3nM3Us/dZv9LYx+3XfWs3hGFh0
r3UXp87VF6qQn56z+zWYqMb4cnPntgrrZvd/R7uJCKbyO+8YLG1PLlJb5kaiBrt1Bx7MeFHDYhU7
YHdbJ3/4NLNN+l0SXlL1rVQIsCtA9vQIbeKfetaPtrybeLhQzVhlnTfMDqVrM18bzaegCMdojZqq
2f03SatkPwYoH23rCy3zmqFEy5IWSXnBJKLBj/Y3Odwe8AHI+eyk69oO6rWiUNeF6b4LsHEGOmGt
99MsvDgw2r6OgfXv85h/GpJBPH3UsKkrJPleNhGaxD7SCvZvEMQ0xT4PQ9ym0vS++R0+A4g4Aprj
MsdPQ9msChLHVi8beCbRUGmkq1Zxrkjpu1vgPm7rleLdkogDN6jnHAYMX1B9WJ4xDounz5LXHAJU
vrGQ8yHP9GgJSdi6mwuvbqFCeQ32B5jmxMwCR6VAQoTN/DfX4vfQmrz/L3rmYu3h0OZCd7tAi3Wd
Vbu/asB/m1Y0CZHKE7R3YcJw8XTiiabKiOgSpq/b4RSW995QvtIOMSRL8otepAeuc9u6mrbd15B2
GeKZqXXBPdHauekPBZjuF7Fec2/91r79HISr4jxWW6ZJ+IJQ30TdCU1B97vLr+KT/73vc9U/24E7
Hf7g5PLciVYVCQEP21Ho9SzfQSPNN4/7r4K9GDnqVtucTbC+VIkGlfWNbZvrMhynO6CJiF/ovWRF
0+9vK6CzT/6fN6ndCIu0dw4Wv5BXBLla0cYldP0Bg12OzKzih6T3MVXbRVvHxCLwoBQknw38fpqq
ABHBoZYnHZDqD0gL20I01a/vmGeS501NmeOTKo2kzM4eEh7BOAb9ve1UbKXrqfd0p/4hQErhfvCn
GqVcLbA9UTmaN8CCbCYCnOx9sCLcS3sLA6VmwwyusKEol4MhxmbLbpdf6VyVPafrxF6Sz/cnKQQ7
wj664cIH87s+A99aoJ1Ko0Mz/woCC+u443bS0iu/xG2Hb1SxtcKiyi7y6rNHwk/NlBvf3WaB7WOf
wypXdY37NLvK0Y2c6APyBReSr4SF3MdWIrngaojMamfiD4oRV0uupU3kqprz7ttKdUxMdq2TRj2H
UEimhFGFmCwz06NKYatn7qynB1XlGPb8O82gML0Fs649otrH6vKM0sZ0i/2aWstKGplKLCwCSd8C
+ZcKFn437bvQu9GPkF11s8E0uKAoCSHKAPdKTn2wI5aJw0Q/j/pLcIjKZyFSiD2J1CLhL+dR0SJK
jvyLla1O2u98gKWd8i/Ge733psxfTKRuIcnSl+omDXyignV7fElCLvTF/xLJ6e2T+BYDZpGfNTqU
1EXI6mDx99od5AFjR1YxQM2jom9VlUfahkLQ0ngj7IE1+HxLscMgMF6ItUlVL4ZYeT4SF+NCXDih
ldRAmBQqxLoWh9OCIQ+roe5yd3OUNFH4Ox4v2ZYl5Ch4jYELmd+h1TGP9NhSKKTM6jRIf/fQ+lJa
IhqUY2TEkvnK8+V2MYtfxtQoVW+FjebPjj+8xIyOeJBt5egz11YAKVYA3lq/hNssos142zbo6PfG
uujlrKHp3+KuMrK/j6CsN3+TxTdIgsicyk/wEUkV60/s15fE1digIPRgOD3WggwpRmRz4WVJLTq1
+vaUEyv0RPEWsDTjJ6YnMHWpCdHwgIAgyWjO8tPxWs0OslrGpaq2Y5c4dkKvon/xEudJeTb9xsag
PADIJfTmuBA0z0SjYeuokPaqN/QMowo3lKMqURYg33FJqLEHwHFtjbh4RjiTEyUvPan042T84fJI
Thkm9c35XR+r0HyZiF7wZag5rQZA4qx8iR6LF3tdwyfW5s0JevMe+Yb2ORRJjgp2HVP0HMnig2xg
KfC9OIXaWEAyNnXBjcBrCnJvJMuGUFynmRJm0DmNnxkgOTssyhrAjcF2sPGCacBm3DChcx8yHfak
Y9BSa8Of7zWuvCooCq3eG/HgRWwuLXilWLgNwtmITqJhIg++1OYZ2AIEQ39pELiqaOml2ZV0njcx
QIwUgmzzobq7Z/E1j9SgKRQsgoxHbTs2avINuGm3e+1W8QVOvl8OUXnUaU1YoEtziy/S65x6TNmn
tJu3JzDESUOEtMdduXRZgyrnNWoRWgSDNPVV1ES2u24Mafm4rEnfBisgB5rWhaRpUZG5VGPobTck
HjBgGutyXp94GeoeHdsGmsmIEPwwnGVbkVdB9Qf22DOGxYee6nNcDq//YZGfeu8q4imUAo2RbFY5
ryNPb4ivkD1+hVv0io3D3ujyN2eACiVqVn5WpC8j7TUU34sGFQ5YvymjW3GWhN1+7ByFWZDGsuFk
OlMeHIITipxA41ssy6BD7CZ6JQ+/MFifHH3k8ycIxyhcNBkSuf/L3T3AtMLU9Xe/TlDW/XIAjiWr
cTw/YZjGbHlJMq7BDAmhNvnwbusotj+jISpdY+OG2ZhP0brWaT5l1e3n3wiIfzqDcH1WRD6QA6Xc
ZyKV3SHOcAARFieLAxrbrkTww1PT4wi2GFEu+XafrQRnXL+7HVkEjYTPg4tE5EXsjXSuQ4f9qwP3
JKRe+v201W0p1rnnAkvFjMUaodCGgOJsBlrMvYmy15+0p2qlkcTm+XyCMU47uNfaROgT4Pc9EZQE
yZ+8aMY2sp3UwJj4ApIaEv+Lm9V+6BWi74zE0hFoREsmHM6vg1FUyYrStMlxvx5s75Gyzrf8DQRD
ScqfEmiK8YzwohiWalmeU9wX3jkw+J7OQTOHleZ5arPiSbRTy80jESBxfy/R92u2VuNnOOPtVjO1
hQJ+gO1gLpu/Nfs8v0BJ9UDy+LrFZrpcVJeP0Q2dz/SzcReAJuD/2cNIpf5sFTn020zdHetUjqkr
dUmoOWIOq7dAch0QirVE8qA+k4a3Rz3V6HWe9UIQDHig6V2FcU4i053GPGtlc2qvO3ip3+C0B+cs
R/Rvc+5xcPZ5EjxfOhyZ2xW6vYgIgZmq5C5LUBuH6HPmREp+wcqB5unFxnjcGwXGav8oOmkTTvso
tY+MnPqJatHMYLxxTQkxQTgxXx3j/5H47Kx3vcRXvfYtztJu3P7AQ+pATzV4V4JUJJucb/ogSXlf
C61hchDDjqXNlej7M7/VIkPpfzYOujTiG+9aDiccA29Mi2TgVywixaPcGvzmmkBZXjvcT/Fnue9C
HneDiSGpMw1nPcVC1UJKjF71Zonu8AyKyXDHkSzjolo90WNeqEiOMYIQVO5mwoUktT+UIvPqoaYe
vJ6lHlZA6EJZe8McrFa0Uo8PXLb8r9RKICIZSG7D5kwfAzCxbNSFAldPUUeZkI5nFIvtFHKW4gyo
6uGYEHOr5yoka7ffsypSRGYal8hwe4jaY2aDzhzeJfPbnC6ErK1FbbYbTYJMfIqmsiQ5zvv+nrZ3
/BkVcQpNMEpESeZVGYkoq98HQKmclSub7uRJrxgnU7BgWxBpwTT1gsVqIx8pUaAgrQF6jdtc0ioU
mhBuZwMtoREXgOU/jsU4VXNzL4wMTpd80seW1wgzb5EIMhkscqPvFude5llK1wIWwnY93XgJNDpt
gWoeJyTqU101AQehtDcJ3P59vEfeufLytasmXvt3c5rjv8APgh43/REenyWmpUfyiGri1qcom7mh
15SlqcwDmEO5K1r5L3bTZAO4Qz/aWgjQE9LLs9iR/G9gDVc1GFwP6ldLkRhp5y4/Se1kh/DH2CUy
X0v/Qf1v7BhfxSTR16QndzeVHsWYRqemG+cRlE+WigjQqF7WyfSQHm36dEYVZeE6n+1sMJGcRPZS
jkYfmf+9ApG7vf587UxXFpszzsCNHNc5usFw7fi/cm/mRWFddWI+Bg+NMT8vE+Auu6mE7auaf7/1
z31g2W/gTvNzO/ytl31VINQTEZ9SceAUQDELx3xobeMBaytAZ5CmKW7taVa+YbDcByh9YFF2kMLs
bPDvUNyZP8SZ2Pe5EGQvHLfLPgIk7xVrCTGjonHzgdMdY/azYcUq+sm8Nih4SycOxwPIPF8KYCss
CXUAx+9JutDEIJKnr9yQYWLODhfOyq3V3n0nSQom4A8e318zc7ZDtLJ5je4QFB8Tvb4eAhOzPwt9
9kVtc72MTQbFZXlqbXi3ptevIWPjjURi6n2Hg24IbJM71fxLLKlCCKAvDKNPBOjLvG/y2NTQgyx+
rH5DaXOJsdkj9nfhgt7p0FJ/j2ZTp1ZkZdx547VWjCYBInHbhh31GOwargEkUvBD06K5dFpGbkRQ
RyHc/ePPpiWd4iA6nYdHqFBtfjNEEY4/7s+pdNW4YuONvX8O8w98DPDQcjV+Vlgm2ebRZNFKrUP7
scsRsn9IoVy7KhBFYxP88rrvBcMe4q5dkOlfcVz+DMOhRPK/V3dU6/tcjZfwfLsqZ++WpTLjEiIC
nLIm8dT+mJb6BANJANusLgLB/h0Wk5Ui8y7RHcZCZPtWyW8eaOQIu4pvcRwwgpePHNY8jmiBcduz
/uLEHaO4Q/mcGROrpmeTYxa5bKcLd3n0OAjt56DTTTLIxn9sZAjcY2FLZ6ZBNXaLmO7R8rQvaHwp
4703k5Ay37UVY8CBIukRFJXjiRKZUX68TgTVBUXg2pwalvRos5z2mOPYeluUvN79zqNILfeReW/M
0sMAjhexPr2vhjMl5gPuipO04ifLGNgQKspvNEXSVlY+yTcwfH04I3NcH4J64W/jxduOthALortl
bnEZeQJgQJVNr1EbPus9Y00kkVFEbOUThgLKwX/MEBKlPcG7NuH0Xl3JqAjRIEhhiYACJ8OqYVlq
jpQV8m4X3Y1Jf1dDbAmQP+N7XzCmcc4IGnM9lUP+PxIR0v2n9VOUtvr8QdXB5G9J5LTWo/b2EO4F
XJISql3OZf/n48HePYSw37u3Tt6G9dFOiJEEDU4H1qz9RqHdYPDueBZVT9VP8tMzRppSPLp5J8/d
0VYa27HECmqJUpsLuPXo57mWC4cCQZvIXoyPYDIhSp+wzQEB5QxeQBWDM3+Hi+caFN1ZqPuL2iCZ
4cjPX3f4HgNUrHQvDkBw5zbzA3FowC/PAQ/9mrLRjZWMjzO+ZAHLPrigEPQa0MLivPevdCA5g/5g
4DB2+acVPtmKFpXTafCSvPdpW6SUGgRcmt3jyrW5P4CxpCL3AXjCWugt47IX3bGQUic8z8vSL/cZ
uWmQWSQc4Ic2qRBHcwNXq+GLpa6n9kjla2byOQSffkp4euaXX/vdkIbrUmwi+lvad4Yg+usum2dK
5Wcr04MyHCdVKWVB+nqvWHs6WXPaGXNzry3SMt+5hlQLe/Hjl606l6NQyyPaD83rME0A8bfGn1jj
M8mp6unTNSIbBzpehutbWRg0Y3wHnVItSR8qvfj+Do2YpHl6ac1cxxNDHfaDfPFfD2/OrQQ6yDST
k+Z0NXpcqOccgYXobFEVnhikm3yRA+eS9o7Pf1sQVUDYgko0BoPd95y5lhmKW0ndMRaNTvbXq7S4
di/zlI2bggy8wTyW/fzbtWymbNz6dQj5I0wYjunRC//qLEt+ilPufI+5By+Bugmaz1FD2+SfdtNZ
RzUSC/rtxvZPxlXJ77mukR2lNC632i528k1F9B6hakC6zWahfxQMZD71vm0AT7Z3B0BToEshioXz
TMllWEMGh+XYdX81M4PFOzYXmBaRAKsIXPSLdK+ofOx4vYYeDbSblGRvBBlW++inTouFN6dPqK4Z
VozUBQeV0zl4fw4kIjUTptRhwZYaLbCYLjZYj3LX0fAJ90l15wgBMf3MmEvng/OyOFcsP09ai4qQ
1YXiUKXcblFuI5Qfka1R6QZ0J7iM1nhrxHFT9aauSopsm0acrgWiepmn5u4+uuyXvW9EIFm2vghX
R4ufL6Wf4dDvQsVcNVPFPpdrDuMHOal3aIKFpIUA5fJyq2vz0MIfZ4JgaJqFjD+tiAWs+ICf24T3
nxpLm9ZtPQpjsSkb8nwcrA+w/0R5Dg1Gkvhp8PIR27pW22m+1VHCfxO9Q8nAlLrirSWtdYvlL5ka
zZtMmurRPjZZGsdnosopKhvyJhTaWYKWSIzoyQWQ1unEOjZ155Msoz5a1wbgKUB9qbIjIk8slogU
GNpW98mxn18lNhrB2aQZfMjFsvygkMmYWBMa0UqRE6eXVIx0sZGFD/dorXOFvKOIKbpmI12hJU3L
Nvl8+YHcJMKw4Nef7VBU4OiFe1iUGfFjW+ri8/0y4UpO/n3qrISV8QpQwsUcrQykc+RVtFvAxoMe
k7S8Il/AOLyVlcEVM7NB7IXgIADWbVy4KE5+zg30/SBiR2dKzg6ZOKYjJCzJ2479Zf6YCm14hK37
egdPv4QzRRBHyT531oSYjnLhk0chLq2VFzLxXnmdxTclUrIP8wArM7pEcv/BQsUOy/zrJEGEmOTc
m0Tw6tz4M1/wCeQgrCRuxO9RB4HFTcajgLUSA1oBZrPmHGT/N8Wa86khWoMWetmwD+yalXIYRuSx
E9SbMut9cqbo1fCDIXuqk9rHhFrjcZ0VPhJTdHVha/BZ+IxcN4yULzB23MDYNGc9C2GdaCfHbhKx
uuNVVV+0DH1cj38I6/HwKQpOHXjewc+gcs8HwgsOgIyUqkbKrGxAgI9lM1KBDXmp6ftG2yPi3GBL
i6KtleXCQXyiRXfuL0nPpgCVXJCwdamJtPprVwgo//TxwsF2Kz+ENsSu+IcwtICS9hcje7YbSEdI
mGzQpwqqS8mrQvErm/vbEjrqmjuRJlgV6FdCUFy2S+So01XyEL5ADXTbaG1kGnP97NRLkDAalWik
sKaw29/oxm/dpVzYIpcMcARWCt2FhzqDj713Jk01z043yu7pw2oJUx0GjlHgcTSNnOoOtYGWbodJ
58+OVl2NuykfVMHFPYsJwcig9txDgByHVR+HVNATp13Au4rjFLrptvwXJXGZyg4jCHaPb+rOgNo6
9yZfitlFxbg55oNaUzTJG0oYDt+UGb91aA8HQQfPzTvYJ4ieP3DKrN2cwO/7JPZJclkFROdHfq1e
yNwTXTBT4YLb4O6TlPW3kumnmVYZv51pgyDG06BMWAECQfXsbkwS0rCG8BxrzYLNwcfoKCnCSrfN
Mc4dnR8magN+G3n+nLu70uc9zCqCGJirAB1dFLAU6aZZE2mrngj75e+lFZZvnWNcxFIQg2nbAzFN
x4uiXVCk0ZUOnquWi38g8VQPVPN6ukDtsMrIAXckoYg2zFf+IY5phTEnk6SKkuwtxY3+SZHnYTla
3iCcZNzMo5bQ+f+iOg7BVj1aKxSMZWbDBlWoRwIhTzwODrS3R3z41z8F63gZ2xVoKSyz52IC0yR2
EgKOB6Du4TiN9RpWfrrKhMnehfOM3u1KsI8eVXm46FWQ1B8s0ZK8urQymqlVgGl3Ox3Ja6RTbUq4
ErX6EXFrF9O//q8ghj3V2s/i8ezSMXC60CCtGv/TDcmbvNq8ozB+fk8wpo3cYj6lbhQAVzr7cqZm
BNvbbXkwmjQ4YmLHza4vj7m79ZcOZhIyoZJczuMexIFDH58R3vMy5I45eggA6PyL992UGngGfzQ6
cxgNNyy2tfcxs+kbEEglInmv+4Cy4Xh0+hcJKyPkd9h19ueA3kTu1vjS8nDFhirX/QTQ4LYWgTaz
XphtbIKnELGKIquCQEWsZL2Bnqqn6KAvjRmfVE0r1NvjRv65Kv9qwqTNhl3tQpbwTviYL7kGT4cY
vd3EPTbwk+1bh2ujY8j5/9lJJ41rAOU5qTUFAUejdzF1N1uCN64CZjKrdaQH1HDJQ5KdktdjEfjS
KayDaxwvdZbktlV8WmlgoBFBLCqawG5HpWp5scTg4jxgfSYQVUhadTTGyzh9QyPIjSx7Q7zf8aHw
U4JhdkURmjDLGbZ+f531A637Ve5jLys6eLBIrry8WWlkenQmB4Erf5jCv9jsInNHWyznASxpZL9T
OJNk0xgN1w6XLlUdWIG3+1bl8quq58DJ2A0iE5jb/iOfECJOC5WeKZgYDjEMnBMahYKJReWWb+Fh
P94ButrXVyKYVY6cR74Z63WkPJl3BQMYUnTqyYEUm3POyftbk5ZaZu7ST4Wo4JbXOZj7njBuGexa
5+CvxlBSm8RoQ2/5ppF2i1mGjGOIwAYOi3mjObeHE645KEqQaxDZPn3/ZBHX69f9rx6hW4s8CP87
kljK0tkKbi0sJ9DyhfMHP/2hzVKBKhksSLCLi8fkqAcmvo6OUdwTBvhJhTdyYUTlLb2xIvz1MSrY
Yq5V4kUumM2u3sESWiShNUthgDGLpzK/ZrosMGsSRmXFRKDQtEtUD/1gcwdMdO+EkzP/WevnngKq
kRJ55oR1sImJQmHdPzPU61M6svODl19R5EH2+MwVDscC3NtTz/MyqfJgkv8rC8KW3T9QP7EwaamI
NZdHtbEzgo5Xz9l+c89jg/fCs8yEFd83mvZ2I8rIEIvdfRp/TH8xVvGgvRQc+9JLwVlywXS5hMfj
hL4hdzP67DK1aIBbVs68o08ZYJ/ZWIdUGEpUWVyoKq0XBO2Ca43TVTrinbU079lZyQZAX9vIdF3F
35WctX/SzrSGzZTPAI0GLtCuKDsYOrxuFV3aCpl6nuVhnBZQ4X23QtRutXjSEgm/f9VFmsrviFwQ
IEYTT16211ihRNUqFK2qsbqeyzU4b2gTu8pNoWbzWxCnkFF30qJGqbHDAdVwGTqRuhX009V8BmJI
znpPHamVZ2G0nLlIN7qkOr0xHzXEujc1ULAxQ7ay2YTHREPwOEAsHXz3r7QmYsLbP4PW+/wJA5MH
flU5FZB7SNkRpmkDYT65E78Hqyzg6vcmenweTLHdfGFdUPbcE++Fk/3XH6MsiwrrOqFesjOTdAjt
BTEZsxKbZsvk3LMW2Jqaki1eN6M9GfeqbzF+pmBd9Qo31vWQn+HXqy6BG0Q0Z/yu8PGGNU/mV5Kn
nE11VlPPvMRB31vtzWJWVPuFkkcAIEv9V4QUQbCn1bpvXyZZt7tHRuKTkNkZdwmgiWcFlu+pQzkV
64LaXRSsib6lIeAVxHMgdNXOhXKPGv9kdQoMLq8+9yHixLv/drbf0Sf/ICX+iNSglogYqy4zCzNA
HB3HQqpw2/1YTYQaiaUkV0R/wIe/+r2k6LjO9+NlU8AiFPar57SITflpIQQmSHDl0wppCwjsFyg9
aUWHsXm8kjzUJsIGXyjetu7PPG3MsG4QGusJZvAi5K0Iioc8WeV+Av8bEzZji5VFm/Yu+4UIRsqB
qxHVyl6BeiFex2rx2EF8doyDROATHiXL7cYZ2LNSvgZ26owWG/r5nH0R70ZdMRcBaGe4poKS2GsS
zzMaXaZ6v8wuwE1yg2pMAOMEYOOpNdss7MCmvRFMHFY3ndNpUrhSpZBDj0bcuLt1oaZJiEobE/+3
wCq7R1DApN01+gp2b/W/CaTBPDgYIMd8sR+G6pNCnMRMj+HdIgolzIshSccqd701bfz7ZsEoyzcO
lQ1XqHD9U/jsIELWP5ODJXAbKBbh25WeFzpKoESheRFuGie9aFCftXpsh1HfCIyo0op5tNUa2xDs
84xFcHav3y1xDOSDM/77mm/3AD+Vq2JEQ90GjgVA1oPUK6EsL2GP3cefCFhAYmkwnhaRodC/pSKB
WhjcAgMIqLbUJ1lSUoWDKkKk6+qo+ciPCCBdZKPMf3c1kbPllgh4m1U1eAlkQNNVWrAIacZTpYDO
gEE3qmrObJJrPOxDJX62ly12s0zVZkeuAEiPEiKOKszkUvWLCnfWu+ebCbuxIx9+O2LDwDoUrUSB
79jvIPuRrxeuBoheDgtx4DW0sGxXBtwEVf+INimxx3wAsoNaAmrbFthBf4IdSVzmGELf8+v3UsPJ
l8xLI4gDXy0P2VhPVOl0a/Hvf7tzspt+s4RBi4zdnVjiCwW0g6Q0hQwGGdI8EyMsgBEnDoN6YeS8
yOqhhmHZhsG+zxpgWqNtkseQ5VNXcUXCna4Uzhk5j7NMkVYEXgsKWXl0l2XTZsYrR4pvrQ67Z8Ia
qSA/MG4bB3wkanlZ/cPOes3qc8QDi1JQnsxeDsFSZM1ndbaodVJtiMKW4KGG9SXMVBpos9Y57w7k
kPeoiBwczMYesaAUAxoOfmS097B81HTwOSdoA1B4Nty/X41QgFTcjwaBlIqv+6VKfZsEDbs3+WEo
On06gHZbr02VWl/HPpZlmbaVeUUF4RFpLGnHzwLoI9Atk9WHAWL7vfAGLUjJunMJLiW9rSm7CPav
2a7EO36tNJZ2YoWYzWdr9fj1ge0rAKyWmXUAOQDjK3G1fIo1X4OvQcTVddIsFpFZ6VP6D3KGyv27
r52fXKZZnEHv75V4j32Q6ZA2Jj943nHUvsDHOVk7w/HXpSZvkx1+4gu51iEP8KNouN4QgD3oC4jq
pJ7Hj8jerMoheGmx4lcv2tGnV1+dSS/dkMEZJBE9ns0kZmVxrsXX6rXP9FXZYSoNbSjAHEwZ7q4F
8OgFBJ5U9qUCkXIl1/tkV7S68L9LJthkYpqfgMYzsVKvh3w0vZXRAOiTLTOFltB2GQt7LILK+xjC
w0luWwqz2qwqlOPFPM5bdqTQjm5yqnrasblgQjx+tqkFvR3fDw+T00MKO9G1eQheOnVLFT9+hVnt
hMb3cyL6BHvt2s3cCphQF4NIIxDoIDQK2dXinNuHcNC/CxUpJLfn3DZM/uYqjHlZJtgi/KsD3S87
TKozFEXceIQd26feRv508HzhElbPQ49ZFzHHyB/CibTIaHuSErC2KYl8QzYsFWWDqFV4r1AGQmnf
SIsu33XCaL64PUS01W13frhjxHNRQuPJqsFpydskP8RpSritA/L/1DXfKd/u9hd49sSEWle98AEd
BevDbQhFyFa0tWn5cUZ6wxa32wt3ciHMzKdIh+jc3q5lAlqw88FPm7jeloxTImP5KFiqfvVA9imJ
mJg9fVE69H5PYgj1wp3L6SvSylGxS/yAcbmKiyv7yoNOPn84vKPJkTw7b7mPYjyZ5mUnsiAQAksa
uyKokUsDJLFWErX+GMrVrbPkg2ZxnOKMzZrm7aygy1IuZv1eLy3zPRxXbxB30geeSio3y2qPjlgY
Q9ynWjGzn/WfnAY93+cvpkOPTPiUEZ5nsDg8bdflR7/uyxaFXqGnNJt8qLBNSiU5Lv/5sMXuchk6
R8JZbBpYirDUfn8/nAkeWpaURMLE1IOw/+/eqBC1wOrCBe0Kb7n1cu+BSAn9o+iFF7HZihhnGHtN
uiRxIFzBuMq7Yvfd3IE/M3tZdsHvQajkV2r5ayLgy4Q/vLI8no90jrXS7l5dtR/VgGgM0Su5nKe/
mZ7yyEM7Bimrthv5aGgtxkZD+HI4MCnvudeUdzMZn/tjUGV0MjG7cFixa0Og9f88JloLdFpVsxZP
wszqOqdKtyPwGDxbQbYczMoC1hRfCDqN533rv+GgbFhHeZb4NaNzorbd6fIgIQliYMzs8MC4UiaH
Rq1MwrdNGX85/JnjD6qfpdUoc/Q1IiNS/ub4JKxt6JW4kXYo0XkDe31YWQOhJHu3PQH8IZ5XrOB/
Z1Uw8UFhZzCzWJaS1z89ju7qbN1ECce9LjRUzsmDSmb5LkMquNQ1ZZa3eD3bzaSB0K2yV4dEdYj8
mB++rLOrq4hsEos3BQMETRaKFuM8/hcK3HkRQAwZuOscKkiUl2wq2DgYfiDMvLGsV/pUy0nFGJ0J
COC578zkEBPgE1vVqpaT0iyPmMx/19EZ9LgCSVyA+scLR6oo/DOh4ichyH/CR85btlxJKNCq6Ddd
EB+MevW0LYPkEzV/ZcOnjmytvZDAb3gJY8jyNY/LBgqRfW6Skc2vqt+kDraDxtswNyDSUZ3FsaVs
2PWlMs94ylcc4IMjE5NC5yD/6oXkqd20KeN3rPkv6twi5ng1q/EWKjawp+IQXevOY5MjJ/3n/dM5
7oDuieptoAcaQ9IBz1bRWin8T/5AisjkP1xmTIKX9mIPPIFPD4VmvlgCEzS+ZzjLXLPMW5OtzZ7C
L699mhXK1R9Fme8yLuYPRlOjIqBQ2VLSE/k0koLaKrZK+xY0SfTZWs/1wQGoFftqfGitoDWpUtd4
WtvcTKBzqwek5cMpx2/JR/aDd5nYn0+fkmnwApzcFCUFN9exECwkEU8YLUq0Bm3y9mWtASFpJGvU
xvQWyufgZRwE6mjrkhd9KWAukjW15SwoiApXM5l44PYZGZmBCx6gjf2W8twA9AYrdaDee/q5FPxi
KN1g23QGTypdpTXWEr49j4CbNpyODmv7iKJmZgtiAJ04g0dyLKeYwOW9YGQIVr3FiZo1J9HuOyku
wxuN+MCMI5eo53yanEM06QfseXNXVnrmJZrAYPy5BkCDQFV82/JcqSvwxp2MS5JKUfetgr90HeBi
OOfdjpbbcBZRGoi1JWDAjqpG0P+4IKCtMkZtN/rF56XRS9UJj2OvSSPmYKBHibTa/HrZkj5D9Doc
R7yd0Gh47pHIeEfklVuBElAZSSUAEcXir6xQx/ZJdITWSsCXTRL0mClpP5IVi0YfyKkEIXRRv9t/
gF4Jsr9lXTRu4fx2YOMIbS4zfXi7V0rRFqxqvLNFgfQccefC8tKFVqnwzBm2bZEMqijdEBxF+lm3
KJPMwiReR1zidLZouqnBWvhvy25YHwWOJyVSOven+t4mja5oQeILVWwgkmhWZzgqhnQ7ZXrBKzeJ
nls9HR2PDeDXk3cIksrp5/Ei/dlyvqdRCJ8ys+r+87mMmRNWuYlZK98vewlNY0AX7qXep7pt//5/
d5C0dT51ITeREegXJ8nzUJomRehdI8dThP01Hgj8dUAY3/wV29tYqKlhO8QgK2Z9yNUNZm4KtgPi
nf6cZy0F+j/chqI61vrBBLBHk6hiCiEDIZFVMib01ctACmtOgeQjkkFH4H/nK48cx+VKs4rqPv/j
8GytsOIzNXi1jspwDDcV8r28+xVGjJGyBRHjE0pBS0gQWJ1XHl0rh8Vubz/0LsX/stXACxC1skW+
rX2WzuzLtpLNtk2YAeUcdxcxXSEfIu0mO+tW1C1YPPzGdRQOgthPrhVdHhwLxpVnj15SOnIrrfUX
dInp7oSHVpQLy3+HxAzPHnp97BYReAU9q+kR/SLjUyr1O5bR9hrTrDkSJoEwN8U0HuISY0GS4Ohw
Y6TZR1dey+fsjyhXGm3J/jtCEelcjVJqKTomn25MgpFfrXisvOF7AQ0GzWswAAcO7oJo8J5iTYfh
vQc6fuW12h4eIiW/NNglm4aH5jR9uk0JzY8kVWanqurz1F8vDuJ/+LQ9TxbDXOx7cgY8GPk/P8C0
rPkIlPqAmZ6a123cpxXuYawfR7nuJO6z6fFqK0rTtXMJB+efi7NUg851A+HX7lvAL5LPELMJtezD
RxELGUCxsqYrPRUzHxc5k+OMeMOvppO4FIUMdDF60lH8sCe0otV/WOS93ZU4OuOtabQvkcQ6tsJO
4RF0gRG8WBnAertoBSWCqRF+WcG7ZZFTWbIoMm/0lwgZ+35oGp5iBBNcogW1T+gjnADL5xq7w9eb
R+EPSK4/AfbWWCkHV8m5mf4K1K4erqntOtr+Mm9LfGoKc2RS8v1FZ/V2I41gwAmcSmyEns+R/iSD
BAA74d8TqNO8KrV+nmhhCo6unJ0ha0rNYL5+KLQZOoGdB3lKAI3dbSftxBFH8swWgCs4Uk8GHzSs
68xMYcxuXg2J7n6NQvg80tHc8aWRSBSC6XqB0YnlJjERlBTC0pBBEE+VqDR2MylnGukL11O+/mB2
jLDNNzaf5EsN/iW/w2SatvKig2ZKtEL35D92JtbpYTcr4Pcl7d7Yy4tyCaUKgPTszU/Tnu8PpaZJ
rO373rX53guX7EvX8jmgG7ZcWiYIsI/I8cNKorc7/+PZa2n0t/VlBuhPKEoHNbh9t54ikct/BOWI
3Ay3X5X/DfguK8Js2QQ4spLHw5jlz0LpJOICa3hco6hsq2h2vfhTbSV4MGrkWvdIPAlmfd79WU9+
G8ew97Yb9kFd9AuOj+ojAw63+8P6PszWAdKSLc4bYUgfnVWz9BdbWuB7ji6GtSFRm/A/EGqfjR6A
v+A125dfGzesfCjVs6j2v9e+AUc9teDIs2pCs2GwOJkrPE2asNMU9dFwTkWqnKoQ1wxf+AywpRJV
wUelUIIX4bqqLykgL8vPN8/CbUTD6l11ZJ6A/4XOlkrIWdIca9/nfJBbs2xA3zp8e/hb82KaqMGG
cZSPN/BBKmWuZEH5r2aYEXiHAM2rhYzTYvJJ435MpcfNUMacjPm3lxZvdsaeoLl7/1GbfL0eVpao
m2P7zzdLo8KrbLbqJwZfLatTUZA2HhsplClmp2Sl2kBhx+BHDqXBWir26qTghN/f0ZVpw9BQEsgV
is9fdywgztLX1mFGoQbnjuSkp53u/ktEpdQsA6xL/jIsuoc+YONSkWQ0Sy7IdCjt1ZumGKzMKchW
Vcix4m4mymJyfPSwRkJT6PP/jNHCE9yaa/GDDLp571eG2qkeKSEWv4+lBrrFdCTj/nwzvnJ+vIAx
jjQqkfewkRCS7QA5prcbKlI+iK0H7uSHozqezxeGbRfqNJpl0QdtX8duKzDAvy5OhLm69ykf+QRP
hVQxyg+VmUx57C6gL1Yqxb2WO7Wy4yM84W4DOBCSMS/pvnToK6qd5wmS3v4Ln3NOzSKCopmoOTWu
dXmMSTnBZzD51rsdlCgdkWnnimrF9d+PS4POViLf43ZBQJW9IiDJ9xkj8qlHU/EeSGVUHEnUa33i
g9Mx7BXVYW3t3e91yrV50EgBtmrVwgwKROznWgyFnfpRa8qM42MCH+KXx1tSEyol0NTehXEgUvM6
PcYpsR2ywXhjc+P6jzZdTpArsbFvU8aBTa2KXFtZc0patQMHurr0IEpZeCUhDI389y0YMFCWvpnT
jIagZs9RCYJ8kDd2IIuA6wyNetSqqRvamZ5rMT3VUbDb9XsF14QkVZEbwlIyfhY2x2hI9lsNWzF/
C+LaL84EPDwaqMMAvF+WFoqjcbE5ER8U/1OBgDoE+phivF53WkffUWF00Wv9oZUFwFVbkEOy1KxF
8QoKQbJ9h6IYy0MtV+1yw2gwePvmbB+EUHzTOygOhJQ0Px/n45shu43MsiS62jngGFEJTFKmBoGk
ooCtJODIyEHFtruROwzXwmbc84C2sOvRflVfOvBEp/U+T+UsWuDUibWuXUibqRf7obxR4z37EJAx
5b/NVUVzs5wOd9qZtSx2cZHgRL074MgxWUIs0Y7HgKGzisMx5DQA/NiwqN4CeUNqmAhU4vcNy7aC
NfPem1BW5OiwdvEOxu1paNCQ0EkRhrq8ummcCF67Bfhrq1x48LVDqGzoHEprraTE/BnUmnOQYnV+
UGMJCcJR0EvlqDj2350cbdbnU/asaBNq+t8QvSDOHFlPrjKRS0bQZYm9g1PLpV7sv4ZyzTGznnQs
cQlQqyj4Z69XLYpNB0BxGXwMLDnuKn1fYatxgt6Ar1igIrppk7BRkAO3Xk0xwqD7n6YBfzdq4iux
qXQg1ycs7mWpaRGqmyWQ9m/Io/jT1Bls/v2O2jkQauqTa4+PsTE9T6KJd//hhNvAXLa2fV5Xmyer
nuuBL5Nvbn0JYr5xxlAPf4ac6gixquBFWbsuOwiY3zBPIA9vFOREsB7xWncWmMdX2dXjvVqX1ylJ
FKHZYoz79778qhyE0p+G8umJgDM8B5shyEqDJVKF3pZiIwNKb2QjLR3qv2/pfvl1lMOlBCWs8gEo
sWehjUhzVRQyamzIrZuNCP8asbxVEYTaZjxvxVH3x/PJk9SS1JoWS3PYupijyGCXurAb9Z2K3hv5
6ifGC4RrZZ2q+EKVLe8Hj1sMYXveGt2Qh1V+uqOqpCDH5Ezbg4dQcLvS7fJ5sW2hFHP7/hd2Lb5G
6FJ2Dlr1xbgKIMQZadh4zpAx/Xs91/xkodvoO9Vj+vs9LYoCXOBHv8YEeCDisYTT6wStWkA6nbpj
Vm1W2kWXb+gKkfPNrCIHhGV2eWumSZTR53mU1bBoaAYSl0W8Pm0zDxd5Ssl0r3Xf/mjxDlpPXMOe
vYiufDTRfUE2/D4hOVfZvMw5pP/1QpyPeSyPd5ipWb4O6PO2bWcMIpU/cOgwrGOytJMq0JlgvTwT
AwXgfMNT4AY7c2tGuXhtb4p391C/8yckHVcFstDPAltKhZY8fY48dkWMYIlTtjK/hAA9qSurwD63
ud4uszTS2GdFRWnw92DnP01+BVfSXQ4AXtC3u1/w3pnRFvMOVLmYCi186csg+IVr7aVay2sqtvPM
TdfELCf7evJrKbYlKngV/3yrjgWogQd6gr71KZEcxChyasHUFYRFQbRuOqZACCyqqJ0Fb9S17gDR
7WlOcQfJ4CFrBmShl8JOu3s7pHKR4QaloyCJ+80kf5v7vbOAR3fspm5X8/0QZnU2nR2EFIXgmLbq
ss6Uz8bnZWYFth15TGe+q2s3KDte7fZutNpPFqHgPy+8UOzDm8jJhPoQzqyJmsSwP3okNM+Nsbuu
JSMIs9Ztlxu341q8C0aZy0cAZFlEPOUMIBvqqXr27gZdZD7YyNrcBk2JocgVS1waeW9MuxAnzXeC
6En3zP2cCFU6zTlWQqRL+ShYvlDchfZkA0DLQfG0LsjbSIXx7qzcFwjIWyWG8cyU69VPF7SLgoJp
XEi/+SOYnwU/cJzhEnO2EeQmUM0sq2wqSl6GTFnJTwVzlkfyY1d15ec5y1aRIAFvxNUgkm1kM4xM
uHWKfsc7V44gs5j7qUL/k5SFSHGW//Y9dTLoHMuXfpXL70+j0/J9UiO4yzPeWFn3lGG6qw5VMleO
xhtEg0WejbmH0/cBZI1maWgmC4qrEelAZRruSeSRfVa/D/67+2n5Em6s3TxtypgJpv9nkABVHeSy
b83rSuY6A5KF0X/U0vQVJvv4STcjcSWd9RjJTSlRzr3GN/Xhwk7UJPo6p+7SAB9GN76gPsDtD2Cu
80Enqq5miYTg/lgvBAWU/iqs9NBSjht+f8fv5tBJ68rZFy0akHKb+fIAGNLqVbkCUFTa7ON85gJb
o7bU3UqXSNGD6gFrYXv6pNl7PeJUyWWIYL3YYBOeIagRk81DDuetXhbokOA/Rmw6ZRUuzdzVkuKc
5nXuBGm68ZyGkkxSI3menM3ISzsN/ovlZFmakm4GbUsjDzbXxyxyNaPc37SJ8rllsVW7nE8tBAiE
nApMswyFWIQdxOreAe+KlJKIs4Y3MVqaVePnZ77O2y0Yt0XdEvzaRlLty44TTwTjJpV9zQ4ibyzJ
ZnQ/35ZSeXTHzrrTUjDnDOEqz1xw1mzSOn0FZdtCuNlsbSKa8VDl2gwzgJfeTJETQ/SkOMQgMTc6
lHfI7fsC3oRSwFhsU6XTSUY6eJ0UjrfJ88g+aPO4qu+vxxptkf3vCEXMIVErMLph6x6whJ2cbtCt
MS4NHHGSCxlMVwXRG8MgoG66UE/4Bd4RL2UpiTspNAup2cYQTnZFM8foULkm1SiOrTov8ieXPZYP
82otCrHwaXLIhgAx1MVXumsymKYBrEogmQn6qR8gQtSzkngPQfRTyR7j3UrvLgnoMVR/WaiQLVhn
+2mMONYVYm/mcLDmIKsS9bLQ3ML8J+dJTt0WoCUwF4dZtQwWVfVwfhmUn1QtFOpmM27J2mV7PySH
F5ftCEn9xpR+aQurGf09EKebdSYJ3SNkt98ysSRskKFab/xsSdc3jj4eipk973dgjvg+me2fiO16
LrewtZUvQucbaadIUdGvLeFRMmMpUXd0d9QGyULKDAIXDHdY7TgSzT6s0DeoxFZfrn39f4S7+4Yy
pPtphu2uPKpGhQqyo3Co46qVfNbr9fNlQX+rNozZn4UVVXveaMGvIpmJrrJL/8RQ1oB8vvHq2b5T
bjKcPee1GA7QoEtbZ89c7DADfHc/uthoDZtum7zThhoXhG0lm/aBIBWuBSh40VmC3UymCi4wLwu8
0DyiWpBADvjegQEJoHgNmac99IRlCc0C+zVGkMIWN5P896wIcExrx46/Y/Ka2sd51YXGixmV1wau
IiX8lyTR01HjVl21Y7rhKNG2vuRf8gV1aiu2rGpaDBqz17g1x9OmWYX4aoQbx0p3k7uwuUr0mslr
+3R5V3JqsDDQADTAs1Y6o/o60hdZPLlr51RUNvFrE4YvhGoogesA64u75sDGoRkd0nOHtykqEOgM
YHguok+IXWcAHjvlw9QGtVPbXPzEzErJBts4q+ceqUcba3M/d06ntNRVpZOf0/Y4BVngu6iUbBYq
c5IoQDPaw5BA4AP94ZEORDAzFrZVe8p1q/GVaBNA0r4cCn6B3N0Ao9OGULnp3NooMMMT5NgxktpK
c68eU1xSU8oB0kllErsEFMAxVkSbI0+ZBDQM9M6Z3q8VGmBo/7uYZrxW8X1wchZsuqsysQK8HvAG
RYVqSRETsH5TBgjn0SZr7As1bOpF7rmJ2BGFq6/Gn0OJv+rMYmYlmeQ4McR0VxCyDNNDPcWpMaeP
dDT+UpH08WgFWclt5P+7NKSu3voXgrvis/q697L7ELqB6a5/nB4g/+wH2njlQ50Ufbln7m4aahsy
o+uqR4YOjp4QHFnnR9BhJAW/bavCzPUnl0WZMWnwDNq9q5eVQW76Jhb0GkZFLaBY/ocql1mlzNJU
KdPd/YRE3R37HeTTM6JQfr7g/RrxlwS67JYopZ6oa1Qrp+9F88WIxKzM4ug09o9jedfRCWO+Pkf6
JkEvvaU1fBaARWxat/7D54QkveujIhiIaZLDI5Qq3tOUz82Mf1wSzJGo0BPoj9ghwipDxeUBbYe/
dp7LF0dWMJcSXgaiVn1XNAPMvfeUbyT9JFVzGYkRiKLMFygttss51VRuuvU1eT05KGG8fYTv08JX
inyw3OAf1v6SZluMaWxLCna1SI6htmge2jNBBUTTU2+wYqaEuAB5v5M7P/pLJbwhQgttXtJ+Hggj
O3sYjtBZ/KgMvvn1Q+2X7ppskBrTJjXg+QHC0IMs0iWnDXyuy/cf0grGJ1t38mLDMGTKM6B3nUC0
7zSgLGj+y6qWec//IQ/86EHgdO2PWK87eR67k4WXfOraBaaMFHvIrBGHHvT51xft1zFS3NTZs80h
unSPR/YAm1xXYzleaEPiZCKPziOHhikwDvXGnMkaTBXI0rzVqW9jnWYAd2MZMd1RlRFoQFGuM55x
9SmssuhLMSUGErnBUFfteIxonfIP8HFOe8GT5dsXMZRdGdMVSZEKvZ+sIOt/gyOBUM6E7xD/W1Vh
ophhyK27ImS5BX4TqJllH/EDzohOFDHhq4/it+o0aNKuhxMWa7G86vCw/ssFnZYSrARmBlRfk9/J
Gjj5/0OfD1foULHLQ7baPMLB1zSpdp/rdQ1RWIwAOYy4SRlMZgrbJd6MLJDk9N75/hR8n0oNmp5b
yZXFqggsbF6mLFU8f7dGgJK50qDUFCpKMSZ6Z513ahGujM8AMa6ouglwTY+E2iaP4/bIRiTm2LYG
NJveAFzrAtGecvjtFOJ0JrgmCEjSrvMUGmTOLodvhed4n2lUBfeX+HH6U0KBGOjOdf9ZtsOCjVRM
HBgM7b/VcmlEc7QHy4sTriD3sJhhxhwrTJ9Cq1pb2Xd9Aogzr7pbtwbAr+THETGH+lLy+BA3vAit
ZdD847xmvQoMS8bGmLydYO5ey+U1PnnE6G+T8G9YZiYYw6ajH+6+497V1SPBCc9U/EMQZG2kAQT/
Ey3RtzOZePSyZf3SEIgSQ1Nw05cSwK7sNJWdHKXMlx5epd92v8YS6NrBVxsOY29DwNQVfJnqjOUx
XTN8xLkFfnONUtyu2TM/GGaXtTQprdoMP5VVpox4ZN0uN8N5RgBFSZeMs6asr76okZykA8Tu9VQh
S+Z9h+5Vp9XJz4bsGooW9iruRQSrxHe2qvC0UNEGxBUy0vBRwgeDPYGGN199akBeq9HBppKEIVhl
p0rAt7m15HK/vjQPdhS+vX4Qtryr0Yz3IVJaEsPnn3aS0fX1xyDVE/9Tqamcu0QVoTy3OvJ2gZvG
wgU26e3Q0F2FIk5c23SXEmQN6VCW9Gr7gU3kpUBTOkf8GjigVivjjmsB7cjHSeRWbQoqgQjKh/nF
dA3DFSbWKWUWYF1IOpzcyI2tM8LOp4CMDm8/VvzEKAOC/26uCMxNs0ScwGu3kbLWGpYeEEV4eeBj
Q+dlrwAj4P8k70M8YBA4YjPJYUgFEkG51D6A55C+qsVPoEw2Hzezj/Hw8fxmCukO12x/5bCywXwi
AUkLu3tTDE4OqxsasMeMb0WN72aK7lbKZX1ajIPC9ZiJ6qQTAieqOpe6qKnyx0b+ED9IElj2I4jv
EEo2Q/hEwX1I78AIOjxpSN9RmLh4LdMS99iu3sTE57o6bUe8GefvwhhDyeljxI+C6OVHhXmG74iu
scwAa8uQIX2fi/uXf4/OmWybAXtKdBbIPVHgE9BWLmsQZ9Jib7DOVreWgWP6jp4Txs2yPY/TZUu7
Mlh8Tl6HZW7zxjnMAo/GgsTkbZuB8uKwvR9/Q3C9PfqID6JjPD29OfBF8A/sicWGQ7uiKmKH80Gm
bwBXSPiKiKRGUqgVXYXmNnduC7450nGljt3VVnM37R4qi8lRwMpahkALHP6m8LAr/pJXAztotQH0
TAdU1r37txkXymvpTIo7UJ+7F5w8XkxJ8cu3d1z83UjLVqwvjsBwUr98D36Rg97OurSa2SOaUvPC
MQnuhZxEYV69W+SUbCKdzG+/dCoivEdKBXXn4tfEEMQcvKsXRHl1xPDZalo25UQ28/kaanBswyoz
N8CJts9oXE7ucQ9jd/C4exbn9rHScVCsvT5dhr37xSgPGH4JlQXMLEhL/9p195erMnTUnJ9DuTGd
xZTfrgzFScx2t9zg04e4Fl3TbnvxLWTMrano8fMDF2vEEeEjNETwHtXjFI+97AogFS7hn0citr9Y
0BNNHzaJk/QUZ9tCHC7bJE32E2FyEWs/M8dS5Q/ZcxnRK0YtLjam6A1EUaKf8J77eFRrOU6iAmnX
rqKb44zbu9tdAUCA088nYvOioV/X+wGi8szbLV8VlWFo2TMmbVZJk/lNZ8FagA5bLxLqYUsSw+Sc
FRjHHHbhg3OcfHr1R4OilcBxcrc1q1/NMWwuuS8/gwRe7fslwg3bE059bt8Gob8VG7zm7DnNxjDx
uLQgzJ64I6ONPEumB3WoMM52rKo+FFR8DU/9Ec39ZKoJuGHFDokUPWSt3+CeEtfdwFSdAzoRX1pz
/O6S4yKiJBo5nm4qtcaYjoBCNKzKGhCeU5R0ydwk9bZQ4IdwjYIY1mVxS+1DiUR2l+tHNBK7tpnW
aq1S5U8LMNlWrwUQl/+7cjp2+bQq4VOk88jbVRIC6S8Zwm1fsAREYr/+0CGOzC+lvAsLE2vUxqZQ
RV1zCdBKBmKcB6imDNARFgTSueQmg27iu2WpZFDsn5ejJoBrQeJ4LQUp3EaVw1GGgPYfYIkiGcJ0
YmBd5rpyzquKgHS03PG2RB+vGISfFDGuwj/RPVjRa/1+dVns4/kXDHt/PNfpFRAh4LVRIGkXpAau
h/Dl/1KcgzCKTDAysSwkifDc7bIX34/MaIactKXi+k32G3XOcb3zvtf0qwcerqtNjwsUKeOpBZ01
uAaa+0R4+4/72oVd/xsY8ngNPW+J+x6NdiZ/Gi9SCTUGJ1fZmMbfm60gzZ9GnLrwtXurKGBUvhPq
bQnveG8O0L2hDLOfDiBsv8OMnn4lieftFxBn1bsmB0wnt8vHqVuHSdq/ULWHLwNFPqnh+esWZfXL
F2X9HKWdzJSqg6+6qc7hFZ5G74ztCI2I2Oz9WaIx8u999b8PCf5/0GUMJopBKKLz4qfsSaCdkKf4
7aDydcS+EyhCINAakEgvF078CCUBUkwjRvpdUJxIQ00xOZ8dfXqfmIrqTYIb9kgPD73p2fO8ovlV
ZVUrCFYbcv86LmXgUngsMWCf9fvJBOImZ7YYi7gCxcXPB05JCDpDYQA20v6QLBP56VhEGOq34JlA
4RE8HZ36vMB5bAhHWA/OO6nqr+Y74pVxk9qb58o4yxaDhmjqJpZ4zA4pAhIAfN+Odk4HVDGW+BP1
J2wMR0ve0GJGd+s9lqCFF8oZtoTNHRjfMrKS3DTkZMA/mpI1eFtW061f7mMcYpHmrW0qfy9/Q1hP
O3q/2IqofUwM0eEYzxyMQfSUAT/uhOimsj/+PHNI833fpH+PWc014xVpPXkDUTG+z7xn02xLTfq9
Xhg2G1/9eHw85atT/EToGUjsmLsAnOuiEOPP19FskIGknN8yVtVW2FBPPT5JnSC77UlL5Dz83oh9
0cor85iyrxWzJ8PdEqDqT71Dgg1CX2WCjJBnxAxqTZe1PlpM2ZA/PmdR6rXY67THeEcwdQA12Lal
jRjeFYdcTPbfQsTmjUQ7CnPuNEMS9hXqWVTr4vINTe/Eocr5z76IgGrSIG5FLPOKBfwcmrbiRqyv
2j+b+x0U80ME2hR5DE1YFXU2jF326+QHc6376DquEZAni4pchKnvGe6Q0om6TztYkVp5k9KuRd5I
VfmzI8Y5IpihZZeAt4XL8HCk19DEj9oHCa/ZvHVFwSLzSsZ63VWSjfrwwoZn3Bsq8LV38DsVCqTT
MQeasEYbQf2wILxSj+N7ZljqprKPNZebPUsS61KlbjJXo66TLNs5LB6jVcSTfhqxiAvcUzq+H2Oj
vWzxtc1xHKVk8o6JL+XcpVAGp1Ff9NKlafJChVpkLIJz3ERVcgfJE1dv199mwTjV7WESDP3fq6Di
Mi+3+P4ql92oRTfCon3T2pmmE1j5I/fHelv37hpGVov72H/F7bzmsvY1X4Z+Dc3a5+4pmBMOpS3i
ohEe6vZ6yU7bKmb4xnuv+SQv8GW4uixdZnIC2Ny4/xRI8zjJTO88t5faMekyGE4riSGb9pV9TiPK
pD41wtV7+in4iYjgTHDhzW5S3YUuHxcvVhz4IBiPzGey0UYU+v1R5y+4MCyV4UShN8GEuocP3nI3
FpAvhHmS5elaL+aoSOcB54zr6xS1X86sFkhIEq8AByTo5qs+4EUtb9dFLsRpbk2ZkBSYCrYHUoGR
7PinOOGhBx10xspIDd4PNih9MkJ9iNzRLDKD9MtnYvyeuJyIEzYp7Oi/4kJ9DjmrP+lLuWRv4ldD
mD8li8t4gx7pfyUOe2hXJLLt3sTUd4/dHrIrqO2/bm39jJ0bu2rK9genfbCyMnfgPsKViasbrb4i
2aoqG2ax0pnhhJoBhnX6xxvYUy7XHifgF9J4dJiz15blT4rvG6JWTjQIZjH+dNgQmHHMZm0hKX79
ZIKgmE3evGc35oH7xxVC7KzQceMXE/I6hnmzipY7y72sZGwPdLMOKFCVD6W14MplVsxyWWVeWCKm
QOg7QCvJaC75CT8LoQmZIzYmRWRK23RfSLqOHQOlQjmRjCMsZ/XwwmXAdeL7/VoZgX5hWsX+9ZIb
GZ/SL4nzhkndVjwKd0NB6gurAbKH+YXvA3rmp8vDi+fgshVzDUA7IkK9RemXIJfQ5CBp6GMcLOYF
9Ub+JsJfo0gtuu35JzXhuF3w3sjkY18VPcdNVsPNG1lqqxbzCy2wejIjBd/gJi+yrVJK08pIV0z+
XbuXD9+OYpwXG3VQM132fDqP1DGsBrn2TP/NFVtHa6lPl4kypz6pk6wjO1SKgY2a97CcucZLaQXE
sulP2JrjlysMz6/bMkq//SNRHLS0+nRwIZSZTK123nOhviBjNfHI7E4p9GyspTDeXw5Y5CYQksxV
H0d/hQh+K+Ot89R8gJmi5zYxzQAksN5WdMSM4R9BBhYqCecBt7ErlVVPWWJ/0DYImqpsBsHtE8nY
6nabG81Dsnph7DD+qgZlHgryQJr9sUuKkTWODUq9ZFZRn3m73jwBrV+b7Qqp33oWQ+DSOZ0OpcpS
JkO/56EPTcAI41qf6YyJ0+ZQ4pLAczfUb7mlPoOtlDYQ55UdT5Dm1liecdNa4PE1DQ9yFqcJLViM
hn1Ra+IrmXWr0SLiRvmBxz2ZSUyeC8rcFlsIXU8jDE6sqvi2aHJfPaAs5NMT5OVYLN9BpkKXtoGH
YZOTMv/fFkNdg1K+oa3TWwRrpiyxtmif0I3oBuiLe9lWA6VSVx/ZKEl69l+P4BSZSsrk/gjIkdPJ
Maypl3oS/83BKfMYOIiHMJ0i2cuTkHZw+1gpUMIN5X6vmGlNR/De8BF2DrATaRtG4ut4fRJ4IFEt
FOa4Wd3UHeAXNYski4AZtB+jvvpa4SxwK7vtsKIPAOsyIFuh2Q28H4cpGRm1L5sqqjGW7yQ+qxM3
RH0F9dC6rRLmBOC4xXgPvCuuACGFUMi5o67pfYru8rgrf9hdSOcOh0x9/mnzbW9IkNlAiCmt/Yws
GJSEpIIFItK5bm9cPOoE4fjwrDOkfCQiXA+nFtuWaaQ3UxwyReJ8CJSb9MISeCkZfz53UzIbuCP3
Eici/+dEuxdL42ASA/HqIdfR2WRJRAYHupL11JMtux+IT6YjbudD9ieK3Hd4mDn1dWQXynbdYj2A
LgSIsQIMJsnRwJPQAQqQVoCqco8emsn1dSq3+IsPRRLSl3EtgU/jpfE287ZEWUhwzy3H+T4v9TAZ
rYXWteFIxq1Eik84kfb42ZxkYww0V+qQCdmnP2LS0XNLnBXXnsQapW1S/U24PEUuoPpW6/8Ixlmu
djqKdy6BhcCTn4QQ3+ylWyYnF/dHgUGLqbmQMcwTtrg4WYbn7enyeEfue1pccs9jAQWR7OPapXyB
OPSbagRPjS9+uxqgk8KB9BlDvMumCSBeRzjG3uULJU+Kmrqb5AR66Lm5snq7n9g3gj6xsdyjVxW7
SUkn6CZ4PIbQQe25e83wfKNqG3FB4ak5hwDwVjbVE5LbehN4SOIfm/XMx5tdtE1OV1u7KiEQTqr+
PSQmdYE81mSM6GPRQIl3hcXN/xttnmqngfMnpv4jDkzgKJqpBUfP2Y2LPqeM4uLV8DJB9gOQPNTu
xcRwk6rbFrI7uPr1nwVoB1sCq9k7g0Cf/RprAmKdiNX8SAzoTsL34kdXLWRf7AvomKJhGbmbpNN0
+XaPVSnjhjAHPLkXv/RnfHxlHNVR/NpEGfnZ4/w99RsWYMx8qpqTGqZXtGneccmijcORsbYIbY1p
TcIFhf13B+EiwOXrtR/ptOAmbgdHr/QB873KKAST6cE1FAr9+4fA38YK9QQvjcKNv2F5SxWZDZlP
dzTkOCvyBoSql1qmba0UM8BO2z2InE+Ucl1H6bMIzpkw0gSHAiO1H5llPda+IDZyuB6D8t0CrouU
VviOeYKExEN1Bmew0fE5jjbHAmLGIk55G3ro53adrbcqHrTcXyl1PDqQvEcxvbA5O45zGXaYZJ7E
L1GuDY3M99QLoH//XV55k8KIa7FeZwPyFlg9Za1mH4UDJtgZSKJA8onGRXYb+StL/DLR0k/clzbZ
HjBzWozwytxy+32EN6zqj4nZ5oGglS8gZ8Bkf03hSqmvmh/XhIKYdv0x84bZDAruhRYTimZanh1F
zdPJ2hkouAp8LmjsqLHf31r+UoNhiGOLR7MRsqnYXkyoGPusBeaMNxd++ySmqw1sHO6/LUsTQOlV
9yIZeCifxfdPhQdnrl1qIV5QB2sJqE2L+MO0RrbX5Rif8XrZhr/OlGdOczIbSc9rhIKhvcaTZO0L
gnRpWV8zPJBtbfSAgj8tkRBeuAjnQWHJgNZh/N+D/KGlW3SOItohNc7Za8bTR6qCBsFcN/UpNiQM
eh8Vw2MTDxku/tpokXcYJVsVaRuy9kN7fxLlZgffYgL09M+G8PzB0/u0IyQop8i/MJoil7ZBAhsJ
p+BCbicMA9GeGYm6GV9gZyL2rkoSSMxq04gGbkhlg27wmZFehskYAiQHfoKQpkISm+YAHonIJ+bD
6JTQBchoacWAds0XQCoog2dbgkWqdaLgS6VGsc1cF0/ipbvDXnPzKIwwbPRiob39/Qbqb7fjALZu
oCZ4yMb6qo2f8KJKIjjbnfhfzjDgXVz93046MSKcms031xGDNIMQgTguD5dn5XBzUt8mFONLTpON
OoLCoBHkzjc+SB3Z9SwKtlN+9eMRJ/YYG85WEu3KQmhfkfC3uwP89spg6V6p7rgjT+n1gKESb5Qr
4m82YYTI4em6RIrLL4YdammDxkI848FjGVveMbO3t8yz2Uh+1r36GLSVmYxuJqhlEnoWxOLP+Mfd
F4X5JilcPLknr5kk1HtLqJHwq3SBIssR+Jd1rKuWQQQP5dqqeo2ijGBkPKTqdfrdUaBbiCwMjZum
hkzKclx1PJ2hpoNkA4s5b32tOdfRVcLwPCTYhKckyRHeogOIF6R7fTOpmagrMYjo4gA2GNeP4wpw
qAW5FpSX22epCL7oH0H99FNT3Opw+73XR+Bg6s0oxC7QkL5QmKHFHilXZQfMwtLVFz4wo+ibE7GL
+Unasxikdkrx9IqIGN/Te9d/2hrO4STy0kLKyp22BVkHYWdhVY4Qv26J6P8x9uq50kIhZqcb63h0
VsD527nj4uCJ/hyZwWV/CQRJSKP05So4L/oa8Lzg0maz9zEErCHC+NoMOHG4LgSy4ArPdc26dIVY
Qvi+zt0hxcglh8zf6ktKWB9yr/4FjM9KWOrvLiC47T+R983Wx/10uWbh/MCAh5cm9Wc8BJLX4WpM
TqDY21h5R0B9LhUal/Pt6JlbasN0HVqvye0hXaYLZJVyDj+sMrO1TyjiFvK/dS0Lj+p/kS9TYQ4Y
i9mF/HLtBXw+TILnGzF2EatVAuq3OvnGrVw0Ky2EDTxXrHHgjvOfx3WT5GgfuVL5cMnurrZweJds
eWvpgZLEC5pAcNmgydypZDoc5K6qzj/ynQGjsHKHUi2IUDqZgiq1Xt+EOCN35OhoVT8l+VTo7gBr
HgzUyG0yIomqN5ElyFvvFIdfp9q34Sm6jJBCaVmjGnAYGEZavNCxtdsmB5+4yVK6axLiN9KEdlfc
++Podq43l9sEcgUqcQd+RNWFvi5Mzp6FeYux3Hnk+R/CoVYrkkU/6EC9puXiSkATX4mLEYsJHUKQ
jXT6hOYwZef206LaM44NGfkqfz3YRQO7sUsdm36m7BtxJp5gwNvWwvnCYBto5cCExHdFwGjhSY34
MTwS9ypjPA+6pyAOt/R0eKy5psVjB/V9N0qcvbzVP9yVKKIOpnRX/gxIpkjdOLtYMFhUr255PdGp
w/JFHwOraijhDnxcrFmbjTw5wfrVoWgXGFWnshryzhVnT/YE2L11nI01sohf36fR/5QQ2W0ryOL3
9iYRZ+kdplJM0Mzpn5NIZh+P/0vSAw1b+9sDFmJN0td93ZsOPUaMxgw3F4YF0s67Lv4YDkeXaaW8
nPlQYu6TgUTGxRHaDV7fRCr26HY2tOF+t3lhaDQjvNLm2r3kte7cfhw769a9t9a4PO6pR4KaGBaJ
mEEOriLNqEyCUNYdtlMDHMLSDlFeIwVdZ6xejZl6wyjyGceOoDHxhK2/EnWspa/x4snXQcGXdonw
3ZI9gpqQGKSDLD9mS85Mho6Ia44JTI6nv6phGRQRZqrQvjJ2tRCtSQx2kkJUhz98vwCx7rasLNhJ
Yj4xgbNC0zFf+gdBAIBNT+ih0gnbVSeiKk16S+HnlA6YZQzQhrYxsDe+3JRYHZi6EEjGBOUcDpJl
NBI5+sB6741duFnRdbNU9+KUJ2EDSRvWuQff3I+maSfm4G8nRWHD0rXP0DfbhCa+aKRLo+InCYZy
iLhcd2eMMOsHOeVkLTY0k6597xWrIN2mvCwkpjj4DC0qf4B2y36DO05oB0DqeVIBlbhXRabWJQCw
/8SUSY8nvowlpMvUbEgr3wiVrN21dS90oeDPQ+CwpaMBfwwe0BljGGURqR5XqDPW7HZnlA8W5+dE
zR+/GDPVA/RJzD3Y6RSup7XJYVoJ1vNlnILLukX1VVWyWconF2qBzLS8G7ImQAnOaLZBMWfE+p/c
bp4z8wEhuhFJ3MnmOa80gq8c8KTIjE22Zk6AUHYjiJ1gKSwSkKYm/2X6WVRdpmm+iDVbrq4YUuBs
1lafBEBpCJSje4PVzNyRKRqB8urS4xOL2nCOvEE+13Q8w0eshMvdTD5cHt22rwGAxdOpr1yAOYXB
/8InaHHlM4fQGmW2/oGwPAuVgsih2UEAH6LnaWyp1yLFiuKzWI5Veb2Od1cmMLimlIwtxydFZ1Wn
CcztrzE1PsgIduAmGLbrxjLktko1XsSaeAaUYhbGzY/tcQHgXSUceMKOPAf1xod56tEpcheutVYC
bsQm76nTedUOEIv2nL3UFZ/DSXerLHmpncuFDmm2iaWpxY/L0pJJdZ6QGDRNRe4MMpGq9pLE7ozP
A+o7epBHjHblM6818in84jrghggWf7yf1HjJcMTDKe7ZYiFClDYConVuZXyGTayFARgBrEZN+sio
20DW3qzx2MMaApFnl3GAsjVDTrlw5IL/QN2ZhVvPR1JRczM0uFPqQeaEHJdCJQYYWN+H5AbmYery
XxO2M9yfp0gFr43S50wF6dBaT7usWgmKXSn6Kh/OAK7gHUtLQR4xXCCsfqcKHrhlNnDfqQtaEF6N
Gh6AQxfSRF5Mw/2MN+gj4qE3lNXZm7SJ2Bw9FhpmCgTyX5ub40R4bmQ+8kRvEpgOGhMkk7AYPYHq
60PJEUH6C6a7ofbwFlPtKhLUAYhsVqZWygha23VGo1TGcjlGv7Tj5XbGwlgrhnh7wO0ssvTTsSU9
Y+iqYvS9Y1l+pyn7w+YzvztWMcERcm42qy8lV5c6OIXESb6Umn2v3mQxIN0IEmYV+QRx9Erh0LML
kAb56jvq16j5rkQbDk7hbUt31DIHZxbRtslkcAtXUjzsSzUGb5OB87RPDXyozvFwP4bNWXpi7p8o
nk32E4/x1ekYkujdroqaVmQZjvcOLqDOP0aJSpgyFEzSxlE9Syh8DFfD0AjNoR5llpesb+/XEj2+
+X+IlQcPXzsmJM8z3eb3QwmMDKb1+49S39W3/6Zcv9FPWDG+OJmo/+QwC4c1SIAGf/Chy/wR83Up
K2gjEBO1AHehC9qEpWLLSbY6dEbamWsNRjZHTWNsUc+k9jGJoFXI8718ir59KtghjA4RGq3Pvdqj
Qe8dPsuY6gAwnQ2kLi5x23rbPw8nkYImedVaUn8/2C6N69NvR7PjFS+3kRN8ZFx4aXrBIG/7TT0S
/v9G4GbvJy1qcfnI8T0lUFWI+71qn9uHzXD5+i16buM0KwNA7Drdx41Bo019RPbKBGJCzmMY3V1z
EIuOPPyf3qxkHGKp7x7VA3ukNXMKeObJWnR4bPYDZZT7UU3o8h9XMgcxsQWYJ08WghW8VdzjR1bi
3paKzWeqasNRI0eeacLGC0QQVhImWBanOPdKZAmb2S2bnMPfkZCmdJk0m5uLSTkbMZk6HcQidf5q
KM3oPgLmG8/sNJ6rvTNEB7EWxZO7r45Te6J0yPoa6E9LEzoYkOGsriTP1jA5xlTuS9c7D8WDKfGW
6kCk+EoC8zLh6R1Ek1i08JDpQ9cjmLJ8njtjp28Bm2h5EPwstcWYaG9OIqlz+ih9YnoqLa0LCocB
2tSHQ++f4NNZKgZPsx3j4Q9N/RThsgM1/UF5Z9JXx04a2lAVYguvJnc8FF8x09CcdAISyPuibrmr
E8TKtkWddWtBDDkixlN5irWo+Wqy7ywEWpjhEpk7ABNgJ7/g59iDdWvKCe7wdDfOzjoCKdoWiWeP
1gSIVb6Wnyi/D3kGHJM7xZtJ6tnCVLE12c2gFLYD9yuEZ1tvWMII13euW5+/m8HJW8d2AjoGCgkx
zyxhvq640pUdqgLVW6fDGxyIO+czf3ICW9/mEwLcbEjW4/bbyA1IfbBfkrKiTn2xofhY1q8Xz1lA
JVmxaYWAjf1kRwBMHGTTdELqeRGG73NsUR7rkehI01LSJ7SopAA2mxhJpbr6RAPOnRbSDQAZx4sW
YRzZI0gLCXU/VGaSSr/r/xwBaTnpOgeeVs50tGg61iN/UE4y1Zm/LVABK+4UIqVNX8B5ZoVJVY1V
rDcl9OTKjm2MS8esX8m7biZAe6HWtkSeLQJUrd7AvrYoWpiVQhUV2KCBAReqIMk/NlsPgntwBYwC
sWaBISr2cmVmPYo4CIisK6Cobia9xOUPUJ8g/rzyB9n+S8o08KEp/NcmE3uyZBGwZHBWCAo7xTri
uuv/wy9VXOfhtvaW7XM8r7FUdLVrFJUsV1aCOey/OyvX5FCJnrcYPzXjRZDEzsLblvRvtInBrihu
+jCwN//KiUdWyVlTQ/CkpDYswijcWCNbq0s+LF4bULizQfyfxlSamyL2N5RebPoaOBsiqFbyQmWr
1GA6x9ESglfFh0MyE+B3tMLiOLs0ugR8AoErlEqHOfnqSPOXEc9iyOKPttAYFTApjW22J+sK2L6z
3WjeWTTGzmeI5lfLBONKaFJoIxgiu0GfZm7BPsxhA39w155UhEmu1a2gJHYYCPYgk2Fs+/2tTRBY
OOC80V0eg60BAVC3ZcA/EmuDioG1y5knYIv2HTYD/VaAefJqd1TNL7Ko4/5taZfD7U7SbpkRNJCK
vr/gtmcBo6X9kjjS26NWBI2qJO2K6+O4iWv3S9czQGRhHqfQbnPDhZHgO24MScJ6+94GS5/Hp3c6
L3JowVwaQ2e4SGnCJNN3kot8Cu43ydnrKmMx53hkAtK8xZYqniEcz/MTWVj69CJ/KNdg3KHujV16
lwxWtYYqOHAX4Y5Lc3ItEfg3VcsdIy/SIQ3rnZdVmTTGBBXODUN5FWqRxvNRAiSNEVT1vk+jYhWr
Ru63RzLll4gpm5bdzQQkOTouV9QsnbF5jAADQufnvN2ylqHRfD/z6PoqQCxXovV62pyHXMQNDLHj
pBMmoMSr5STs/y6BC0+KWaFY0B25+5AtwYsZKakVM4exfRgNVY/IbZEcITu95b0I+wf43co+rXja
Sn/V4svwpgVKRg+wQU9+pucYhKGceh8Fnb5Tu5EurXRNNHT5Q818eGXJOC2akgh0b5A8g1xXZ6k0
R9cVBQy5Y/gfzb0cmyM5qaObXz4ra8vteofXtOmfgi67LTmbyOxEaJ63HCOADTt0Xp0fN6Dp23BM
i8UI0dlqHFBdqjh3ioTTCJLUeFuKA5cVapJkCw1xsTnJroX1nJd85qXCYjgfRKctUpkg/H7pzS4H
5PpN+OpnHc/ASq+my91ylXWLt2WZTlJGnJe+JtWgBEU+wKO47uOQb2S2+sPwJYquJUuVgJSj/1Ga
Nmcb1IG4qJi33onDoD0OSCQi+oqTx0ifutQD1CT/WGF+GBZ2DAL1W7XLzvilTJbRT7g0wAYuTyHe
SBxyugb1RQ6eu27evaAUZNbPKU3lZvEVFjUEuNrRhBwpOGP+07BD7waLadiNbBWvzyWN1+7BuMRU
ABoBACk9Nu9gE8Hul7PCwbl94LQFXl3sfcPW1IjiAJDy4Tye3LESJNWA4n7DRIKhGJq30ylGhF2k
w6eZsSstOzsGVaoRVvGjDH9cOBv1G6+DM8hmGftOQnPdRy5oDdk0pIARAYzIi1SIcSYpeoZeDP2j
m/IScybbkNMbYwdV3XhwxSf7//qCF9fTR49fAVKfGAonsC7knb872kFb3H8KSDb/GLo3R+7QgWT+
GPQTRH41P35+0Ab9NzLfuC4ffXQHeaaScrYZ9iirEOoMTQnG/wH1lcjnJRKnfIUTcw1eB78eS/Dy
Dq6UgafdYb7p0/qCEWDN1bYYyIZ9Pt3sl8N41vrJ/aWOTZcIErnSV5SWgRN4+uGfcklCvZcao9s+
4K39Bt36AWc/QtD8I1SSHCrR/aKMHt5qR/TYM+Yh2VvgaZsl2u3iVpa4Q1BhzVczBhhKTADsIy+I
0bLGj8QEdQgUWDX07FSFBL3gUq8o8B3yUqPE2ihe3jgQgZr2KM54u8ezmHv04/xjQI+1Kfgm7mNb
/ti23miZsApP/ZGoB00qNQXHhD4YN5FjCXKB2XWHg81rUK5VwPvMwirEaBFaGpXmS9v3LW/d3TTs
599mg/yaleexBPN2JCIm4NZ7LZPkvsSynGZUSuOEG0Ws36kaeXztxhQqDuDQzhFk2TXSW2Du6Eev
qOrgB1v7VjjKLtSj7PnozzIUi1LrhISitA2ZH5BcobTjEUiK3rjFr8YF52bKvbzcAXrnIJJcL2Yh
cG3V2Tr0wfmLRqpehAUgN0L/HkHi05edy2JYfxQTW8gTPS9l/2QGFiv9+Q3h+FiJgiILnO7wFIZ3
ipKVqQb75IFzR4g+wWj1Ifmb+SCOu1tc9BPW93KYsr+90Q1EH6TyUDUFqJveHWUtE24LJ5eLk+Gu
WmInI59qgJcIIo86nTk/+uaiDX94Jfiyx6fSOpy4IFFfsl94Y3ZsOL6n8ifV9cy7e/OrXMB3sovU
k03asetJ+bX5aYenCTMjOZuDLeqh91TKq6NHl8Md7lXGcsCnwJB3x6rOB3VOyYjwR3zaArFvtw4d
kOLSEPF/2ld/bxP/wqxRk224IsWel9QQRNCzVrxj/FH16YF5nuKpFS30T52co9b40rMROc98LyF+
mNtU8/ea4x2VC9fTGfO2d1q5of9t4IjMuBYK1aIInPP4Ve5otpOzReQP3rF3/7nbG9dSJP0li4f/
10+bMGmzz116dIsQ3Uf5GHLna/Ce+LIvUolmmwCVnLgivjGTjmq0pQuUVIaWq1sxjAZr3Q7PFkw+
snFkM8XfgLZXtfoGHh3NkUl9DOLC7mHplk6U7N0+Qe4YJlfUUWFOOp/EfyB4X6k4+MpLhOqRje4D
8ym+VXLpyqO6Tm4uSkNFJJ9Pu7bJzW1pnpxgDUFDFYHVscZwSjVPI8Na9+5D7A/KGN0+02UblhF7
mkLiDSbNvyO9iKSa/DSdKdYigr1FTlNH5xEu6pK70adI5lzA3NjSk0jEfgg/OOCBEQZLjhFVI0Di
NQ29kcKly1pJQrt1a8D5LBoCr41HBYoHg5Okfb/iOdO99f3ssKLfQJhi1rvtubhxngMioyvMqv0P
h0SEzR+XYCZnRYdmIhcNd2ieuc+4e2TmRoNt2Lyzyzqr8Jv00/m4kRBjgBJrDEiePhVajNz4yWqy
ZNFLF7XydnLXntV3S9EC8mx4P33Fti7vs0JVRYMD2W2yKuCuGqlrxTin68G+uk7Fngu+eKIE1446
M/I/RCoR2NWDwsTWySMmy+SI+jAzlUbc1A2cb94SahR1dETC2sTdR83Tfl64NlkZSVOZacYzEyEn
j7Kr9UmrcGd/g2IrYacX6RqiPUyY1G/ZQWu6tjilKxdndw4bvztMFH4ddm3brC9eh5VDEFcvNS16
tuP++1EZOIJ0nISU2VIhW0vRpaOWE7eRsFV0hRUknJrC9LqnxoV/e5A8pbzODR79iwH5wxP2aJk0
807XiZ+YJQyAXlLZqIohu4XbEFN1jcxTSxtvwvkfuksVtRShILyVErL4QAHpzLOhpGRFHIQnKq1+
ARd+3LJMzrE4hSVGwlWUVOEbnVIALzHYxEKHeaV4vMf+zDqyrH/B3my/SSXli0mLnBvAidBjXMGn
QkZrbRXm7yHd17qdV2w00zlrBwBtQC44ryavTfOuSmqG14LE8JqKZdTnIb/0s1GeKofuvTY4WkGM
RVWeflFJvU4sRRsq7mAgGozyxYpLhSPI6FlVfxIFDF2Y4lFKyFcxmJcEBqcxOqakCpFpZJspdFuX
x6xnMmTZUqYOHOwwHXlqDcKOUlXISZMr68BdJ4U4DtL4lRc6LqljRnzOhUGUyov2jeBkHVV1oni2
jCWlnaQ9x0ora01lABHgj0XAs/+Id965MKOEsjhUifJUzXXOlNQPufwajbsxS21yIN+exu7IxSIg
IUxwjLKfQNBfB6M7q0oVLJd+ZvSA4xFVj4Zn43gaMg3xCC4rdoYvzYJ6WauDpphKybZUJrtf7fnQ
Jp38+IAiNU8zQ2uJ+en3j4/jSmy75tiN7MgcSle6RIM8RRZT0ZKUqd0gpisgEwcZOYJFM+yNzJpq
7+OUjsW9rADbcRIg6EFhPrfm2h1C1l3n/ud4wFCSNKQ1OCe7M7sWvXcVUMfZz1I0c9gFwtn2mj4K
60dveXEAO/dg+LXwRVM82L8nfbGhLhyHPNTpPqM/mA6OYgcLb/LC/v1v2yh6de1GBwMv3LwcJpHn
pL6vwye2MyoTNWimQ5X6dXIp64SGTwGgqKtH0GuFhNHmTxPKc+wQbmr2fRl5qdKYfdRsoL58QSFZ
5+ME/Vnr8o/vMrJhgkgby/33dNt8F4i2VSfDp7uuGUZvOwa96Pm/iL+wOTtXyTDdeCdJ6tXshWey
iT/s4hAKfpA7MBWzWq8zdbjxIZyts2wGxDZvOuWl89q0nMlcO59TQGmNgVdzFTsxPk3lRCmv7HcK
OGUrQO66CxOamDS04XCfpBKOiKPgy1c4N42r0K+hGmPk0dnMGClfeCzValIwaChSA4j4Fiq43uBq
oBXTQ/1GxLAQqEvZYMmZvcXHUjAUQ8g1l+Aw6nE2Z3Sf4tXcTEVLguyCrp6lMu4WcjRaxNtqpRt8
TpG48fnrgkaNk8QHhFPL14Hjoo5uYdf2MfK+pVfAWX2cpLChW/+BKzMSfg6ndYJM3VHldugce/u8
zikDSo6neAGQcC0/kj2KLrYWf4lYgk1uWgj/GN3Hf0DVu10KU4kabmBb5uk/OkjgFUTsQHHl1JF1
UCjx58ChcKsc3vnbScvErwCrHfyhur4RzKHFpPRVKzxYyltRGcyEYUKr6T2F4Y3PdXiLS9HRxXii
lohdOG5jn69410Fj+6Lpw5ncRHeBt1dwOR0NVMlYOnoa4YRHqdL+webzM9+kgAJ12KFpUkLldCZO
6/xSs0A4emc6RyyrrnO7iyJFE+u+x8VbhHacLf/BQSQ9MuTAorXkR+RKhZxggPO/LbNvxhDir/Wa
3zg02VlvkFlMVZ72WYd7Ggn3pw+6Vithy5KsapbbXPgda8/IaEzwQDihDi1tjWrEYqaMFgQpEARL
ZINd80AOypLJNnHWdbFoEzj1zemslMjaJZ8d++cmbEc7mgPY5EYETjAPlCHcjgwLOpIas3EZjZw5
yg7U+ZR+YwQxA8gco83jj/XP2dmFmCWo3qA4arpr3bV+zSsDX62CRJhtbdvE84DMAVmkjukYo0ns
WXU8//T5oHgliPE8rbfAf9Ves4aqj2wnbl2diCST3Gt9RdWx+GULQbjeuMe+HAmys+OdlggPD1tq
b8TxxbToBfmTwahEqC6ATFxZ685tm4Yaac6kEFnG3E0EGLYwIQbAZ0LzrKZPlBxTztZWn6MlSE1H
Qwt4u7rEEls5BrLOyRxzP6aI5Wpf5BfbATLE2ypDgT2/7U3/0+wr14Yi4NErOAJIWmYf41QuYw+z
MI/1nt8tVE1r9kr3JAw+gI8H5YVCCkS7KNE3JITMfZFbFvA8ZBvjtmxFQWkaoXW36rmg7d1o3kbM
OP8ajd8eUStdskvJGIaE1A7aahx4/6So3DxjPjrf4sIx5YO69N0ie9o9G3PJpDPVLDa/QOhsjK16
N4Jt3LTDYP2+GRnsbq3w2/u3bv6efCfWHVN5u33QcHghA/pLsxVe/BfiJqmV95BOyTHmk6jG3I3A
MuUvq14ar8v5UrN5hTYGTBPhmILrmBpiUfgQAjNTflu8ULLU6UXpTVgWN98nzFk4+UDd7oQHGK5K
2Hckl5Lu4GnMYRiLLnE3T6LKHgtoUJrHWEOnyPKG3BQBFHtMXYYylUPlTt0sKoGypxaC5qct2R4c
9uWmGOex3jS4PikzAlZB/SPHJrWL4036/G/Vujw8fLmXRcZEBI10ypcEMCUtibJpKmRqZjGdACml
SxhCqf4FToaektYig2vpV+lBggC9F/1dnYlw9holBMYT6IW41BXItH7BtZSN/+AiCqAj2+NT/WyX
vym39oD8oK0UBZNf2vlEd6PwUckw0Gt1v8uFLd1jMEh9l0uIUSV6QfIjfnQlxGuSEOLIHh7tyoTq
Wbc8ErKRrexmCk2n2B6Cz7XZ/Sv3ofkPwVj0AUR0LvkmZX1bTRMb53aLwRnnLOz3Qens4Zp0fnko
YIP+rfziQEt9GsfNOsxVWpm5+dIrM9L7l2p7PLtFQiNRvGOwRvsDgaEaAIO1YL6IpHIpgKXmgOEv
DAD6z3vmYSIQLks15C1lYQc11hcskR6PlsMjeRVfrxzI2RCxnCrxhvub4ZU5DLDxgtg9mqn0jw44
XWQOi/dHmEsQoUABRtBpZO4gt12YHQNJDfPRllyWmI8NT6RB6760945IFKpcykMPGGuAoRRQnTRb
oB0gE5ZBT1aF590sGVR6ZopbQL9ZYzIzW9giNSzlbXZZqO9/248L8aINg7lEyfXwHib+0TuYX1Ln
enfGxCEAKJX0VdLNNttwsdNnFfyS7FcPrmumaaCObK7CKaAo0Ty7rSc2vhb7P2Bjp6cbAKYp1gZH
ek+ynoNKON1AHrtwtnnBUBzVp87TD44ynAZvGaBzxOabKhL+BNh6XTwpw2/hmCrYwcwtXqxJDTRL
zBdzdHhpiiWE4FfMoDElJZjf11kv5Qy4+1VsbCXBgoWDQ8OWP2UclWcLiiz/UDOPeIZznUsP8Jq4
tnK9Ehc+pZLix4uQFluTEyVVOHkN5ohcDjSo2dH5Jo7CMqqkCHe5AgYchafYR1qbTq42wFwdtfAy
2cpd31JcK4Hm1rcDD9z+KSW0duhTxp+W0wLEr/NbHIRnzBKHG/iLTZgTSNpnfX8OS3p0S7BuJeU0
wDZs7LJFbEwNPYnZAPisP1y+k8wsNP2g4XwLZ1Zqxmfbo3Il56etnnSTPBMwyq2BzVGDbj4tsXTE
3V0ETL3JROApmq4XUcKXrCz91COxJxGtHlyfEWNdWiYApRFiCSSd8q1DQQhDYBlc1XU1I3oJsTx8
XQVfYAWt6TmxGthoA5wkGtR2/N7v/y5udBszYMfaxl0of85UJ7v0sZmXYDT+8bEdx2Izznm7xtHk
m2J7dwHYmyd17gX5qc2wBmwfGgv5B4MmFmBorywi2lULQ0Kl7TTdpp2gSkjZGdpRV6SAALG+m5qJ
djkezyeuugbXy7NfH3fKhA4Wg220cHZQG71HAZR5XZOfBg6wYYJLBhc5D0uBRDz8phvaHBo7vsqO
XUrr2P8h9DC86oYZfWrcErwm6E8p6AlO2KABv1ykdXVDg5Bgug0uWaD6VLdQurm6m2s2irlyxbm/
zotNdvWtkL8jwEMsgT8nZO8bi2WGP1C8fd+fwwBiAAtImHrDKqxUaeU6yRt5kJCLnu+rKVG+IqES
Hmbx9IGXYwuAm4zIwkLbHAyWZyrSJEp3z71ZwMU6LRLSrh1RDbWjL7YzNE+BDMwgxqQSB1DHBpa3
tH6WSVetvswDSfV1nIj7kWpXmVsU8U0ag9GwMRO7IYuzIXaNaUT8V+X65dnd6SsWc/szrBf8BP44
kwd2AwW77ZSjBdPI1Vzv6GYafUn/Zp/Vgnt2n2n9/x7RA3KtqfjMdeLI5AMfeplAxcXwQYKfa7UN
pJEbwqRQACgVH82Ynk6sBYLHqLg47wnmiU4SRzLJx2PscdLm1hTaaTEqM0gDuBh8TIXh46j7Jl/v
HQ1S1fQyFwazMnkh7FKjt6DYE8Ch5pmkgoVHEUjgHs7pLrkcrAYWQcA3mQxbpJpjlwijrrfYI53r
5IKxWCTIAuGDL6r7zrYTBXgW5SWfRB8AM32LjGaD1Ddt12Gb8OcbvgfAx+ZBrzeNS6yeg32VCFC1
zm20YBR4xTT1uFHy/vTBsTKjpurseB3i45wnfGt4twuzs3ieSujzBlrVdYHuNcR6B2eLwUHadGJy
uty5s0mxxiXPEoPGoXJi0CeZmdDiiO/bFur382izPA8Kvk/mHan9k6M4jQcrbLiZZmu952HqF6sW
9DK/4uYT0BdhAPchKbC7g22j3c3Ei8++Sk0LB/atFJRpZ6y1opJt3/Kgw76Q2glLxmTH3G5iXhWP
+C7tBtM1+MOYyizXXDAnHJ3NBaNMmLTBH9np6W3cbuzx1Q44Dm1tFE2Ii3fDJ/qElIoXUP+45pSW
91Apf+IDllTFetBPclYY1RxQLhHFpohsz649txyXqED/FWXKlXiKhq/+jnRue7yMA7xisdPnx1J8
Ne6cSwGpHvuGfGs3Ba3H73YorTIc6AAd2GSivge7lCJHu34grynwxNOJe/f5DtfcM6/btmumk+B5
QLwHnl8nyXbRWQQajoD2NOAk6FBDVDPzy1YTHezrcf/ZCfTZi9BprY+xBOLsV+vS5y5KuJ7JisUq
9SWG2lQSRt/jdSpRSoW8swgySZFK2gWGTnsRlDmS48YJt2Q6NchDkKUIC+pekWuJfrz1809ikEGj
g2ctPqLshk1atYI+MGQAUzA6hkp1v6/sJt+UryT4gLbrWMXHvWhD2nDKTg6jXg1OxSdVSzD8crYi
664FlRgG9No5mLu8AFvaEn4KIV/vGlgHChPJpMKIoGd+OMQpDRvnUrz9EN+WVuJGxwr6j4RF3pXd
9XaOdZ2NUkulNp/pzIXu3Uk/2fOmfOCAl9LrIM9RDVC/ABSYZYrtRVzpf3zbRqwcvhqwXMKgKvf/
7C7rGgbUucuJHVjxLuaLKaMgasTeoHy+qJ5yxGvV38W2its5HyBusICk49RF3BNIcJ38ZjC80r4y
lGLHoiiIIerq9T+7p8w5yaVP+er508EWyjoba+8mbHCyPjz5FE3O6+HU8tSYaTypsYdqhqTn0gZN
0pnB7lyPX81lG/KE9JWJG0Atdv3IKHFdnCekY8BiLedf5XvUw38QCiN+wHPt6jFkWRFC5A5PD7F9
YOM3s3QctpdnqCX0q6HFwsSKZTu5eZfy/roxS5vbGrvmerGppVOn7oy7IQDPHOKZOD1pKziqiBln
3eoa1IzEd4fYp4uYpvfjPgOMIMfGvAoKIQ5TQPcm3r59s1d3xateF/HAkCFlD2RsHgMDWlbZankE
ONu8duDmu0D+JBZrEziEBrQ/hb7YkwuGJIhnygvRzRsxtzg2nHScZLlLmDdWzncb1yb4qTpilBM1
XXh92z4sDUzyVBjlFYGvhIotIy8NB4qTb0tjSHUSavZDP5jaOgyyKwISIl85cR3XGtEUqLfvsLgX
zWaG1RoPxFpJ5JdVmldDJ5eHk9KZGFBsJFgqd9HZkXL8Es+LkL5zLru5C1bKwijdC0MjvaDsqQ3+
LOdwzVZk5VPgb4NGQWIsaiz+35+q7R2eHggW18BggyXA1A7P2IA+Q4hqLHl/wiiRyQmnZxFdTXiK
rHk8KagcQlZgtL8V4Uj2dYi1VZ1II0XYqLqzj9lPBccZKtmUFHvWoJTWZviDQLAOINa+dBK7FVwB
rtZWJTEyr154kyLz8LJkC7U3s1qJi9VrtrKxeLQ60OkwduTW9qy04zjQUr9VcJGT5HdoGAFo3Zw/
XvgHJWFUdYMwihLnj5sCrEm9eju+nRojM2ph0TulB4yZ5dA5rw6mrXF6o4t24rdFDQmZpUyIoAsc
tZewVaN0DusNU1T4VEwfhArJhfCwvMUD3VK3UX07ZRaQy1C1l3cv6Te3KrTQnAceaKND5EJ6OiIS
NFwYOPgpU2/WTfyIvhy7aBn/1kes+E79oZ2CWac3F81wwcMFh4IRO1X/OzgmA5TDoE0NUvMFC0sY
brovPGGnTOoFlDlC90b7xTPkpyJSvLMhW8DWO0Rh48dIisxhHr02vGdkgYpN1bBQSoNyLKGwONhK
U03UQQiBmp/v9juhbhMs/XogE9r2RUf19DiH7tpf304y/q6dWLLkfr7JFluNWnis+W48NVfStbht
5Mizs+fNuao3bLVHdYsp7hxXG9gxiHypJwIhSdNpb9AaqYg/26NrRd5T3Jj84Mku5GvWZ2xixEiK
mxt0ltxYN58tGwl/xTCD0du5X4t1eUTtCcx/s+zH1QVPmderOLeeJyKIzlDdy5k8moQdvRCpPb+J
1m7c1ECncv7LmVNVR06nl5agujPs/DHQSZ6kN8TVxoG+GJtSHlgqm+w9oyjDV1g5xHRj6CUfjxNZ
v84ctQGmzvXG5m+04sMLdQGU0aHdj0iDO+Nbvps6n+fTaqNPPY6bfSBNfgI/uaOwaVritxxSKjC9
RDbHwGRGFG+ZovRNBBrbr7LbKERULLYds/TEEwVy9Xxi9Q7mB8NRgHgd9M/lPRDh2k6dEYEKSPyd
0nEMj1cy479NcJgBeXQY3nUyhjKjluNweOnenkf776SDzRAYJbN45Kqk8i82z5oSkUa41IfOJBC3
JXUUL2J5wRN6/hnB0/3/bhWakI1o3FHr798VBZCCjJ4U1ojB+nQqYrO0b+ZcBYnINgW1B9VFrxYE
vIk6GTbOuFIymJyo+PiZ6jlovjQE62VfKznGgOq3mF8tBiZ1u6xSxpzAYAq2SiD2Nl4juPA3Lp6u
6NvpS8DTo58qk1hj+zs1SkfheSCIXGDJR8BgkW+auhU3zuehYdRTq+Wra6wsN0amaYt1NVT7S34r
H9YTqWXWb+cD9njcA2h8hpr48J7H1LK9kZuaxeBq8hXcyjOgrBcfTVJCd9AKTBtLwO3AnnMraoA5
jt9LiMReAM91sm/3ICU7t22fGPxYodcFrG5s4H4CiJF8XNtX92sey+M+Dd68EhNog0t1YFsDKQ6x
RDg+k/30woWEGQRsFn3O8nHJSTPCua9xjgZs42hzxcvciI/QT9PM4qBbyRmpx+fozV0h+DU/Te6d
wiMb5cn9Jv4puTso80eaKNkomcBq0uy+cc8jaQp3wwCUDYWuX+VIGDG/Ige9bBmipP/wDqTPuXq7
bJYPbRzbj03AC5uIo+Xi2TkOyFg/j+mmM+y7O+ZhlyWMTMY41T0aVM3KbYhgg54G9KNqjGudXMPx
hpyOhcMA7DGPOlnKpBwnmp+mt3/kq+QKg2HBsLV2B/R+eidrl8OssZ6nUw/1gMgMJS9D133DXku0
y8BRfFZ/lUO6KEk2HFfQNwhN8K+AgfgeYGT8pcUgaZWedfCjsx6AqBDlM+fDO8ZN4e3JqmE8Pk/T
pGY7tOE0tk2Ssf+qOsPv5+MC3eJ8SVxVuCt4WxbQktwueWn/h+gZcQu/MqLmr8F94nfi3jlw9EQa
2ssg/1dPbRbOv5DRK2McfiXzNzpRcK3I3g5JbAqmLNiF7QeIoPkoNaN8dhgU62CCnLgEVRiYQoD3
6CTZd58qHEsu9/mcKfBw8A7Ve90ixIdGxbPJJ3n1j2Li+09d40B5qJUHeNsa46o2Nd0VK9xfHVuY
pLMeG4s6XB1PHKcIcvQwoCQEjcJq8cl1k3Oe5F939wsv88lg63A91LSdKxg6d6T9blr7hH7bG0MQ
Rrb5VztXuegUZDI1sD/4coKJGxwZNzsLACVFkkWddwIesuY/5D/9qzVG+tTBKXJ4NBkXCbxtXHZn
o88x1Uk/4smcsSvAeZLwVn9dTskajQWSZfgBVJRDLWHPwrsIbCCmPAX2WCqo0f+ZKGbC8bbJ/HwZ
Y8LUOrWQAlzetjBXFBF9cc3v5oXG83hkp9+zJV6t7RS2ErFOhkTQIALF/4XoIa8f5I+MvoLMpniL
OdIVhkZkSRalexIk4ZwigzWDU19yWSEoH3gQbu0KpACDG6ciB95SqmPE/HCaC7fHtFQZDtZ2E7ra
W+/2yl1qdoUV82UjVItpMUCswf6pFWoEuo0LGV8M5zB7DOdOSfUxJ94+yfT3zIkQ+AxveX5s4w4Q
LP/1IjZy3cNnJzMA+mKRwcc2tcBfRkV7Z7bK6Ig7X3TfZjqc56PV4vjFFlJtq5HWWYYtRuYxDm4d
01AxIZwcMB3j6T6ebdt2YGSu7G3s/KOw7KFg6JYhpEjCD4hItMlXjqIszNKhhQufTUL1INoAXdlA
6uJWm/d15mYq4vUgtOckPfgroTmlE10MCUEV7qbiDbkctENK6WSyLFAvjokFHSf8AExJ/xDJ+olJ
2LbJwjs+mLQuC/NDyRVtjF6CVAcVdu9+sQMXHyTL0+uDU2l4rXMZpPiFYUKakeDMgfNm9YpvlJCh
VjzX+m8Av8HCxv78NjdhgwAQUQ1YyNo2QSkBVF11YnLWGAl0U6YgnjFpEiPwKyzYq1Z5/+75w0i9
7OBq8iwV2eb7gfobQ+JT5OFsITvxvOCoDfTEB6Km8LkN2Icpraumqv1VPu4xNmp0iz5Zz0eopjFp
qu8r63nzgOd7h2EcJL8351EVrq2ilGmkyEIozyCiGZdNSZmdl64E7XF/y/bu9Zqe/pCzpykk6Xj7
8/scgM2pLSEgWnBe5wVXgvOH9+FGpc8+fS6FoCMcixEYlj8I1g2pL3rR42DcONeRn13CbxGbv/qK
H+UFPHqPz5E6JavVbHMzemCavTRMmA0Pzf9v2uQDNWKm7YJUns6OfCbH4KDYEuRwNDNOe61C8PCB
4X+KgOdFcvZj0dI1NifP2MlXC2vW7+Y+ewpULQLL20K0+Hf0d+cDZWof7cKL7K0h9vFtcybCz6Sd
y8aIUXyUXcSDAYHt0gABCftx8KsIJb2SW4+4DFOMt5ASA7swNyi6u1547EhUy+xK5X7J9LyP67gr
RrfkQgYvUDYbpkQ0Zcuy5trEAH7sSzZUidbBsRG+Jpgm4IGtbzyWQ6E5Mw4NvofjZ8i8vs8duM3s
P8YXr9zQ4XfZ9vJSUCDG+UGBwWVn8rLraKknOAQBrLM7vJ9KYrp3+DmDXd7mzJk4iPfd/dZQA0Tx
kQrzGsGxcWzv3FCLUN/Jzk8FPdfnpodhAoOeqr92Rkeo/PGTOeNikavEMzWnFKQ8ONKN/ccWxAfv
99Y3gtGUr6juJXg55KCm9dSwzRLek0+sRc7wTDop7kZrcBxP+fVr9i45Y/L/7zfurTZsFUAMD+FV
DHpiC5nPV39kLTV/kSR3ZCuaXFlUnVE5z9tCgXAk3BiuU3qQBp+H9oCS3Mf1p/VValvq8nd3xUSf
AZOPLMCgLfzaCQuWTTanICZO5/f14mNSHK2mT4zPbD8BbMyj7qvCWA7Yb+54wrK3L7qCUTZtmfMV
qXnHLoV5rqU8eAwfpHDZX1vM6caIBgqsNcpsxEa3F1uYvtbigdyp51fJIPtujRz1tpR/mjVUz3ZV
DfpBPHu9PSWv8NKQvQ1KEb+cONsEaThSAmH+chNvaTxoB3OwqqK0Q3Zw2L+Ju5OBJo2Yq1dwJlF9
0LCYKcJS6qbxzT5jDn5uEVAKL+PylY3p4LhaVkUYmRJR1j0bkqzwuTgd2Is+k93tqJcg3WIRzGY9
J+rjisyRPYgj/4MAtj/nZtrjYFNy20KvGc1V4Nd0oHLjeCsdMi2hWdsnnAEFpoQvxmXnEw9Qsd0O
KA0mX1S6fa8cfNS5BWpEB16noGAIwA/jQxDaHbSAsk5ctxOVbWBJBANzbBaXYNRdPiy9BVPJpQ0l
ncX9cYkxpm7Zj2GjSzhr3LtD+Qu3QhdY+kQ3QHCdfRTwXHmMUNJxZfMkl346rm1KyD7OVIDRTvIe
T+78NENKAV9HSGtSxUaoA4p2jzj/hslEUhMG0b061OtWxsnfjPdhAm1kc3clKca/6PUFo4ZRp0LP
ssVA0HO1NlczDWzPwsts3sF3XRTV+evQ1a5p5ztHzTyWBNr9fVcn7IIqPe+U47Fo5BpL4PAkDNgd
F1QNWcwhD4eP2WRgLj23OQsF0lTzWZztIyeMYMWxIvLXwGz55vRMf61MzHqppo6a6bK2g/wXaKYX
pSCz1ccW+zN/6HPMxKuX76IA9MYzbyTIQPvB32yR3jZqrd2BWii1mAMM/dsvqf3aE251S+JYMEia
/ZsC7pBoY135c4bBWcDcPS2zTtt0df5iRvkulk7PqUveLwKNcVdxcd8cleuVOQGKKcgSo28x2lpr
f/yG8vi+I43l8WXCS3gF4VUYFlkOhUbG1mzb0El9eD9m8DHLSs3KmDLToHHWsENHddSBjiTDklZC
P/T/ui+diq1ykUngV3xE6VHmcMJuMdXIEHF/cCXn5bQ8fXyw3UHI6IRyCMHOnsdNo05AeGWyVPDy
nYOoD4/0TpD/vQRjNkZwcXDAiDieiVotbWCCjThUHddDWCAtNsorvDmkLhG+TzqniiNbxTCAdeEB
PLlGkqYeBZ3LqozFhCxzijjAVub+Edlu0MwVP/aNmCTdGF/wNIvaPXf25e1raCsjU+77GjIgsvI6
WoLYF3oQQ5Is6aiaKRXwKUoJ84YRTsNsENMAfbzVZCD10f2nm4XnnZ07Mb7P9DHB2XI26pQHMk6G
SREqp37vpxvY60esB0jCGkw4d8iqw5WxfZQXeDpweCT7hlksGMBVqjBhGKFhlP95pcPoTRG2zI5T
cDR6bOHbrfn3LzgXFoJupWHOr5ngKpFz5qSW5AV2t/o4+uctO79FfKsj75kWEr0rjaM/w9cPN5Wz
MT4hT/vClQJxSLGE4J2uVc5lAzHcScXuYXcmsOQ68R5EXc1K1i/ylasAsyRy564XhdM+f+NTwPip
+QF0x09Zo0Ob5ao9+bhbMGNJ9WBzUECGzBxAzPdHacfKCpY/igNCPxBXgwJEX89MqZzY5JQOwv7p
fxqTS3/tpCP5PjSsLH59YkxbXy3RdNOBEnK2Br0xT0FPdHGbhp/0lfH7HhEUfJJzPVsjC1cFHlWs
e8qVAqFqyuxfhMrRuZmolnHaUGFuldrpAQGOBozEMYM6XJT2DdmQkpGnBXIaXV6GSg62WP8CcaZX
2yeDN1UUHEAurBKGLcXfyZeeGtFQHhyHPd85PkxvQ8gKs2ZRCp0zMUKKu4DmRO/B+Pfkc0KSiNN5
xusv4GsNJzuedjuSOiJ8L3bcKqWuYOFKMPu9SmOC7lP2TJE5PVYlfxbFz6VPe1hzBKRKr6r8kTjD
oR4GN+Se+3QVeqIxsr3aPhK9Qyha0ZQQ43jpFtZkftfiU2JiU8ubCJIoFfRPL1q1h+O/x+bXdldV
hJLbjzFLz7EQJREqeduVtMhjSpXZYhroLMixRYc5RxQRnnYwb+1tP7VDsE2+KIrr2r02dXFl9uhr
3PjYaEtHR9zc8adg87o6N9xEsQUXynDcV5aBGDWzsgD+HAasq1WFlFtGDbTvhwrMog3NIeSDjgwy
kxO8Du4Fr0rcwWcUNI8zfPIHNn0X1lwB87DR45ppLnR6cRQPV48xtUssyQbkb/Qqtcwqk2KPVwaj
O1lFW8giu9gLr83yAM0oHesqoSjSTKyfLCMLtylmIXjgzWhzeJWqmlP8mA94j7VQbXsTBh5blWV6
x01R73xL86aVqp5bLxLFBsQNgSnY62pE8aYkrlAfdqGEdjAabHBaaQopMGV7MNsae5VRa8zU4J4M
dpAIVE4Kz1BeI9raw0HsmEtycQCch0Hzv1u/rWhaRZtN66u8JMlLnMk9FOUuBheOmUxPN/T/fKLA
Vzw9QRlDCB/kYyOWlc02okvHkPeZAQGkUjlRgLkA0h5P03lcHS357iTGEHV8SeC8V4BsGKZrGMHn
PB1x+6E0WbZ6Oig+/5HlGZwC0vwW7AMa2V5OSoZvsOmxRMfsI+DJQzAFmjzqTxbF+MoMqPzIWbyR
3HDGtXKxIKZmGEDaJPo8J+QYOedMles/0PhVg/6Xw1oZXuX2wh9cMjtWxLSMeN1Hx7iQlI1/VswQ
ugBW6HXXzvclYUp4+Q8BwPjtG+lpnoQ8MEgGHHY6uVmfW/eNW3wR9PH28ylTlkHD8GoYPZlS058K
t9B3jm+iLFfk8wVGoE3MPpwPSr+kFEERfTBhCyxjhLOy+m7OMLrJMjlJAytmWZKJudfvWbGFrLD/
5DtJwN6IA5NcpAWxe4n5KpzfM4Pi/g6QF8k9KCq9h0OphMsx07MfrV9IKVT6sqFhHWniNp9PbY3E
vxOaR19rmS1VL0913cxXCFqntmtT6pVU08NfpcKjMpN73CM0qBBufIVz9wjrQ1aKP9LOiSWt6no4
R90gyrUNcQgs2CdjiyFe0j4PVumgMANT0vkZTiCJSqQ4o2gA5tZrGccyFImIrmGhQE+dv/9SpPlc
xxLjQW3BJuxmM7UBHxHd8RNSMXnT3swHD/8qkbfvCl3BrsKo00wzxM+VNVviJWQ0uKhabGZZwFwJ
7cNgdkeCA99Y+nzh7gi9nl3O/PHvRP6f0Q0THWSrjQGxx8BAh1IFHb384B7NbYFeN9OBzP6b7kXo
eeTJvWwRCiRWoMrNCWnXBheN7RDXXXs8rn45RV9popKwIX2+5mVS8sRM/bsI7fD5iIx+sSAxv7F1
A9F+8tyW8CiaNRL6m6HXK3+DqNJlhTIkngWtok/JhiodTXDlehNg5M7yB4GkruXp0useK5URzQEH
+wizLFy83//0ih/hy+pXySvVQrjIbHTxAUf2DJFDoBjA7c1pidtmsPFz6hQMhxGxb+6z6KP98fe7
Ga3yHecfBwc87pEgPo6BwQGtZ5LAs4m8G4epWhcTuv7JBwWAftWGNZl9UdooOtWeR84Gqb1AKwhB
JIFGO0HGj2W3iVdLf17+tFwETjTZ1tqVODa3GvAz+pfUCaeBfBpTT/VtN9/xHW6xhHTqb2r/G4De
t7KxMmOvGcppaNvIqbgEosYsrLzRPBqX02IstTAVfTfnoHb0e+7I7Bmc8Ru6wn/Msn2/sYt82bvT
+wS6uTcVloP7uxMB0McIQjoExUEWvrFOUfT/YHbVAK0J4Fwv4mSEc/RxcpfjpIzlZ2KfirMICmFZ
VNXS8WOVzygm81FjvKeBo/cBuXsOkHSEs5odP2rWaqzsKirMsOey0zJ9uqafURjHEwH4sO2+0Ok8
wLxmormp5KHOUlgUV/zdvmxJXmLttjLlj/NTDO005EmoR6k0q3VEbWoosfv6WMnPQeCdKall+quc
bR3u/JuBAXpyfnWpZ++zJq+3f5jGclCwgpBVFP0txs0z8zaoJQRn7G5KNhDZdIQHphy8Xt8QTKFu
/sH7lULRPDe9J+Y0CUMv3HySaFIxI9niOhsZvJhr6jPM24VI6J4lh/RKgySJuH7Ulju4HKuVLJxF
PszWkPrPAihEjvXIFyrtTB2I2tpzxrYTXVAOE/MnCwSjyylalwxZD1xHVHojM4VcIvScmc2b9Ii8
hEIwiIh8eiBFf14Dky0JP455gf3F9gxFUm+rbTbzEVfdlLqMe3swzbyqhLvWWCx9mR9/+8qZ4+o8
X7dz3xEMHklINxB0uI3bi9HXiQmoxDPEPdDWbIjVv98pexN1+Q0T4t0TW1BM7R32+rbGKShfJkU4
89AqK/h/F89DT5tSOJWlg7tPyNWIobSmTXWxbLCIcpCrbAc365ATJ4dWFmdk6O46RY1zNf+dfdvy
kkHjJNgnR9ytNKRn/dgw+sHipmqitTiQ9PvwTWMccstUCw2v4h4KaMrZm4EKCaM1Z3K1CPBSlPh9
phlfE2DqIAjWqQimCghnc+K9TKiPnNWLIbm1OPolOVBBhswrM+2RnvfbFPhr+u7c+TO1deEauWg1
RP7FtHXJSzO55hC9Vx6NS57V7A1U0nUaoUkpqsABqvmHpmdVLLmmeFzMRsgs2xH0h6nQnXV1gWjo
X/n9DV0xyphEnZGGRQnC/RKnmu6+lLVETU8iO5SHlBX3jQIRLTmVud0V8nWdCBPOZFTRuyKu4xl4
CE3C9TfoB856/3uxxW8GIZqAUfDzwvKLLChdP7XwzdrHKrZHRU9gB5miyzfw1QwvUTprFilg4lpn
bwEs57hjMJpl09XAecJUC6NZSCThN6TV8wIyEOSxke0VgJvSXgsqkLP25GMqvgfZFPiXBMYvQYwx
BxKIrJWjuvuqpS8rXr+XsPBYzsY5u/KV43Nt4ogdzW3gGAtTCsl5GjTkFohfsjDUJyz9pBVsPA2A
HhhNEYhegVhWc0bXYNYEFXcjNM8ac5NA7Zz6UdFgmSSM4RpqdGgv/tLy4NTAig6gBgFARtoLDJdC
mrH2NQwCCWRbObmo8lGWqSKYXmeP3csp6BNXrwLeWYMmPDyo+ic9IhHjIY8DfhS2gnglVXnZnnrS
Yv2gMrmcxuKs5e/itQm96oIYvxRAYPNPs9tfC8+4/Lo/1PU/piY6FgKkH2JbC9zTigk24uNyiO4O
1WgCGKbD8OGrQFr1kDkgQmmUf0yub3Uju9/6s1LlxzEvwRAJA6mwDUi9ITeAzwt9Q2r4CU9ZtG3C
D+j53djV0jMbE5hojd68gW8BbcTrCVpUgjO09lUHn0dUZFlrrmjRVCUB0KgndOSUtz04Ub53wnI/
eKlt/D7UpSq6ju7Du/wOMJoeHLfiMDbgyzKQCTogPC4bdUFRMFM/CtWIRcNF5YCBzok/YwGL7Y1R
/bryR3dNfiisV5QSF+1Ta3/G6FJkA+iwtC8WKLU58PtYXIL3CikQt7/s0eV5hrwxjK1VCZvSP/Gi
PNEkhrzwCh0nLb43Ph6TKLLiW71rzThqx+4lLGJ4S0gvvTD5GnI02JmhLlWj+PUUEvC/km987mqz
FDvidxaRAxRD5ly/Ta3gegEpXey48jtQMF/fDlYTp+tjKa909AJHB+B8TbobHyQlKKhF7tZHISs7
p8tgHgglPf+zCuO7scAR90XqdXwMFNuKnYPkCUqNdOOnzIHJeCAwMa2muNBoTnuinLW+VdgMlB8j
t8SejO9humdM3o6wvNCz4YweIoN5GudEqm2hoYTZqFtrZ4GwGdfKuwgFGIZNPx3nI0LNZj7Y+7O0
TdmAOQHAW+LhlTiRFuVpJdox7gAOMdFiYfwVgEVJyCe3g7/DL7+43YCIiqQIqc+UjM4EoNWWNOg4
qN2NtA6neIMsNpFcwkfLiDKGoOPiCLTvpPK19MG74IclwsXRPHxd7Lt9YMDdk5PY4+IYfrMJc/5j
DVQT7jKj9frELHTfhix/ohBHWIj7xcWPhHk+Djbkfj/QwOrRBkudpgQDIehP26tGTaA8hb+hW9ag
U//Drn6yUUz+5eOO2YbGhXjADILH36NMAgCxSFB5iYMVHUzG6vpfVB8KV6LndarlPo1JQMSL93cv
iojCw3CKhl8+A6R2pePd2qiwN0kJUsP2D4iHCDUf+DPiSjny7vF9hoBfUI5SmN72tHC3rhU3n1Fw
P+J3B12OFk5NL2yQBR3zDxrIR9zAQWSq8Nn1NAqUL3Bttzj2ibzFiRDMkG720BSf9sGmaRenz6hv
zmZE/oag+ACmqXK++P6HJDj96d9NB1Beg7fvvnorOp4rGLlsZ/vEFd/4Omn3v/shl5eRRzXz0FL9
24rmfA86zjaoLOQvZ65ZJ0E1T9/hqY3eFRpJ0ioe+eLs0FH23bxYMyFuF4FUFnaZ3Q7jdb+z6GTE
ssYu9RdrtvBzZ7o/WrcNddRIgCaP0M3iCyZ1dfvWA299DDzV9CuoHyd1gZOlGDgmoowFZbvZCsVp
/3Z3MwSBsan+JQv302Bqv4V9dGFJrLGDot0Zs70FkVVNmc/1MN36SF0aJYMc6w4v4aazCYdhGmfw
lq2Rox3AY+UUj2RLz42eExnOz6r7reGvzVWtWNFDkH5V8o7AoX2r1BdQoBWNyQo3egMxcarW/uaf
2cS2LKjx2yiIyN7vCdY7wpslU0v9cYEbFHgY+pgwanyddQscO8apfs9ERM8dxt1I0LfMmhB4gAdL
UK7zhMCbAIrM0tc35YcnHG7Puzv9CVzrqR1a9Vc9q7mUb8KKzIzuZ/s6MZWAkcAoyk1UeA129UKj
l2IeM/JXVLmXcKVmjI7yZZzcKAXeVxYB4N9OsXPFHYRYHeoxHLxXTlBrCTWD1XRtIDAgDYmuI2ea
eeXl+Rwee8VSQsjMYWHsy4RvI3nX7RN0QlFdcM9YTK15/0DWIchdX+95JD/zb4v+OUswxI+mh6Tm
sMG8lk7sAhaPsnil0wi0xobNUJwa4CcI2qb3XUsFfamLKPjMtCUZUNELVU5Yh6j7LzL9vRmFKdfP
2EUuiCK/+srJHHe8c0b1q5S3m+sW+rBbS5JoLXTfZCqxnsO2jJOjreZRm7FDwQ4buTEjefb+39BB
L1eG8wV5rq8k4rTdGwnIcQGFcgqsPl+wKMC50Mm08wDyTjyI8pgHCu7rLgWTXvhMJ/S6zFB6H605
XkTGOS33S+uMc/2mjKXVmcXxQfEB9QPpiNsDxx/seyH8kwEXlr7wNf5S/0dCjW7qzYWqlck8jakS
AEtoJs+iXfigHrKLY9J7Y+Cmh3jPAkYlEYEK/ihPsvwPOocrKjZVuWZn1QxSpBQuqj/bgTyrDV2J
ussI0pK3H4WP4fUNYAeInjtT4GBh0ZZBlH/EHPKaPLDbcCijenP/LTQOvlPaA3Y+5aZH39eQBoSX
QA3TKCFy7f5Bu3QpwKHmWyr1jt5ipHkwhoC0AszpZ6aQxU/ALP3ih1p223gp8zUPOPfSf3sGJ1Er
kdKZveI4SmVsZjfuA5lqjXsSaSB76m3N5Wwmrr/H9bchAAKy9+kj5+QGNSMVe2rWy4wwmS55WQzc
PeIJHH3wa4GdkGkTZK3rWCdFUs3v3vmtyHqjUQO+bhswsZ4XCwUnzhgkB4bdb2jTQSm15mP/i5RN
c0K5YE8It/mC0EZXptP4MOY/+KAlV6En2BZfz5Lem1LLyyrwyosmo8cVbdiJR8G/eKlbFTCo8LFb
nsAtMOKXoFYUlWFSvsdVBH4Y1ec2FWYfCfOiE4ZfZny1PwVJeG8JjaaYK6bKpi4HGOhKLDcxyqTG
w3q/QLn8m8XFuLzGLlyeksoGEP4v9SHvJT4hWqaMr3omB3xOlvIwx6OSBU3HXt/y4aHLbnzaTNP6
j3Zgx5Qgtt26BCavPZ2pKTLZb4nSA3032qEFJIJPhCa+JnOU6aP93hZo9A43VGyvEvuVkEMdegp6
tqyKFloZ0JXJWbl6OgPJwty69hycQcyJpw5cgLqR0fBC+w7TLv3FfsF7+XMW+eiEsODpgfrLvjKs
D04MnYUPOvHDpYH9p1k3dNzTVrmOfCKpwDPrAmHXyRRX9Y8ZcxZAXV490QYYvvMKYhA6oTrS6lSp
OwFrzI5qn0AhnPq+2OcVGFKRqQJXU1tNR99QMO4x9xQknx7xMVNWshHGK6Gn8FtrKvTASgZNyxr5
TWMUvd9fJfvMfYMAgYZ/r24dywJXVVhDuaDvyuJ7Ds8xaFoG4/FnHGTbZZfgZbFSH1L/7sDIh4QM
QkO4HFQyD7SeHProzC8iDnJ53uHNrheJyctsxlbFUh19TiRXipx+9AL0YM6QOS4hd/sCd3woj3r7
CyiGci69KymGo3l3HVbEP/w9Q+OAf6pdBp3QeYqGQSz6Cknt0dSEDMd55p+xLk5AVCtgqbsWFAgl
vSqtmLBBe6jxzRMGaIepoInCCs/UkBGBt/3HvkVRWakZX0i2lpB/Vl5H31fMHCnJWdMqseWTPfiT
SZzi1CYqmMVPtJ6qmuG/qI/WphpZW1WFP+a2ev9JxBTWQOFb0nwQs025K5UGzBp9rrqc3duYYcSY
HdEYs6Wp+FUTbwTctS8eUtJVNEWjP7XH2eVqWLEf6TwGPwIVVHRsoI6cD1YCA639RUHka/MN8cEx
xNc0Gd8hQ5J9LsCKXDk6qDaQV1+Dz2qjr08Idqp2MORpDeT2lEbL6IklDA29QK/LeyTpbXUBelHi
As3alnhDnQk2rRKeXz+IOWEk4HOB/m3imwtI9HItUzRw2wDxAbNtlTB7a+pfYddBcV0IOunAJL6h
gLoEYrL4/4/IdcMofLpsGveHwU1AtZ/9cJUA/dAvpy68iMSIPvDq49QcPQmDSAgUDRzglQ7dS0pj
JtOyvcPTQut2+8pSKt9JN5SkSw6A7I4k8sLKijlweVGG87keQLj23cmSC2Zs+CDSsb7K/HLBmmow
rQn5IC7W2SCcMzyyZ82RamFpCLYN3lkEcmrDbgGif0bGTFXvpIrTq2igy3p/MUMrUjRJk+cOCafo
0sOtKFMiiFZGqzMZlKf5Oo7OpOArRYljwvutoynipmHAWNWuea76vN6YL/K4PA/caQBFTY9HlBRu
/Ols9Tad6vRl1dMNlQVwtgZnoc7OCNW1jl+gk0ssPEAzeVjKY/hKKBPAI+E/kwSmD1OUfWoOYco+
JkAB4iWmUGK7oNUyo/9qoCrJgEwtbOyE2hBqQJ1ttLenTNsqvWRRfaGAVFkM8zDJeSYlix/5YdZo
zOyOTir0l5EidHAbBCjTB4H7GriBoJZxO9QoOPbjND0QnZLIAZ5jQV2BDUZgyYPucxfrO6P/C6xb
fWyEFra4mTkBBnmxWXur1LK3FBNnbiubi8N54wiP9zOvI0UXLvUR260ZZDvdUvKTynXaFY0sDPgp
eO8M/N9SSvXi5UaxnQoh38lBVcPWVthA3dcHQjTGqMPDrNEW2QxGcf/SFsm9T14FAw7uFe4dxnm0
FE7elJSHM0XMSN9g9qpH7S9MJqMH+hKLJ+jgyju/swLMaKigDSPbstK5TmYGDUX452+Qd9FrUtM+
CFlEEiZADLLBcJZDnN37MoDxiQpOnB+ogsCu2jQq+ripkfPGE+RhX0eeOjrv+NK5LzkYAYRmYWIv
BkTfqDQkCs2VkAOVRRoqVC3yu6YnYTV9Wfsy04tf34gr6xOj3hzN5zW3XmnCfS3VwYjvRA5evMRV
mIY9YR/pLMklUrMM1vKtVKJaES/ujONZbLauxoenASPYbMe4hUNCoVfki0k17UJsQBsJuvcjVmHH
EzsKaAcv3aB++g0EBweMED6Jx87lQ+s3i0Z3SkdMZg7gcBEGhNbSqILjfoCqs0PgUbUjVXVSDhuN
qAk2ez+s9heq2jIQ2IVc9gc72BjxtNO1Bh49CVGwwbD41JLY0J9HYz0I/L5IN04u3q4bnMWgTXYz
AvNwdqBifdi9clCrr+Aokll+6Lcm+3NrmdVSu6OXqlkkT3gmPg9z5m8eWlK6MUV0Q1N02Fv/kV0C
zMO2dXQD9t1+2s38w5s/hA4zMntM8LATWWAC0dRvG2oX01kSw9n6MM8e5a9gFOrFPKJMdpBXO83D
I00MCK29pM9KYOlBI1YUQEAiKklmUGOpBF43TZ67MIs8fpIlILLdmBYjQkzo7/y05+4aWzplieNH
4Uvdq2R2t5/qv2z9UWgqtGetv7ntSoM/SJZ//9pn8O/3/KwpifV4D1JM06JS1aKGCylNbBU4ZlUs
sWDAicJ+I1ZxuVfLVviwdKh4P7YQ+iex5Q/3NXwZ4Z09klLiYgtaZreli6zOlZgkwEYjhIG5npHM
RjNyoqBxSE5rm0Jd+xlKMHPLb4lLTn3LMmBfk789koW/xSABo74ino4jFLdmxVbyOUkBHP8DKFCk
Cm6S2mVUy4mPCq1cfOCbwWNAd3Q+6H2V/AAN2uwk0O2cto4lzL92U6UMfHW6VOEk1X8zseoAmfar
FABSAMyMjgL5KBfCWsU9O9P4XN29rXuTYMlWgqJbLwfmJn69DcDsWbGErIcyJNpBjQbRTPDKrKic
hmECjnm0YNPfX/dRx1OXYQPB3moMmygUylcjp1RXucR0DoMIDpnLbfjrlZzQCxF5ryIs7TvMJ+/I
0C/wAV9DprUetlcNJH4J9inT+wIiDBT6HuS1GmPRAgkjXKVD0uu69YV/AILEMALmFhJpvhSZ1vs3
g+EsDzC5nXHTPcsKOHkrgRAcCL+gX03JsSlU+QGxeVzCPfc8RoERHlipQ4vx0YBKxLMo4QXyLDT+
n+pYUM+sOCuvG1P1gIolmCxuZxP1L8nyrA8qjHnPN1LHhhp9azV/krO0Cr5BfT1UmL0/ZaYLSz0r
mmI9RcRy8ot33brtcjfEE9m1KHHfeq0JBCmO0VjA2Q3f1stFQyWKjQ742K/3AsIQvZfCpunHjVcq
XSY+27d1/3B5doKmYOoENs2K31Ip3s1NnxN3wgQMkMe5rg2ARxAn1CRkcChwCfZKkfNvrO9+hamv
eMq1Q+wREH3FqJtZLNoDm4L8/+OTIcKKooqU3n65BFjvfmdUDhjpXB8OsqKcZJV3+jQXaq//7njL
U1HM0JXfP1ypYZoMA8jleJwXgUKhRELh3XTdMXCKpnEuR8x+g7Gh+h9YTFrRr9IjdhC1qfHsl0jk
d1w1FeW9E6i3DfPOVpWA5e8SHM4ml4GwkGeGmuplwn7zmnYiJhzfm9M12xiEmYgFEjV7YkwKG2Ll
iWTbE4YXF87aIIEw7sstBBjvWSww1thbIeZX9o1MmH3PepF9go5y+Bi09JYGQTNVi9pUOM2ljIK3
wdU4eYpgz7IP1DRuSlj2WCROAVxKw0bs5YO6Jb3VwYELMOye3IEcNRfgLDY7Zjs38CL7HpNOVN+P
1qy19bDFfIuYZy6jbhrh5LVzBEREsc2s4V6jtQx/zXRCjI8SciQDyW6D/tRgLT3kkVlUf4ZeI589
KFojDeb9HwDVfTupbt9z/caMQoFHOCUWjW3Vpb4Oi0ZS3sIYuK2WvSxbZhdAPtftU4H0UDDfF0lp
Dlf/9nBv2pToembV0FvE14JKxgvC85q5D1F6d9qIn8JS8dV+Gzd3mnRokamXZYDrVSVRQybc5snA
EZbcfpEJnddU5Aa9ZRwnC/q38MDmLhCUo1NMoLiT6UENP6d3VqW6oD+n1d3h/UvjjAwkNhVk04Yo
nYxiVLGwOroMCU+oqlg3S4wx9pK5SH+kXthwCJljddcienfKgU99nxx4uI694y/Uehv2nLhAooev
Yr92f+1Xa/Dz10ltf/USlsNQh3syDTY623qOvZKyKTscGOE4Ui0ahkkVvFREC+GiYW5JvEiy1vuu
99PiG+u7hyPYPxkF1QnlV3mM+oykCCmArqxB1Bb9Gw1X2udbz0inK1tzTqEM9Hz/e5R8NVYPkQzR
+bdmaX4uZH0wWaBxBjVqkmY1Euj4CJVAlTLIEqwC0iCaRInjK0RCBIs34I+/EBEwbq5v9G1mFBZG
FxEvmMqFD16VxHE8xkSymyGiuDkqYzHzPIpyJyHMrkeH8qnvc9J230sadvgWsBXAGUinxNjK96AH
dzYlmIZXVGUAxJiJxAJBmav051U7rMYQQVrdIKfKiPRi45ITu6XQE/lpTBbC0pkodgqRAHDUYzOG
/HSTPE5VNWSROLwJ93Eh3Z6T2COdC56kvaycoEhzYfxrqGtJurty20p14QAhsybhcpwgLB/G25jR
/xfqVD8A/mkUgL7BNogahopm597eyqT8ACd4HlP51tS242v4B0+PIG0+HrHV+UNhhggh0ElBKBAO
2INCYd17/rQsy3N9jS+LqTSrqUau8oBYizBvq95PoKJ1PHaAcu4zbTwUfCO2WAkPEQeYC9A4AA2/
wL6DJchPkp+l+UtYRNKaF0nfJtvoWpyzg8i8e/jXM9/+kYQ/ZzP3elXQWM4hunWHJzXKWZrb67ft
XAV9ho1VxI2GjKJm3P5KY7abSMYkun31ped59Rko78cPO+sZPoGEkl2IHipp3nDScafX21j8monK
kJc/S5FDWnL1nJ9IDRMLjluJbQOM/7NcHxfR3f8QqA4kOVIkE6Gb0+k/dGBf2B9WW1vFclavL6GY
n/6DOj/ziO/thIgM7rTNG9AjnHdE37sMQP9Cd+FdmTVgb8LVE9dQyfN9Rfpdomit48vdHY+z3y5x
I4vctN9vvl0XXIOyHQETKK8dnoxY3srMtmw8LPFoUQCpTX0zmtSqLJQpjg8fJsRRWP7tl+/5JRdr
B2ETV4P0DMW2NB8sBn0Brdg2i8Tg3V66rWhIGnNyGrGQteTXflRL+DHb3D9YZmVzL8koIbuGAiBW
tAxZY+BIgXVzundKrWKDR9ctjl70PmYYBslXNKfndhhCXDRIijLbLEejuZ5DhGEKwmuBUnzfy/Dc
fso663vgLXN2C8pBU80qzU3UJyxYnnHmM4a5KRYTu1mw4JY08I83ghoac7ORpeglybX/H0ROchoh
mnLxt6uETstNrKoJ603rKQW3etGP+leQgPzBoZKLpZEujZXTIBSi1rGLrf55RCGrzhI9F4Aeq+X5
b68FC/mIg3EpxNxIprKXCFPjyLhVxQLJ+nHJ2AfvCutSTiz22wPjw+48UfdjO5HoC2OXtA4w9vBa
PV4zE/iIsUevkyU72gzLlp+2H3S5lB2lWh5LiiFn7Nns3S/ZCmhMWTt54D//F0bwSMQxBU59HKQw
egHYJ4LKUgvnJRwF6yD69YvVIGchksUdIGY/fZuu4n03P+RU9f1K2FcKWvmx2ZS9fnqGnEfpQrXO
lmdmMV6Oibk/cylZK91xuD+H8kOLYvvN0Fx4w0XC3h8Qwz/raH6+V3CZMWdUCk8SdZb9GAGYHT9n
9glqTZewvtSGDJ4uLzuMJAdTx0XUZykstrtnOLg95tuo6V3IlJ866IL/6ZY+FZsWCDfZuirE3oUW
QLrNm0CPFd+2fwXUpLsxgoP7MhQZuLxapPij+OpfmnWWqFhaGT9XgeqqPvGhkPskWOXEEXrp4ZIk
dyTN5qWMUROYXwgOuERgr2IILVkpNMvxtSUntyCnAcdNZn5OzrV4J2BFr81DKw7rzvtk9FHYMc6N
lgjbXmMAzH3PtxhvDy1I8GSZfFN/LS6ryP03K5Mtl5S3rRORUc1LiBeKblj28NIXn5dQucliiSlG
PTHLD4vrm/Rb0ER//mT5tCo3oOkuw+wK/s5pzu8XiXGP5m0kE58FaucbXXEZlMe0C/PTzkt+9N0u
q7EWWBvExXITAekgtYAgCyw+aTZBz+C5Fb5deJcXmX1FH99hTwxyMr8hoEOljJzUwDAYD81oHRHx
9NWMU/VU1zmErEVLZe8hF4FwFZ7FFL3WVbnCBSVLH6XD2vBIDGIBEG0v+pBJcr4f2RbriOstKFCR
AAedKDDj32ysKoLC7I+qNioyFdT7X6h6MijwfPsE9a0utqmy555LwugI8rDIxvhkGgsiobhWQZgK
u1gxmOmm78DACeGGs1V6+J7mBhh563oyie8Ep26psbGLhSW01c1YPxv31gsn6BAdBz6GNmsoGim8
31gt0rdUfiLQCpEZpSW5JaAcZ66E7G3uHVql3cGbPk0G0LeUwBFDvkRnjmol/1Ma/IhiSOoHbL9F
kQ1ulWeJ6DCJDjb5asavAS9ybFeblZtech17mStt0J6IGlY+ev6GBgMSRhd4oif7pbPP9rNaguEE
yqX50YOx5WOn26UyBfmjgo/puOrvNcT51GgFHM9r8zIbBsPfvXjIphsXSTvCgzeS778oacpp/A3l
N+Uib4lbTJ5hTIcO/eNZn3zwiRYGHDf6kqP1PzVYTbXZHPXcPTX39yqjAsh9tfd+ae1mzQ3atsJ8
NECzhe07Y4ql5XGMMCke/GMosX+mB3zo1HMb7iY0XSBDEWo7h6OLEiOzFzcu21h4wC9dNSydWTKi
yHo7vm0KjPDOAOXelRjILJ6ISbzoq9ZZImsyUe5rou59xFazOgi32TVezZv66m6fVzmHOBKBky1o
9gqXZ/QdtKZWsvt+EAsmIO9xrZ+iQVu//EZ+J748x5mqF0yG7TBvRGp3XOHlGxnbo8E5eIlhx/tR
qxfHkyVJrM1LX7/oTJaoN8MWSM3QgO/9PCY8UrdCL/lw4mtbI5KvEn8/AEiq37i0TWTX9Px58wfX
DjzNErK0zBGAnKhF4UvbRat7/DpDGzsd8AxJfQPQuUOHyo51hm8MQH8dg6fy0IagRlpBZXb/xaM2
VWMeccB7aAvojLmDx9+272c1Dflv0VcBQ63CHGdm6a87u1gM8qFatkngVvxrkEzIXFOIZFBEUhjK
WSsal/xwA47irxwdPj43a8pJU5ymNTKnj+vFqzwORJ+5gg3muSR92WKWztJJgeUQpTRJQl8fT3L2
VXDBx5AJ6tZ4+QbKsqdTE8EpChAFWhw88x4EVL7Kqr1utACmULc8F210R9KeKWsnNNF/cUeEs/wt
h2ejkuU9YFLR+rrZFjxdk3+njpb90dh40tTaVbMoifZYFrz5wYEmcKjZyUPMOwrmf4CXxj9iAsOX
Vstl+YuNeUXhGOp0+ocE/iEyGXdshkG6TKxE4dgYTp2oxQeEe/BNzMnB6A0otXU/TVJUVZRNKY/9
RVF9xMj2ww0t1hWjAk9Wyu6XQ3qaBS+CPzuR2H7ikfCJWmfVXgEW2wGkmY/JbmN33aP/mwHmk2UX
z0V/EdPJk1HKmAvmAbUW3Cf9Q/3zq3XyMBfIUkdA6JBinsUaOAv8w+gzuCiO5/g7k73oU1QuMeky
U9EFn2mQB3OKFIIwO0/65f+itjtpJoyCFtuGGT/6j76YCKwq9qmNDEWZ5zkzil+E+VxKK2nblC0+
JklEaeqbO1lnyOGFfFqszodHw3jTRw6oB7+QPV+WTOFEjWDBnldVbMlsfWXb+FWT5OwdHLR2S6LA
LWaF3iR0AjM/4D2oOwci4o2LBS49fC+GBCQX8bIvW94AXGNZH1YxzcaGZ03Zi473RwZwmrP2ZMtK
F8yILmYD8dIKlsjB9FgSkM+xM8QAMcR9Tot/xHw+z+C3bzDKHBhHbgF+5uAlefGThqCLP8EUwXNp
4Jg5z1nuEr/vfAtNZNGdd9VkZ2uNbR17dEqXP0vO+qBl9qjBdE7ieHW4g5HTjl7yvpwb9+EG72A9
ZgHxIcGwuh9CqbUxecg9q6cCD7M3GubGX2nZq2630i+tqId2+IYrQEHMCNWVI7UP2c3RuYbZyPND
c56HzPbrNTJtV1Ik5Ebv2oooY00zHoVAm/nLZBNyXJVO5Txm9sOFTOg3NGQA/g5n+wJPYmXAIVnA
RMygmOomsKg7Guuc1Z2jtVXl5wIQHLZ0aR4cmcZy+dMWB3p2FzEtSAsP99M1ZnrUaJZuTWOkz8Ey
Hc28uCF7ynAe/vlT3SMDLnhqfigV5y7pkNLZV1by7w5AzlpqMHe5CaMo+xAqufwOPLp6UTONvTyF
l5pCQS/5qovAKmVZH9/6/S2QUoVRO0coLBDEm6Bu69wujIDA5GNKse4ONXL2ZguEnUfVYoFDUkCG
43OTH7UHOB7RDHPJjjPJQT1oGcwX0vY1Ag5bSa7hLnv43492ld64YGEcDeXCvuwrsFVbcdxySEdk
0RwK2K3knVE5F208jv1TIEHMaXANweFn48a1qioIBaZNyCVFn8MIhejKeGjgpZX4MloqiOs7bKfM
+nze7cDdeVQUIW4uE7shFPuT1KfWahLe/4hmO25JkcYm1GFccI31R83C3XXXBAEtvdq51vwmD8pk
AmLwptsE0Wwb0brrHSVmBzn1S8vWGawo5TADf3gO+KYFBSQj2KXe2Bv6g9T8u30G7TRP+uSp3afR
Ldu+MgFGTGjwYdtXf1z1QPZRYcv+K4U6oDCWl2mboNVniUUryq3tgFerOD6yz7GKIDpQ4wep0ycR
FijkHCzgouks26+kH+KC1WcXLACo0PzUHs5QgLTAe8A5fk7y9ogKR2mAfdcgDbdMtrtqcWOoZV0j
PLirfCEo9wRI5d0DMvyWHY5Yu56fggy4Ay81fRWhDRhf66zWCZQXJuq1Y+4O3BGiqVQPKG2KtL9M
gQHOiNXm8rs1iVUoaLVDPWNQxraAiLz4+RbGBHFtDn+JmWS35Oar/0iQYUgl9bwNo264jJcdX9W/
NMh5LWuOneFywJ4BAG0GW95XbpgOZjhUiZWDDCpVKoVRpg4cxmWZUtpTSpeSpDwiEih4/BfcO/TV
epGcwThJ4h3MX+xZuMp2KeC7u6t54DOEpHcd0Ka5H9lBIoJwkC+x1KvaObyuTkIj2tmjpGCRxyWR
X/5ZWFH4t5oQWJg0rpgkn9qPVcno58WC8laSmDhQby2vdQXlZRZXbO2gnoaYF8zX8B+ENEVxD9Sh
1MqMfldA88XwhLgIDVsJNtESanXZENljkH+jJlWF0TSYW0RrkUU+N9TUnkqymDRgENMG4jIUBUgf
W8gkgiDgv3nQS9kRixlKqiQqAkyAUa2a3qrsDN0GU6QLPsw+2MQ2Dr1usQPAbZB+PaPIMeV3wPnj
IxIjhTx35I3DI1y2AvmKkGuxikKEjH+mxmBKFyhXuFrpnc+ehmrTmGYGNEInYU85NPo+AS5rGA2I
kytaq9liaLtNBTr4IY35DA0V4iQLdG/9SmEtrX+b40jVkvvhNVhN6ZVhCj/HnuuYfFA5YBAwvPBK
EvfN/T8EsCWsGh0/6QJu8y5QjQSDWzzd+BPWf9vaE1ns35DQzueAWK/lDyzUybv6tZWG/xnyfkVJ
B8RDL4Wfs/hcgzLWXxrKVdgFIWx1hxyBr/T4bLY1IkjHwJYCkcMEDVUaGU45VvsmKItbksbgPI15
iPAKf676pq6dSXsv5+MZsLpay1bdFNT/NcmK0JZ3GWFDXeFO675tiKqvX/6sLEC+TRCH4SXxVekm
uEONOh87LWYQEgnujahma9iUMKqYz2RBC8/7/xr4cPu0/sZSHty676fY4dvNv9Mc50p8GiN/djOI
VkLbK/6gH8879Y9QxRNBddq1/WmDS61Czk/wwANnfGuD8GQIDsqBeKuI8ID7RqxhnOhyyB1ye3OY
ejhNcohpi/8jBIzcWPnmE8hsYD3dPv7v6eqCaTgVAYIcZ48GA28RJAofN2DR5JqeNrYJaUcBbGiD
mTmIPsOVDvE7C0CkRG8F4zCW/MOTTQdy3g2nAv/ZlbLNmQGFx1A0+TnaVFQVSIR7mdr+3TZvBBaK
Inp909g7LYXb8iH7O0toq4at4qYQVTCd27WVi2vK8UJbM2vO1x8YyVeAzmJQl5bk7T8uzg1adVtZ
ljdXnixAwkObyvDZJZqWsIety6yYTaQWy8mRy6rzwi2YRbZg9wVtY60QLVyENnX1C8riLND5lwU7
7hxxJapMsSudig1+6tyTO7CZ3SKkTo6O01GOMZWJiFjbcUQYprgr+Z5MQ6AnR8nmp6hd9wwKo94e
mh9uIp9p5cMqq2uDE7O2+qQ/OzkzU5T7sc1aTk5QjqwoIwcWe7nWj0aRQtBtTsfPYgbpalFODmDX
IamKDCtCJ37PgZMhkHmC0gvAQ8pW72CItLmJECpSRP6iMd0GH2/UzRyf3/6kuAFsqMnVB0YVhJXs
Y0lp0/GHjMeemfBRV4yP/b75ACcvIQPy2BUZgH+2xHOSihHVaakSJa1fCIJHViC/MeBju8YY7fiy
C+hqix68faCI8ouRShBMMUZaBU7/VuwPhSk4EsAnu+3q9UcNUdGMvl58o5j0+UUbQYeKTxXnZP7w
xNR7+kyyD/nR2SrMtX5Fal1XhBecKM5xEv2xeLMJrBRFgbUEg7zjxTg6YTX/3Loq3bAiYb0lfrw/
o4dtoY8DWOYpenAEon81Jl5SXu60k7dWAD3Rt40ktt0yhVO5SgbZU2dFyfcnGHZ+Cu1ATgqqSgQo
C8nVDQ37DHXB0aDVdpe6ucsnfUceAawIpMdksSz8bcuik2fBO52hKpMOg5W313Nxq3M2bf+RUe1Y
fW5w+0gXYwI8B5s7XBWx0ZoMWvX0JyL4jXL82U+/FP6CKDwQpZHnLmNUX4ayd5z1giHvSKDCnRfK
XEdPrDcS3uCo/EpMhW5eU+ePsjFJKegEtInTeVqgTonZsvhY6sOjS8weHr7/tZFRwxucrnwtOGPI
Hm65T+3muITgLXYvojDgxDvZupuD3VNwAxHswFtlGx1U16ICZ9j747v3bnXXNn1YTdWSQzqA0Xay
fhMySJd+kBf72l6CxKsmtuszBeXKCiK57MCc4XQ03BvfmgKkMDFXYd0nurvFbsEAvI9KXx/Xeisq
/3hcKNXfaL2fNvakfC/QSJ9wvacN7IPIgd6if+cj64CMvFDde83nTqW1k+zFYcR6qtfnT/EgiYMv
CPj+q/LDxCylmLLFKUPJZvvYo/WNK9wU6ngbewIFvgwHrkca+1bBtnjVhb7V0RUZSP0HntzEbxd4
aSxMy2nznSRzShf4zRKrUI6PTZphKO/gNECDx9SmJV6r4u1Xi9oNvu1LzgV8BSYderoiRkWFzfh2
wZXGqnLaUDiLlNBijAs3MxrSm05bDQb5j8ZrzPeSr4wMSTy08OFRevv3TUS3iqDZflka/YM0g368
FiNMDXPygb1f1sZx/fPiofgu18d0afG07eNjkk4sCTXMwZnzbzGWWwghcj4o+UaUZxg3w+OS+QAW
9ma0S6g7sgrhC/w1PMEw1uS8VwqWNBBi4PEWi6Q7sk84U/1v3wEuA0mKTwY2xZ3DyMUHwqFV2shj
7c8h8jNtnHh4QrWOtHXK/DQx1Vlvslu3VmQ8ZZCB1eSW4ecn8/6VfLNTvDHQnb4sew+UT9DXIa9S
7GEEnORqn5Oq5blXPwI8s+KLKdcBDbH70X8iPtcjWLtDkNedAPn+jP3qNRBHWLeb5IE5WRLnAKWd
iXB69dX0GnfeilHz+wKFaIdaNru6M/46cCRt1Z+Je49W6unPPRsmLLxIQPcnK7QmOgI+fH3ajrHH
yxYEw6v6Z0FROlmUrI7K9VWCm+0Y9hjOOB67xefrfglThq2/AyqDBydvQHnmmkGIsiwf42ymz5gD
AjTOP7Yj6+pRmiQHnKQSIWf2yzgek04U3gVrDCivM/szlgwf5WA3LOotJTjilceM/LqoJDz4gqZv
9f6pOlwkXMgOB+EoqUH6NaDsSbo+zHhbG1Ud3FBuX7oqTJTp7VUd1PmqGbQ06n1MO+f+p6DSpuHt
wuPlDGY1Jb53uqgL4J+JVVQ70JpUBeQhy1Z1UbUI4XIXPpVG2jJWjIqycLWh4eQOb6jzt0B0thu6
MfC1R8Nz5EP35iCALAj6ysGP7D+8wzhgaPWzoFEJB9BkDpQPn41LLZQRieu+klwh+ck8u5mg3S5v
3IHMqgu5mMeZ67GR+OR6ljDjfCDluOcKhvXNjTO0O0o1ICVuyqTFrvv+FlS+zAz0P9hdJNM7C5ma
9n44qzjUPKncjYtvEgn+vFUQJAXunDTVCGOUbjaM7WcsDEqx75zCzbPuLaJCdz9bqSBfnj5hESh1
6+mcj0HkThyJ1c2YxRY0iIPSv9BtU/DMbDKwCRVB56W0GVuskGxeEb309FK2S8+w94+PoWrayUh0
wolU32Tt9O1mliRnpduzDUX7118XRX3Oarnzl8y9+aK+lhxdBxWy3Z9/9r9HnTtCXSiThE5D1mkz
Sy+zUZHId2cvpQp+e/eShVEfSw9dn/Zx/+WkdvLOxkUoUXoEUnOfER+3Biaj6+qZ4V1EwwcmfM72
bt2nRDFgKW8BOFBE7NDgu7myyYSMFoDZ8wVMvIbHH1D106rePo074K4e31JhJOeZvtCWmFGPZbBI
fWpsJLe6UB/LF6fDnxT6ABNYS/p0TEXB5qi0TGUItVbo14bBNodnvsc9R7kuEPYh856s6LqPlEgJ
JIoE977PCd6rAX0mHBWbnQucDCd94YVgJsYqCpj4ghG1kct02cOK1hnzP1ZYcF1SPg1lYZFNConY
8hJ7hdK9ZyuEwJLFCHf2+p0TqIhYc2y9lfof4PNIpPX6If04eU3cS5xiHX1DCHE9uIT6QVSE3VDX
xfe9bgPNKnmfeXqfWFnFPckMdyeCZFq3x8MD/bgm3mKdUEv7c7olF5Asx+yFGwecEVofSvQQVkjq
qZysnYnLiu6ayySPp29XwNioYL4MNfdNHU6AVlxI1O465aSA2WanN9e/QaVVjoY7zymaDgJHWvD4
1X1fc+Td6j5o/cB8qYRVS2Jwr8sMNvvUmRG10EDXv5HXvDKrDQ9OPOewCuCPjGpZ/xY+nl/KDlXy
qQ5FXhZHqBfn6JD0BIEVnDXF6Ln4EebOlG2B6NUGlbbrCnz90iRkUfdIuGnJckr4cr4SP+hW9ord
hR9fD0pDGAqtDHq8ebsOczadCdx0bnd5pnWZRl040cufGent7+8ZLqU+seEeQ1m+GTftx3Cd0aHU
7HPHPhcp+l4YD8lp2GeutNHagp0HEGMnZ20eKCRzz5Jxleh8EuJBviimZ6HWhuXrD5qXhZ8TiASp
a/dLznRvdEi3Ynh3OAMxxm8WCuvqWno1xg6cCvcJ25WFN8fl6RrhOAVwmMSHOkLZZnFtR/BQGLQP
Uj4IJ7zGhSSquMWinoFYZXFnaHMqh2rR2d7M86LQLhnB0cl/ouTm5pAYqFmV+Mxh8Jl9hhkfz4pG
Ug3SPqCTUrRqpF0EcBavY2LEBRwzOoODyDi1uGIc7E4fZay970aEPKZzyxupnyYXAiiSzdGmxrZm
p1te2TBlW9sQwP6wTWUWNsHlsv6JYq0Zcx8MElHwA7gq4j2T8pvMfc7v/r3RrUvKola6P9HJqEDh
UwDPwju9/T7eBxL3qt//0y3G1OFLuob52/aWcRFGBwbwgQKLSTyHXNYWr2Z/PGPDQ9mXhEIl0elF
awSprEWEWaVR8Igk7vqJbrI8K+Kxai/OtxB6gdnbr7yFtW9mvvwiFZEwpU2CuUUK/oNRvpyIGKwH
TrMILTZmBAWmQM6ozH7GhSikMIO0CwuIjscnIftQPHsTK7i8j/LboUPS05wsKnm3d6Y9Qq8O/6mc
tuFOXJyz6Noin/caU3gk3keNgDu34b1jrXjtw724HarRyvVMgvH+LVVH/iGi4TxV9Fm4SJnkWDWC
cJSW7Tmd3+Im9vwGkc7Z5c3mutM7yJxgmPDAubjQDuza47ITDRhh9BsnKny6+yO1E1kNzL2BNvsA
9N+jMuIuYUH0Ky34+mEIil85HGaPkxIimS1ZNpH9JB4TzSkHZ4KFzqb4pMoT11izuU1U0IgxSf6o
1SgKLYhGqQPTBf0cDNmk+9ql7jg8T70AIwuN060oCuImNDZ11GesCWAOG/z7hVGwa/3O1IKywUmH
tnPvsuCyd+9FK/Z7YoaaqNT/gHk0OnfHIJ01ymriVUxkqBn8Nn2Sg2AYlmpicLMmVseHVdqIALdS
0Z9I2za+D6bB7/1j7ePSO/SDh4VmGp9NbdPtOA9vNIokvqMXlFuxFAcq0OYozDnWs6B4Nq0889s3
Pi7SbpGTZAMWkBFAcriChXPrDnoOU0cWZfgBKb9yGJLEqerldWSJdBF0wyXerBIugqF5Uwcf0zne
kjqb+1BKyi16KH++kE20GVpLQWN48rsaCZC2spTKgv83i9cR7JI3DHcrxbnwsFz/P67rEJbQTV8r
SBC+bsJEdHnyAqNGjufHUjtOIMbpV8/BjQ20gH8iwZlEiqUK76wHtFMEE+ONMjl+s37Q30UggVhg
IDo1u9konF9UUOL2dKYdi2xibBdzVOgTeXPDbqmaPucg36zwQXYoWYoZKE4rdb7+YJk/ix6A+bKU
zXNp2VMBQ/12rv+j8vxPTtVZhEs4JRrr9yscPg9f4ukH1nZaxZ+BNMdiF/cmmSV6yj+YSfTeViEb
KuaAIo916/NsPSoUtjCrqaq+9ZNGlarEbPQSVe4QgW95ltKSVi/i60F3tJD7A4fETZGVYgQrgG5i
EwCuqZgK8zxvOQXanIV+3spsrDwPaXYSY1saUmnDUdIGht6KYuMMlkdBIsSWN6oJg0TleQoYin7f
LaqfI8JaEo9p9tnvOgcmqljVNNoJCBBGbq0HwOWm89SeeDZUh9V22gnA4a5euSLOrJXcX8d1rOLG
nwVmZIXbqBBo4sQBDPJj+i76GevziE3xl618n6rQULfN+spVeDBc8sOqK1X7rzyU7dvxwx6IpNSc
KuobhSBo4zFmV/XMOO5DCPU/nVIoTd+uy9rnN1fOao2lYYuGf30fpDbITKSEE+pg2gAIYjtAqdIr
SbHNGAyssJt++A52clsSQ0f8QdyFRvHn3bwgE4j/gSe01kaqvk7NS+cR4QZMl/3sA8hZudJisZpe
ewTx4ERF+S/qhKk7esibKJPj9y7mzFqhKGjImeGXz+PcEaZEef1drMgQH124qKS0q0Kyd60tHzBg
c1VealK16dTexBaG5o3P47WN3/Zad4Y5Ee6onyRMN9ahd2QeGLecRiLzJRJOTw29/ZPtb+DN+nHG
WhlVkDJmr96OD9MDvC0UqpNNzTnmOgyPSaXuOyHJpSFWn7ZvQ0DK9lryVtBwaDY7HhSi1kYHX90w
nhduzwoK/f0Wpoei9FzkHSPJp/+4/DJ5SrQo4yF3iKGRVqCkg/XXhRJRJEMGLqoYLcxKnCtnVZma
BE690qZ4gyIqjcuv5XPpAc4rtLKRh0OBwO2aODljhUGFi5srx4vwHZahvw2UdCqZyiID/WCuMJSf
PKp8BMCYPE4LFD6cPlzh0/P3JuXiCz/eK/TN0slWG1bD/uFXNvI8vGd86yLxoXsCbV5vdllkYWbF
dF9MycYrFfpEgYF88Lh7yr9Kq4lFw/q4mTAyZDLUbMPvcX4rBpbWmsYCZkE21QUsB+omF8bSgXYE
jVJWzohXdj46VdR+JdN9D7VbJrYQ235OP5RTTBqSgnU/wWzfEwQnzyGpLfBEQfEAZ+YrN+I32DkB
mLwJNhl+CeWnjeXoiSrBG8mZvRGIajyfZpMWDPofwBRADVAFt75fj9jEiBGNoYIACkqjwa9EXt/s
2nrtojWVRXPwfiZE20rAfjlppup4snpRcKtlmobntr3gDgKHesVBWgOuMjODXpZFxWR3F7fYGRCk
p6ckFZtJjDEUE27bY1w7jWXooBS7vZ3Jc2Ifg64H6YsRMYHPOH+IzvJdXDVDyrbPQ0wvsveKyra/
P6a7AiKzRdAs4VTww1QltkpJs1DRHBK8Wc2UYFEb8OydzqZLm+E6U3Ka7iL3wsLeOl9Q53rOdpAu
mDtKGEl1GDGftQwAQSkCS7eZ/hbTQOsK+2tXK0z/DBRCZsPn7cCFppKD4hlnl+icGZyetsM8gdAo
9Pj7sIblBzztouUavrFT1usI24gkH8OT9rEVq5oia3C5u6LqIIGjK86flXIsdWyDq179eIVfK4+k
qGHuh0FD4NPZqugKGSZk1QX8bpr89tHTGEGvA7sn2VYSgqQnLaUrImKp8KKcZCaMXM1bT5lxy1F8
kYozSg0yXK9LIvHWO7g+VoZWIImApytKfLyRyNCGHENuRart1FDIrry77R+PwrHFXO6kpxCKAssf
E8ZKqsWL4rLje08ckQR7KzrXKrNKG4Jlx4wWpKKVaX+MwN2JgWziq0iowvaSay2pqxixelNxAdUs
m8S53lCT0+KI92Vkfc9rViDFn1PlEvm27XAtkbVV1ach6ZKcdIfuTulLZKJFeTAMQQUrPwV6XZjD
svdHLadUYqDLMr5imv1BAHIAGjbPt82rq1crAuUA3W4CuaDm86MGxUBJrOowMcSKVqrBAVPofE/S
52LiEYqRzlo7zxdWmL3IJ0AKqNSzJVnkql98Fo3zThWeNhIs7Cg7G2UdpOPwxvoUD60uVnpoCOq6
wEv25oMl93KjwRExpKhDWb+41qJ+SvBuzzoXlEEVbKJQ9xQLp+a87OQWFoL6CXo1LObpRKVdUE9u
9Eb0R/4Q/QSEEcwL4+17tIHataoSH9VvAWUKhpyL0Tk9XWQi82y9TcRzz1BeMh4atnLOXcebWGGe
CsiYdfmbtqDtHXykh6s+Ms74A1ulyPgf5HQH6KkHZ5IPRU2UlNPnVpiZ9yYvO4d4UuFoSRMaoH63
a9LDYK7b97S1de6oMghdmN6d/+cCqfOU8j3cSC8Thv2EeZ8BFa0rWHrH0T19r2oj4MdvzmRTAGXa
cpfefadX8JFoG9l58WhMzT2O8kaJynGFIu/rubedFNxgVjYKy1hQqqSY7j57q6r67jIYKE1bd0je
2MnlRVCXuRFe7oGMM9bDooGjGvpxE3P2kIbKnBy6lXjlhBD75HaG27XrNM20rs6uerb+Zw2azsqc
ezhcwQk1n9mnvaEUR3SVfUDN/kYy7FXo9FwZmGm5u75eGn3z/YD5unIZlmy9Y1tb49hJP473ZWDV
5MmsivlbjC3uDVWvcTuRudcYeMFzsa5PM36m524uIT1xpXPCOUUkHa3Sro0jkXosG0usLDbt7aNJ
vnSH2Z+QzIy4KIzwHbbjJz06X3sTP4NsZECcoD1MPcAvFpZgNhpB0RI2k8w2r9WdoyMbYZSj8F1p
LO9fnd1oso+/h2wzNdlBATvYlcZnxXf4tDBIisZex4PMflw+UFQs4JpsIeyKa1OuIE9gaYNgCcgJ
m2P9ltvUdz5snw3FuidAWNC/PlK+ywD5lePBVWGxyGdosZ6HrotGNXe4Emmi9+tcWyCTrLmFRCAG
aotHeY/QmxL6oux8oXQq1tMdTSeWOqV6H1tXcT7sAUEVLMyit0tdB/33+cTUcWIkcfkWmYevTD9K
MH6abRioFHPbMgnNuIdNdFkxX4/7yLMhdWY26v94HBV45FOOmJ6EX+sAK4cbswS4gJIP7Xm39jg5
ZGqosUNQn55WPAK0vdSl9AP9QPNoxSyV3fcZYSQcd0jZgNKF8IN30c/23lHTvp4ohHVWF+MEPTjM
reaTMqDmqLOes3qmXDS8Bgmf7Ct1rQNyRiWscwX7I05H6/tH/P4oDvr9glK1oXIJH6RSsrupE7vs
M1YRHShba/Ef+PEryHtGubkbCOivqFBOeLqiHc3AFuWoeQPCTx8Qdw6HYm0HOKWVODl9GL4XoAac
Cv7YBnHSjaYy/H3AM0joJRs2ZlA3dpMHGOyiTuaNoTTyGbWYAAgLRz3SNS91RCETk/2VTf96xWZu
RPPeSZ9G0Z6auVHCvt9if6hUUrypAesHo6jk//RmdeYqiHxH8rdUryinvlOfcdMk0l5p2Pu0KYNx
/OukxrMX4cN0WoRhYMA4VvF1+swauGhkzdng4bNLc8xBIgWSofJPfTUeyrwX1DDkK2LBuMkw5x+0
OV5KNmkW8k/EFhtIwstDlSurqSYUPYUfNKmCkreKfSgGKVih1HJczmAWGEEbiegpXl8WIsnMV+He
nLGE7x5IKpTy2/4RdHXxwXThq3UvJzyaWOSRemrXeWN8UWMxXSnrrjPaflMq+1k7gDZdSW9Dec5Y
Z9PqVK6dKczQp9lXa05EIMov0P5awTPTJ3/bQUiWC74UbaXWHS96VqaqRm3ou5DtF8XBMXTQHjZ1
qZ3zFtT13oXxrInUeT6IX/GFcxE8cyKwC8p4FSrRBEScLtbvvAQTarDlW6N5xD96QB5leb0y0Jwt
d1KFdFQ5jLM6kvM/ZJTJC3stzu4jCpWva11bPC7xtE2Xgn8QWbcbA1MTHbErHyG2HR9BeInaA3JV
QjI26W/+YH3qd1519u1D2IwRj98XjhpHWvxhVTtNQSvUtHqvjC+wgCvDMmJiSUGcqS85hM0leuLX
EBS9clS4KSgSKLRH2LEiQEMeAGtiMAdy0aA+/qlj+mVS1o1ISDLJLj5PjjK4+jqBte3/TNj327u+
5fr23Dv3t+02/vsHmJQ3pKAAAlPgyoYcYNuBoZmtsDErll/8gMqXrRV4JoNe6kVuMMLlVk18UhDW
DODEUP6xoDSZuFihwil3R+DjICc3pRrIQ9t6TcKPExU48ze0UBBnKy0/YofXso9O5/3TWSr7lXaS
KhIF6QcyIMCJ2+qdAHrepna8A46WPRSWWF9sYxZbqoX2RkSO1yO3Avmq0dZgZlnn6sCq8GwQVTZQ
SwMl/P+zpYQeHA/2qU64yVtKEvjn7rcbdVYnNxS4ZHRE8rHihVbV9ch+ej+cZUQSLdwvmIoi5rEk
08F+0QvqkZBq+MXxEdpaV5mTlrINgs+acvKMgGwISgT+VWWLwmBb7gwjf9uV7ts5eosA8sWKGDLL
qynkj8sulo0LDUweqIRpYn5kDyxf42APSbuqs74pBTlnlPvgOqP37a6ZbNoHMBcoTtpETikOvtkd
IKxzsC2AJqB4QjutIDjb3DYzrOvyNI1Ax5BOr5l+y8HYNuwOU0erSmdtEj1EP6dn38s9Lp1mwRQj
nBmsum+i6ZNFG2p7gL3GxKurPdggTNAtD3z+Jhv1dcYa+9UH9Q2sJPY460tP7fAef1O5ATZ6meC2
/VeCkLl/74qwUq5olK5Af0zTxAh9UfpltNxOEHffOunUE6nU2cfxNqPva7InlGOOWYn8OLBg8n+x
e+/edRJ+clyL6VIQj14KBCgx3Cd86V8uTAUwoopOIeFyMo1F5nf+NdArN5vdCmWirKk8H3V+Fo5A
JUqviyo8WgHAc4B2Cgt4acN1jaOU6dhkPssoc0ldUb8OSav+I2ylGjolSbAtE56jJKeLKn8oj3n5
ROWTS5BlaUAJhZ7gLST4UpGrrAzqGL0CD5pjhyiRU4AMudi3AsjDbo/TH+1cJp47h3rCkXwLIFBC
rJHV2vZ+F+2NrcCBVkdcEUUSiHuVjhxL3xsc3YZA0kPIMal0vtt51Dw6/9WnGDKd26yD4rmQl6V+
0SmiBkkAFq/j9SBE3wgoscO4xh+9sDDe0xbYkdqPwl4/pcgjERMCbWMQzHn5QGfK+m6tfwNOagr0
hxAMvW3CEcBDXuSg93Z8fUAN1vUx8yRVwcg/ySN+8HjrzctvtomfO8vwCTlfu/mZO5wLBlLtSpg1
4zM6xqo7tbl0mprMNkOwBikbWq2zX2PssXW/KTMm9WTds0iiDUk3bFwKzD++J9TDDrFi+HeoGSJm
v8uLAOh8dWEKoQsFhX2x0ImXVwEMgkTloez7m+US8VjF/BfoMT21QNC2p/0jJwaF+/1kYBvzHKe4
CtcAAEwyYE1rszVaXV+AOzZ/k2wZx87Mw9MSDCQDeiX5HNyhoZ9YktNPtTt/I19aBw7jcFXiTtZ+
do2/vwNe+2Ot5T8hlWCRSBHohKDxC4oPz1W7PZTYjTCF+UxxQXHzLWI5ihXXaQlVwKVrN8NsRoNr
ghTgceDMedhCbjCMFw819h/nz+5GVXftII2jghvYOduFBPUU1cjWr7D6Bq5ktPeXU/GcoVmtf/1R
830ITlQ0x2H23G5BK5shFbuS5yQxR2nqmwz284QpLeU+sz3VmzJPOMYT0cjfSO41WfFTiVI3tqGb
hQ23JFRgpg9Qjlwdt+R26L+EtpryG2TLA903O9wrIjfmZ0T4CGE1yP+wY4Yf/qb10jWU7is3YXII
94WAOa6BMkDFWe4Jx2RWMufMO+BCI7VaT42E6dqAJ5fqgDzPyti0rnTwap6wy+cqBvfgRUvi6Nrb
bYHxBof3hOKurUYjkzPHDyfvYx+F7CmQeTMaiK8VAyWJVvwYGLyghwbvIhGVu31Oe22WLK3j2ESC
tjLX41zkRijyiu0uNgUaVOJxnRCqdY591ZWdRmfNKcTtcW3J5h7XrPbVvKkhqpJnIRinAv804jd5
mnB7/0b/xci88O/5cTM7bOIFzcT+TtoKY9uYl6tD7CE/fcLbf8teiSdLF9da/lLTskwM8Oa+zQpk
ZeT4cd1u8JoCSVABmh8wwWlHqU5XNRu/fjhnQ3MBbZXXdn1oYm31OhwvrYlvOc0MOYQWNqeTSNYu
XQ0CZxsec3QKBOJxEO87NwOlELUNJfxqi9Uan6qxBbnZF1dz+AVcjQFJMOOgsOzkyil/ng/lz7KY
DVfvAIUxuvX7YEsg+y0sKKmj72FbK1CPRTEj7LfAF9tmtvK9qR5YyMguwjTiNU9TNntTnh5nzS7d
Kc576GCNsVF1qmoNT1uWn2OY9XYyC81kDRateKf8UOIdqZ7RWsbqWqwr8KTvNWegD6CPMmno5N81
NA0hIFkdikagdHHr8XKIZuiYvAsuythD1w7jB8+Az5WRXoRwhXYUV20dCFN3PL29vSW+kH07Mrsm
B5/Mu1alnvsZO4QoC+e7akhiGmr2hOsCKxIM/TMVEImIg+6mTtjVmuw5YrzdPXwGtqUCP/au8fh0
QxEGrvjqQ+wZKyOIjoHw8wgcAr1TFVOEo+1dCL7iKTVgw6XsmKHcpLKDqZ0JDFw2sAkuKDdP3zLe
RRDFKDsBGcZe+Igow3gG7g9S5IYSBYNFhkcGpg0bLru4wxQ5PHJsTyu9lhuG0F+/4IfjrmVljj2/
fn8BzxZ0v+U7GiEREXQV+ph7ic7RxHmswqQZbmihcN2sg4AbSBQ2go4QzeKAwPtLlyLsxS99R6/O
mr/n8G89fcoCrnxnuZgdAG3isseykjHvh24/itMmfLLmzG/jwXXJsFUAT/iNqZ2Tg6HIIzxLmMEI
cuKrY9dhBIKPMXJuolp/Esxt3ldYn8TJucVMZF2I8xPWIkca1ZSCbPkDkXXE+iUGYaKHlcjsA/jE
w6o8B6WUAvynwL0UMZAh/lCBJH07/JMMsmlqhoQWcwagySEVywMdRh0NpnMI2qExbDVzw5iuMoPw
8UV0coXuw82eEbiKZwMFaiPeAUFOmi/yGvtf4+S7M3newDqp6EfXV5TCGl6nB3TOhkTqyONr045q
KSFgXiWEWZveDtOYV4CnMU/EhAxgP6Fjm4ndrS1qI8nUBd0MDFiAdItA7Sd42NmoZ/Mr5YNXysHi
Qfm1BnrbqgT3B/VgDu80wBFgZLa56DPZZla8jvhCahAKM8DujD04J4JOV6N8hVWXkoRm/VcFQuGu
D7TIbfx9YG5OUMpdSWh/sZnkAR3awRQJmlyguLfzxCQhAmE6ClKVXX5bQtJxmeazAV1B96hkEDjm
vWIYhROJQ8Ms2cTaFSgufJyzQwk+ITnNUIAPES1oO/Hd151UOW8ZcvWwJCmnDLo3xOrEfzpFxZP5
I1/GguATVWX4whN/uow/JehK1QnuQJYFbCJlzaBzNvV97XiT2mxtm7UAErT+aar3Ggt1oiCFE2+3
ZHaAKZ9eXChjly/a4bOk8JoMPko1vt1CI/eJBaeBB6MJsga+rCLbpRghByT4WTKcbglQ3IcH8V0b
hEtrveNM8ZEF5J0MUs3SqVITqlhZqqE6ppWOb13gRrLBRQrfwWGCB2fOjBbxL6O/dSR5l35CLl0o
noznrvg5RwVkLbG/I9JhWWBJO7hfqpXr3BIH4PsjdVgvid+JrhQDrb/mUUVaiBpwVL9DcrmKIhsh
9sxtI8fHbb7T9Oh4eol+sbFf0Qv5PyrR8uHueO1r2ySZfntzVSFGoXpPkND8Ij3tgYvJlQaYAlxx
HBgQULKoOdNs31imwWbLY0pkDU/T1M5GN1qRrIm0RvFius2/r83WCVLPcUa4GBeAxpxxJpOWEYtY
YkGEON22yLJx52Rhdi48m3QWJPWUtXgrMeDBcijg+vddzaZ9HRS+jluRX1ue2rMlmcnPzHYfd6Hx
JB3V6ntqQPuWRIwKFvTp7PfPK69PEFHn8TQd9JRX0mNEM2j3OaPkEo6G/UMJxDgsa+x1r1o/4glX
91Huhl05EFO+NslmzCm6z0M1t1sIKG+Xj+Xu0XO+J6Wean/+mSCuc7e/2VY61Br5O7wuB2pkVILt
3jAGaJS0R3yzWvovK3amwG1JQ3WIQgImC2AVweeSNwco0pdXBdumcIPWUrzy2Hb09iOWZc3xYEjo
pfVJLWJ5v85c+DDLuwc3Q9Yn80opQ0iHneGWPwtub8cIIZ+0WeKOzVaiJgWL8PN5hylqQq+HVypj
eABSMVhX9pUKokC8QBgo8vNJYIWaP7s0lLjdW3xTwMg2r7n78+wg0sVb3MXyDylqd5Xt0SZWdtMA
LCbJzRE6JlHKbtYGKSapVOF7yXL2CWjKQ8q0RAXVvYjluLVb/DUI1hXyeGWjVqy1p2cg/4q4yUat
ltCHYT9XfQPC6P8Ch/4fq6UcZSX/08bzO8dvqBfeQFwH/gFO5MedeM52I3MHqyPsXUjObkIIU2LL
u910I2jpd6HGO+Cse8h4ZnctGqlcMadnPHQG2nJRDTiM8hO+c/Rutjs1R30zFRQMzlhk5CSURiOL
7ep2PeRkqjfisLxat/esHOdEo6EIvkBOIp5yomOJr5RXbz0OTnZvlgyMKYRltjFOGDhNstNF93WR
K/W2bvoV+xIPpAadvY1kkieCI6AgnDFEYEnxuORT4Ij4SVxZmtvwDMbFXSWB+qqwUW99g7hmE9nB
BRjpLOBPgpxWglvcovJgIlI3GskmW1DEqSXN2tBBxDcbDPzvKHlpzD0uj9JKOMb0OaAiCEL/1Vi1
PdqsNtVYZVaUo6qsX4Pc7rKCgl0a635LQrSgmslbQ18yM9bD6/TbVByp15YaEX7Fj54V9jRyUNcu
anMLjaWoQdwgcrLVkbt5pB0E66WsVKk6vJ8V5tX638CsOsDdE/stJwg2SqGrHbO4SuxmXQjPVs/j
Mrcm9Aoa/5yw3pUgkcs6osIY3qye92/PEkL9ywcKNaC0IYtxSuQyZJvzbpMCgcoclJdviv5ao6MX
B2Ekw3wGC5JNOLlx/4ktuAVqKx/OWvd7TFTRGd8DkuouJY2tFBoTZ615CgZl/YzBzs5z2+R23K24
qX27rj4jGqDYN0Tpootltjk19rCJoAWJ/GC6jUU9IwIlrJgKjXHVpgNkM24jZXDPC/x17Chd3bVj
qElLMF09E/GR4EduQbeJGirf6RD08weyrfzTFAKMfQvHQRhiUzLkLBk28NJR+2NLFEOlQCRX/iU6
YBcjXUfjWSuGu7GzZKeNnLQyG7aCJjJ5VM8H9Mu+rhdgr4dm36Eybse05LW3qTbQ/cf0RWWxP3Ba
pzXRiOys5v1bQ+sefSS47YJFju5yghuWzlDEocxH+FNcAj+YM3U6cE0ExMQN0oYXtdE7ctiHeQJ8
gwpC7dsTiomua1FCVt4RhhsehoQ+hsCDsUjyFD9e6vHM16W6M0Prlt9WCiUAzRiB3KtT4IGqGLQF
RSFcTW19WhXzqtXHhxIXeFKgqtsfyuZ7Z3OhkmfEG9F7on+26a3MBY4K9Ne35XFRzQXU7LAfop5J
H/U0z4WF2dQvZsg45bp1uar8yDSSr6fL84WxqPQwMUfdJ4vQojnvwxqy7XWvxCpw3YHGUgr22s1s
qfCLLlYJivlBnVBuZxc+WXXIjjO/8DW4FJhJCwSrKR4VKJEDUTDUI8dJbkGgoSBp7SqBGiobfvTO
ZoWsQJoqAZATsUzRNzipmdwU9tPuPCIcdN0x9r9m3hGfCtmSPtaqfh7ZA+T23JvIRuu3bqj4joCB
fB+2/o4pLUfENh/169fFVyGkjkI1BGOOv6e2oqdxvsApGfmY0Kd/C9T+uqrYyAHZCZoFYIYIjRlN
48ZltdibqKIJ7c2vYrgHaLla3RAkQV6y4Ax1AaBbAAnkMHYVbjx/cYJPXM5Qi1H7Sx/d/7cMcQs6
yI455e0g4sJUlVKXYzz1ONy7t3UAEMqjbXEoXqWkhRzHXfB4fSkQNvJQuYv5m0UwSZm98cI084SS
8/TuS/ra1X6zuN7zk3Cf4ClbfYH73P1oWC7LrtW1EeMD+jUnwmnLlc5a/HPD4U0ge47QAhlaN0Vn
bR4EkBiFqRgCGqJvgc6SM5CPuod6gYE2v+FmomH4a2rCqBbSGBkRMC8ydPE02GJXEXa9Xtkd9B+p
XKW0AWDhLsV9+A8m3G9ZkQ06/1sFFJGZ2Nf6ijob+1z4moOQLa+2VznOQq8ozwZdzfyw1XRxeKme
1PKQPw4ejVriP/6YNhjYM3jOxGkVWhTcqzRyOOTqmSYE8RAcqx7Nd3JG+S+ksDoJ1T3iUubu/dJD
4IigT4DqG6dSJ9UDVmEraOFlYtTfdf41zo8OUzFWpoyO5YR+Ns3f77MilPPTC8vojIWA59bTV6gJ
j6zwE+W1SJvz4hJ9jXOnwLp9w9CufzhnP9fulbc3pyXfVx0jNWLevhADFRKgMt8wEROSROPFBldv
9GzpCdYXUTNc+DZUCeH6jz7JHuPxNbSY+JLIgPqW5OR1PVGi1OBx2tCm1YYsdhNyWlLKVfnYcqcq
asXyklfEbwBeuR87o8pJJY5KAOdRWHJFSTTdhCyEVnpzqENYAgdTrLkb7QezFflaTl/ZdCSKcODm
n3B/nDW31Ktms4WYbefjGeMnGNMQYJ0w0ABQETrcOi9I1XgwsKVrrGzNuuuaKgNKcN1awG0s3cnk
CMa5Rq0L6AA9Ijn/KKmqwyuo6T0AAYo/+iV6Eadllc5yGAnHCAeZ6h0K0F2Aq/pBeTXwo0+Er+Ws
dCZ4ZI/aVsQvGNtW2cHAumZd0SBXqePeTcevcT3KQ5cVLXs+gUMZFfqjjTPhygtJD+SndF3T18zR
d55tlHqMSv9MVNXht0BgVYaZdq5cohJJmJRrtTFk4W9ZZuZWOanWEvhbg+mccO1g55nYxj4LKNem
0ctnoIQppoquQ9dl1KLziO29W+zWT4dUXkFK2tuCqG/pYLd43B8hNvBzwj9iaMTogAqb5YecA7A5
vaAJwUw1MJwvCdPE9JIfVpmYqbf89YfrWksQEp43M34PmS0bZDhKopYsV0SDLj948C8a+uw8qWIl
ya2nJJF6xGwNdWV0PXfHdOzB87vyHyFsATZTkww6Fi+6YwtGa79LH5T/FApb3uCKVjR45geIXwNk
sA1DK8CGvkEww1tOLQ7/vBpAyo93cSZIcUdSwHEBQdhw+28yzxDBHnlGnlLuMf9d/gjHmbZ4xnLj
QeYoPAaXV1Ti+tYjFrl+NNMrnkoujyAtJETJcgRYwgmw3LVTDOp/n8/zrWOzhrqP5ifJ6EtG9wnq
VjMh91wkqhrJ3Ix2UrhzBRDnOyWcaPMmtrOBnGKcdehIsg3nv5v5dxGhxeuAcKM/YUbYEGKFZPsb
HzPEUYJMg2OsKGpq4HXazZ/InU9jwWEqf1lL6AtEKsa36IB0PFyIjJmanzD1scyJYK/AXUAny4d4
TmOPNINIZ60fWblsSF63de8HFF6HgvdP7yjeDBvmr14gjYjKqsYB7e9GaO5QD0PeqXnkKGQBIpLw
7/IF73N4eoCHZexjlrlrrGls4eWkzNnM3TVhFATlZLfnPB+nCGu+AjGjefKyQX0GFhXyD3GbXzCW
dRFoLdUPFz97Zee5OM3GWm8O2XtiypIpYvU1OaBPrpG0Pj/x4H+3MPzQgBPth1ia1JW+0TqMLGNP
RZ2btWE/LKvTlUnaCyu4vVbWhsMgykvtVdjyQkkUh/mn/V4YYWLkTwV8lh6hwCMjTM0RuQdnnoUx
zPh8jxU6OWxclzPh2nskt2rCaOzw3wSX8yBc14AD76McIpt+vgNWpYF9ESliINM1goZasuAhVNS8
SxKSSv4IrMTxxAJX8LZNvK+gNxVO9vJpFMHF/6lwhwZibY/SmcqWFkXFNAXV0WqOwx/YBGts5oZG
OCQ7PUEHOyUwo5TWD2/RSN2yHjtHJgS6rvcuOh/mK+iqjresXYR1eclA5mZeA69gArUht4JcqIEx
4Gbb6YCddZdKoVFPzJY0Q/m24kYD7NesIgo4mMW6PXLX6OS1AR/KbrIoTpqIFbwUEYE/OJaM97Hw
okL2pHWuu9TZgG4eAkY3zt4qxwUwNF0LKasq3GUokZIEPcAqdeU9Gp8jOuSGTTqgppHs575Vc1eU
iMWT3PIjYfg+f+3RNGNjHg5yNMBwA6pDoONwwIE9qCSkuSj4iCzIi4/Gr+4mvzZoB6wZtH/1mIBH
DJsORFR4+9dlPtk0dxiIWT2ZM8u57DG9vTgH5iybVHydVP/FwCBoTkjY1yM0MRN2ZrKKXKoRabvX
xFl3gi9KiqlGnCIv61hRbImZ/5/niCxIMt7YyGrM6HpG7gKtJP7alhFKmODxsxxIkuxSn+0geqDC
6hbmf5KC3qGrSMiz+JwKifTxqNsu9aXgzDBkG7r9un0/obL+qYkVky9bYfLIcajYvEb9QdxH1Wvs
ZFsz+gSsY73T0njF89a8femwgV4CDHyl+aJP2kpavhDwjKxzXW8Kp4UGP36aYmMONprSBk9o8h91
tQXE/7n0+odme6WelbaHiAJlaCO/zFqaINaJVl5pAG0RqgWGuUlgLXrJ8Gd1im7didWeLyVf4CdP
+4biIuabSISKpjS/PHFEbeerY+xHSpDtyM6YTG6mZvXb7x49SrdtZhG43ahJA2c0Tr+oG1MeCDA3
l/A9fPntNzTodf4hJzmrnDp6NWbG/HIrx/rjz72+kmmQMK0wWer8EQPEqkn6CpG6y3a3dSwhlKTk
b4jmh1m44i87IEJzS4/VeCLXY2ge9hvSJa+vJKUcAicXDC2cuQn+rU8kFz5jFWaADq3Fn1VnZNfQ
5FcJhSzsqZwclH8ZEoo1kXF2Zt0uzFcU2ILV2XWPkw/ypCLqwi8WJ30lbhgvnYejaditcJGl9DeK
N4f/lbj+hQ2V1ff1mFThTIvIQivVxlHT6yGCCWIlRDUqt859fd819R0wjRnUff8UiI14ZYefUSy7
6UH5lJVjS2i8SrF7Fw4njCSu2gsueFCRs3PGvKU5Gb4n5WtL7V+Ky5yQa4L1sbo28X6zfJQXx9Kt
GItTHQ8Vv+sLrMf7x7jW+XTIycsJOB6mh0A0N1UE5fi7wChbQdb3ygVv0byZlI3GxMW3s+HKZ+RN
uJnRdZkvdylBN9WmmAYkF68eCHNFuTZdSAlPkEXhigNg0dZWr19hiNLok+L4OD+uBuYxmOwRzgVA
hPKej3uPWK9/1rbeiybaJfYF1PHXLfiqEEUAm09giPpqBEINXVxdwDAeCAH/UPdeUHKKAMkBmzJC
0v/9/tPGn+ndPbUY0XeQC36rWW+f+kfRuBlNC1hQmGpcXNvnjWIgQCpnHxkj5O5jzwmGG2EEt7B4
J9SzzBBXAAaeeN6fs7tgnHE4xwixGoXoMaKYrPX/surbpg8WOOiFSeHxO/74PNLN5TbfvpwMp4VU
KuEfxuuSAJ2X2PXbAyQznA6qC0n+Tw5pwHneq4W9DmfcWK8SgRLJ61ZI5cTzT5FY4U6nFt8FN8Cs
InQj9DkmnBNGKj4y3ftKOpl7eTZ5WBZ+GAvv0GrItR+ZBO+HPuG41ar+lvb1VhZptInktseI0xOn
9poafHXnVdaIw3WhROdPJNoVHqeHKUPBycBvMbSh3ffJNpJQChxgy8q+D32b0rvMM/IlYCL5ylv+
haAtHvhirT6tTxSWatPByT3rZ8kNfkJFZLzwudSnqQKi+3YB7ASPcNy3+U0NMQ3R3xxMcEiaapg6
KlukYABVbc6C/hyLsIQDBcMiEIT36dAw3pxL7zwDi5GbwGsC+NVbsVl5opv2BdTDEW2m2MwAw4At
wP2Mz9KwmcTWc2WPwuga+2Nrg7X3kWRKsS/DCE6B7FImH732Fk3fVHWSCiVF3JRUAUqUAOmH4p2j
eLz3ANztyAQrv3tHTGSec6/H9kWnRxmH6kvIbmyAugvfuk1RdNa9FU69VVWqc4wAtLsbcd59Rtp8
yjnd4yRz4oPQN25zl1p0LqWSZ1OT+aZPp2xTyGAKNGI4FtJMbVnlyJHOZbMDl5l4xx8KTHDi7J7i
kC/yyDIbI6Jgc00vdu1h+CvK+tiYOglDZ//yTlyB66CrlvT9OGg66WQBfRSuWKUBNvFrEfDGExvA
Dk0rJ13K0bkm+V7t0EPIumEFoxv7IT5OM4NGhD/41OOgp4+WFCnEKTIdN0yCsPAlYpXztfceEQ0E
kmz++WEPpWW6WT2dTF7QNevSoRbjlh3vPkP0Yd5+cqKpmhVeuFUTvrJj2qe1LTacUeJHyXxIYNTL
KKQPe8DE5U702K7oruSAnxVWYbaj0vMTzRy1IXQVLtgp/ERmIL477UMVA4uWPB30O4C/bOZAEZkt
84coXorhsEgYAQ3letYcxB+MDKm6WXGbtQmaQo/pCTG6PmojwNkJT1COdHnQCno70vObdvMarzCg
T2cjRlb/Q2C0XS5uCh5QS2s9z2fxGlJH1VH1VZLVG8NTsHJoXE79KM0eGuWcPkaGkWrscummiQyr
zBYHeDxnEHtuuerGFFjYfl5auspL6WQfnYrldGcmjsOdEG7DakkDicZHo6gbdk4fwmB84O1ygDNZ
0t553r5wMGAY1nUFTkOMtGon/BtlbOUmAJedOW+FRYoE99F225jBrAZzshBVRerByZbcZQo4NYPh
093UqnaA9MG1iBQrlv42XRTZ7wsV+WDBGOJ/V3tfUUTiZZB+ml8O+fXdwk0F2lZTKgYnd6aWtSrE
EnDKwdjotnlCeAwtWB2jrq/zlYeEulcPUzYfyziNvutE8gIuQ79pVbnEt3hHgIbo7mZoA2QtBBLS
5WPGgVCmyRElkUSQuBSzrb8arx24gKs0N0OAM0ylj8fkQMjyJjU2/VveO6QzF4TOIb0zYNCU2u/W
pElSXKHSCBgUp807JKQq9UKaL4oJlh1OmUNNFOxLNTBvyDseZNMvjojP3PpY+PTQjhIJZLfzF9xB
GpMcYoAbi2MpxI5xt5/7NG+u91RWkL7aX7dZs/8fqx0R9tBDg5HRtRSYEOhDQHy9sn/BzewJFUQ9
16jBMyY1wsXwDl6L/eVCg92/CkgVE7cOJbLvxAfyNjBTHuaQ3bdt2OEDcf+kCOzNqr/u+KCnABCV
APiGWLj+1X+J6uDJ7haceDqpnR6uKM/izhjC5DhA7fzhpQm5axpeQJeZhR2Z5ERIdenX/2YI0qnu
vUtMTplQL6WUgWIWNBCmnoIACBVEQN6/pFtuB7gC5d5xUjsL66ZRUMkxLfWWORdS8RKNZcNEapAX
u0BCVmj0c3RQdruGlGdKyrkdzNtxpozd6Uxrcpvztnf+T1xN/vdfXChAsBDaOyK1uTTWg3stfaym
LgcWfwT4biqq6/tCMUs297VtC+1Cz2HaWccq/2jMaQBiRsvo5c9v6jTcOJwkMNVEEAeqD27MApWr
QYlq2YYQzCnR3dbfz2LI0/RzLHYygK1KkDOW1zk/LLdBUZuoqq9laiObrWScfJXFOlYWEAYR0+bl
ILZWH12D3wtJAzMsSWhHCDsC/LeYWYozaeWQjdZx3SttkVp8eKgKmEOK65VH+K6Y4smzZ/tkDfFM
s2G8ZarqD5TFgFsES7nsvgLSuFwJIFWINamso3KIFIMjRObxTLE4+cJYlPSbaXhkVmC+Dp8VSoXM
HqahPFeT2H71uktB9ZB42L2vhafNrRbhLwa+wZcTR0GFAJmMaW/zLMnoWHbn53olydVFUpLE6SNL
NSeeUCvFDehBibK8u38JMPXA3KZoLYe5qXTMqqXQXNAIP4wEVDZb2YuXGIstVS1z4Mn+7YeIEKmZ
01BfKP+DcCVa9Qzg0PAdksptXmo0tvyQ7l8FOxcT80wthd6W1Qpg3ha4RJjZeLUBaD33d6iifIlb
vyKJKLV3F5CNL1HgLdhFrXHnklKjhfgh/tqLZxD8qE4STCGZdU34Ujs5F+hr7E6bSg3/bPxkRhpq
0SFjuqoy/PqYQliXXFiX5y9/Rd4QkCPvEO4Sra+vyLlW3Kzx8KmRMr1tVvaeIqhj9JOEL2t16nCA
kH8JEBRUBhsK6LQkKCjAKm6FiqjTBCjcMhP2j9LfMdVtmxSIvINS3bX9VwokB8TJDe2ZsR4Px6xs
KTaJUBQfqKhFVUfYo1vktLyu20jMib8oS6VrKYB91ozdsMoZK6MjooM6z75z7cicBpnZqvnqStBw
jw080BbWKMdRIjr9Y8MgRaM3V49hFt/v+i2fwEmMZNUJyI7XF81nsaLu6s+h7B9kfcFuVCFRuDWw
K4LXxqeC+8wg/C9ufET40GW6rqlIxEhqUd3eXgBlN6inbnBztMBF2ivTVKJr/UCeRXrA30x1ThvJ
9q7tUG98tvSL4CMsdzeVZ6UMyXNdKeSibNm5KCxkcVflB8rKHDgsecrIcnx+P6a1SOmwoxh3zwNp
Mt0BAFesGMyUEe8kdaTy/nLQLY9u/HU/n2GJzoNGELpk3ohE11kmxV2OSzlWEJmStoucj2tt3dtK
4wXbXe9FFxBqFkiCLzuCzy04pn8EgiMEt1ErhQHRra4HD2kF7gSyY1WvE1xhdk2mE20DhQq8FPgc
sza+P0cXZsVj4Lf577+M8P0cUaRThNdjflS40Tt3ET3hJH7KYStmuqwt0c/RYW3hHxy1hI/wSXeV
5XXvJ4JR1a2eEnLBKIQ/mk5JGgXg9neUMgHPafkpQC63V1WkTn9C/F6qiRGV0/8r+7QpUCOtqYN9
0U7hb/3Dlp0EYx7BBvv5y1GEl40l5gAP52ebKMPJAdyQ2JSYQjRNBWukpyp7MXYSMuzDmkEGPhWS
gHMCtWenEzfiWAC2htq+RQv5q1bCBrTCe3xzHA97d/YnjCLHh1N8Ish5JNwnOYS0zre56IGorVQ8
ADcpepRMcpbhoZkU6igjYfZu+ofjab1jw5J/5hlldfX1zuKT4DHnHJhrbet9bxB+VkzYPXxtD9xk
JIdh/WM9RH2shvaqrPOBK/2jAqft0PLrcFbZ87dP1eeSPxxlxUgcbxafW60ju9P0ufWwBt1pa+yv
8SuskEhNsSvlzRl1/y/E99ZLtXN+Nb/ZhC/UJuM9Ga7uvAbvpCl1q3gGDtIi+qvFvjjJDEbmDCu5
qAVWM04d84RCCIxDfwoZNhKvd8BxuLrrP2CCQJvRXepwlh0P/U8VRFkn7GjtNRv/tQUXxouPiQwv
Rsq4i3ByXkAc896y6tVCjiQsrC2cjRFL05HHreAERTk1YVzpFXJUrtPq1tnWIxlmauSucHUtZCer
GhvbIhb7b8932D/IjniqNYkIzBGexF26ZWsObSQDNf/GzcEoQrwT//AT5sMDnv8MkKlOI1yVmAB+
b1dNmIbeM2Ucc2HzlOpDWa146AxmTl4G6XsTi/PBhYIMnZaYdNKGNLr+7bvH83uv4j+RvRlh+mNB
UhIvnb5GJpAPDZowcgX5I/7N3nhae+HllxwnWsoiOXb70NUblyd4/SwC5oqDbYn7k6ywntutGR6L
+ZO++SnRgZi5rLe3j/II5cZ8INlhacU4OEEobbP2QO0/D07djD93vnDDjjAXlDytClmJBsWiUVQw
eM5gwdtu+7pTgK/wTJg7HBWBv/bcQoCa59btMtSmFtcuJswRxiD/8Lj1UvYyD1qEheVmOaTZf8qW
LoGPeCiozF9vZYVnDgO5bn1gx/Wkdmf3EniqimpYo56wirdrBPmUa8yiSY0rxylte2qoGfu6RLXx
SUL5CCoiLF9H7nip7ayufbKpxNtpA0WWIJZRQRsFDjv7ym6HmdYD5jMK1qlFgxT1ehUt6CiEfTcz
MDjgmnKztMRRdc1FwytlHV6uaB0+fE+7FYbXx5XH1pjA7CH7WrZbyPE+9rQeOUrlpCHhm5zA3CKn
V2WUoCunyUUEuWRWBhF6HmJH4lZRitNBbBAA3Wt1O4Dm9CEIVfi2t8uidiAwKDWK53NbRHLkGuaH
g5+c9jt/D5W7SuoVjHC9BYqkUDqhA4mJ0hXkbwJLWU3tqoz/70hN/yg96CgRCUvtSB0CLmmsJpQj
m9cpv+F0dfMDxYO/xMTkTnreeEUMkFHJyRfeRPONv9DqrBSYc3NiRor7Wsu0yF9JGuFcf8W0NOeG
14Lmy2aebiwG+LAhXOU4IxHjBQ+pX+iv7VvtVl5xZCQovIGYYcX3xChvi2tr3DU/IOSYfKnPkfG6
j772ys05m7hYp1XW8kCykPBeqW/+D+ftKx8EIDAZczY3kmwSSHp3Keh3/pQT3vKMbHCYAbDp+0H/
UaQA/igHBxtl8SKu4QuUskJ0Z9DqTxrh44wD/1NZ2ckIcD943hafMB+Eb3ptgi56DT+uA2g2ydYV
fCBqFR5Qm2LxyOrn27PLoOSjppjArTGinRRUvfA5V99CGpSO6K2JePtqG/A4Kq4sj+7KgWnuZUOk
zyh6dVgZBGlEqzSBpmyqvtBFh5sGwb8IiKIvjclJynvg78Xub7GNgEp5ly96PwMdv7+ovP26NaJ5
UuqDzkv2aLSOqPgzy2sXO/rUapNgENelO2f3sJiWL1HRQ6XMSdzKr9RrQveoUsjowkxrPvb+JbGn
ERXf6LgbuIGvpDIZHtdC0EgLqPMoYmO6iOJ964sYV2QPcv1vHb/t9Gskmwv+ZO67PtPZaJsJe4XK
KcUZNQoWt7DRMbDjn1OtPvp7sLXSqHI5Ms2KiC2c0aDmWcefOQ3TT1qD64RU7inklw240ZisYK+M
SS1mNLo67YwflgXEP1HwdIp94hRERxRuKqDVVTEcmblJ+spPKe91Hzz0eWUkxS0RV9WSFdC2gRSm
xxUP9xV0yUXkvcREwwHtTmXe0f0aqHRESIBABFH263Snl1dG/HP26rVYVC5P5d8qRjJISUoc6pbL
M0kF5KPKV0dzTChDNEIPKOfvE84BauvNfm/VPs/r6dn513sH2f5An6f19K3KrexSP/ly4qx0FTNL
Gu0sOKYEwJaOGxDuJojTHlYWYrTEKWhLJB+WgZICUqu5zvp9Wki4pmVtWNR0tXOD1wIdTyo3PGzk
P01YrV/a7JKc+Mbx2QgO3VrWyqFHNOR1ClhLSQ0qBcruA6IyKICkp4HNMWFPWhxsYmeSMomuGPIM
Wj43tfDB6J2TgYaSL4HUD+bdV5adtLeMdsg6lVsO3u+D5XAW/ToE5nSnO0spS7ClhDL6OZvu8dmc
551UTuFdgpv4W/Ub5Dd95WaaQAJhIaMbNva1fxb4r9/BWHR1QvMUqoH7j41zmhxh3bxr/4478v+I
zu6cdokAkdNGcStAzc469V6DvJeTuwfDkOdGadxHsIEjXaSIM5U+lrlvsGXJfrCVXIOusS87t/h3
GP1IxZ7+yFPHjRms6w86LtaIUNGY+gvli6w8C9m3qIV6vjBy8pFVt875ClKdLsBXa9XHHZZRLYda
QRjPo4J/ybPtVYXGgqSsaKDCzbxB2bsLsuRFJJHPidr41UovYXZ8YRyvBShOPUnGrL5QLnjZhi0b
ugBwJGRyoTLj6WdDid5VEvfGFDsN17nGVSQDmlWauCzWmlOPTjHpfRZgGFOUuHsUUaAjYeZNSrAd
VbEiLhRl82yGpxqX8xmm3K5Dj0UUVil1VlHok8KiAn7ctZrk71KchoiLqHrz3/NtxHWc/ja+fstS
ceeEdV83AxawMhySgRwgwQSHO7Orm+/YC5nwzK4B/xn3gQv8+A3jDLaKtYY/JSgVu6+es5zPkWgU
mgQdMqvRvLFjJ32M7nj55sTjJVNhS0HLPlSPkGMbaCR1aw4iILmEy884nnlWRiDiyQKqypJ38bDF
RolVwXmOwVEJfhrronaT12iB/jMLpfORr1KzJ1jAv5iO/RzG7irY/GdeyxlQZtJYIiAMRluijRUd
31Nd+TxWRdYV0CReGzFGyyKhWvnX3dnYLdIwt+iJrUUumSb+6L/XBsWa+8nwdCkunhQLArkw+Xg9
1QfVLqouOVR4SsMiWdp5qEk1fhUhq+TKeAylrzaPCCo7M3jjfHYA+8UspdnUqrD4kBJwXSQnSe7W
FvsihlN6tG9VFVE5zUkmamvQOndbj7R6RmHk7Uu9QEVKKskIySvkEhisPA1brsYOR+XgwXntBpNU
oe+Nw7iepG/lmLNut/065hYn4OcDt34AViu6979UEN2j06kxCHaQ7G/cMSPS0ngw4eWOTAwYB+q3
eBWcW8ZCSuI6DhatLMzMr7kNi2YWjes44nERmO1hTMfTeEPFIt2abZ7O8Zjt0mX8Qh1Ih/ixMfdO
T/kxukZ5SjO1Jdi0wRN9KujSI/JmRo8cj9WFiXCqDGzCtQEsmoBtWcmu8/l8608oZH5UqWAH1ovt
pCBPa7h8lbsjenRuB/iusw8tTZbn6tb0OHunRJJfLQoh6SMOHmBRlyQ1B+7nMDfzIWX4h0tSaXkI
S7/C000depN2WheeIU84XQhHVTZJtuSl1m2YGAGqLrHZEqlP8SB8Zeo1DpXZuO9Z5RDxE0ma3+Kc
7mUd3OJmDaYnx+kK07/ZeTRjkhio+fgIdNgXzYIA/hgZZDdjaqC5HsBJpT9rBYzjnQyWaKxbSH6i
s1ZYpV6J+fI+LvvM3oJevlOU13aS4QSsdeZZ4nPLJNHK7koJ2ksMYzJm1lMR9JoYWdLIMxLyhTNl
5XzqKV89OhuPeNIAPjrd8BZPWMk615TnKWrInHGrqf+rTJwgFzymbqZynK6Etm07Ci9JCFbV1Ho+
XNtrtBUpPjJHXgZEaGZce/pVVl2l9vCX4FKk4kgdYZXtZ9qgL09km9s0umgjETkOo6pLOQZjRnoB
AkDKug2L8T4Qb7XbeFUHrQg7ONHmkUdUXVi5EH0HYLC31Cv2oeR5v36GnjlGTm5Tds4gN4DMNOGq
wRzEtbtvq3hq31/n7PgRzJ/dJqhe+AMLdWU/h7PzJ7IgYNe340S0t1hZn851Ny8FiEyctYfDJ/0f
Jn7TNeB71qN922FUhtIevVPVWA8WnrGFneItkAjaLQH36Eaj2M9TnLYurBAyl6OVsc7Hjvaaq/rg
s8BkGplT3x2NGfVr2NJlDd5FfylesRofdGVNtEz72FKJY8RVkk3C1GPqKieqjE8wboDpaHDrMxVs
SW4Rpi3UH2txkrROZV0hU/5XVnXR9v/VnoWzqSpof2TuRV4SLmiuXbxrmXMfzuLh5QT8BnqLLzVy
wLFUnTYLgCVUzVr9m0yCfASu59UAnImSbmxzaQ0j5Wka8dZBV02/pdpMohz8/KAKHe2y4G1NOcN0
bXRZ1mNf75eQagJ3QGlYZSr/8r1+vA84AJIVupp7kSJ78c/rwrxCjAbhF5kJyjVrGPQ/56+WMCd5
FKcpO0SsuR/J/Nml6dT56afijj8JQpLhCSKOdKQxr+GypOdXm7YAGYi4AR1HvWt3hhV0R0dKxeHI
gfgH94TDXzq6+GI3CMebVNw6ubpvhOcufrtFN4Opo54gpdSINOAL76d+bZNhCkSthoDrQ0LaWkkm
dY+4eekZ4PCq3nVLhN67bPftTI/MlaErmKzFAoaY6OoENCQ2sydYXbbj6r7wqdWXqjWZHfY+8szY
/NVB288HWNa9aHQ3sepxPM4z4fhiTM2w3KIyMwfyZY1a1KWMkDNNpCATwT7Ed3aeaCGofs4gQeP2
ZmB+fXjCp0ly3VM9FapVCR54c2Tv+AK4svCrA0LqOD4+3BVjRLOTeAmvzeK7NhHnhTvc+u3AheMa
ZOx2OX/Lfkskn2X6bgInSk24k5bbMxAKT7P3VJld+2RtRgXeFdX4rIfaE6StRONo8WXTdIqrGysW
pqUUhTNaCK67NPBl9k2mrumW42zWWsdJ6D7UxVGc4Q8AGrB+ozSoEUPxnO1aV8P6rt73+F8bY//o
cSnIdsLWXydnI9sLHbIUDG4FfRRMb/x4Q0ckbk03yoARbk599P35ruiI07ptbz1kwyPQ+u+YWN4l
dE2YkaZcIrZYBXsMkUn0agkhVDkZ9CT5LzOkAzRBzK3TX3P4vVxOgI9L+7pQho3VBWZWT+aJJORq
xi5eRgIb7pNK9plEVho7ZVFRioC1foVuDuH87uDUAsprHofuQkWuwOGuUEhMw/nK/5dikvdlXI2k
izxl7jA3U/pYyHoedyfCyFsqjiieTbJi3xBiL6NWNo6F5CX/4WoOiszFWoJR3T0Em0Ax+38mvf36
wGQlex6LPUgX1Np9pu947veCBbnHLj38OvOGMFS0NqgGXNrITS3p6URkXkHdSNT2IeDOpL6HKpJJ
nd359gL+DHuRI6fJ/0kSVgMA3Wnksv1JnNJ29MoAOrbhcrvAkg+2HTpj46HzD6R9+YKOMikvHgR9
WOV6TtjjnW0aPe+5ZZNIdbFJKh5OeLf4X0e6KzNRQjn/EoEbxJUfwV7s1fLjUDzUAaum8AP5Vtn9
vP7uN1mCIHnkLet9OY43T0If98/VZb5U9uWdwac20+xaLzXxMrpjVSWZnL6Qv6v5Pnk4r4OUhdC0
HakJtGsrtjEX86H+dBp8heVdX+hUcmRMt0K9WeZ38To6bTzMeSl+HYx3TQEi9XRard25yD2YqCsK
0N1snuBMUl5gNbTB/pl3fm1ERKkptIpEQyaNinaEujiMJPE/oyyhFtkbgm9zfuK8+ORnAsuOmSNj
b6wrHgalO4BLLbbo+1EAQBwXVhQwWAAPEo5iCwe51Ka0Hg5tzUXsCCoAWrURBvB40hyqFnQcUr/h
TTu+xX4vJNaMiW89/r6QhPKQUbcFQ5S7W+/GE78Z5QvxqGbNyjn605Wntz9rFUA9L8KVU7Rquy18
RQa5mItirKbehwLPy/T2S9sKS0tbzaKYneAezOJx6o3iu6VI9BguVGlUVMUFf88HdnRN1IwZK6gz
zyA4f11X3QXU64F6DYxGE70E5e6airEqsKpj3YB/3iweAiSWKvi4yZVXuuJL5th60wbPDxUmDwkr
I7r+NotgcwxAjZUctvkrsYZHy2fa0twh+i8VeWujF1fpJLvzGfhMc0c/Gbo846lL+Z4SqN3RFfvn
BmMFC9UE9wrIJKTVFfKsQoRLhKpzptyKDPBnfUBPYcJvCmK/RYMbccF81NFc9YkpZEN9XrbqugW4
OfWcaSWreiphqYs1157KZQPBIfVoZlC6GnxiLm42+/LBPIGQjheI+qinGIlWxSfHeR6jTmOtJJ/c
G0uhzjjsCN+3zI5rJZ33wM0FZCbcyYj4MFuiQom9twFl1WbPKXMKtJLNPyuEg8oHlEI5YBwd7eIF
3dhOL5a2UVIDSMw10t7mUO+QNKxNzblOIU0mDc3a8z7jIOEUtnM6bKUUR2sJZX+JCjkN44AN+dgi
puSXZAx6FV5uwf3fn30JOw9F+8hETiOOVB6J07tBpUAE3hhoPzq+1YzAdCVB7c5txo4YJTmdw8xY
ErwHgWEDlw4fp3u8npcBtE5kG9ORKWvBrFtxNsJ9vpDBj+7S3AAqW/Uy3sPyLUWa5crp1w9jIliT
Z4zOHJRgxa9yhIHX8prJGylqEhLpB2k/HSAoL7H/J8MMarXqvWBXGapsszdmhtf28hR4yoNtGX3b
GSPeaVST0HG2o4JMwRVFsCL6kJI72UIJkiPHAtgu9zhmbVKxFLsOAVwJdSwYyg43ZzCylEGz8FyW
/sFkMr/NNydbTvHSE1gATDzrUXO3EEvyUyrEwJARm1Auzpu40MoMai0cvvKFeQ+QlKOVig5ibbsw
BxBqfsuINUl2e1ijSeCXDYlxfS69rOW0NnVDXzR4t17MYTTPoUYGx1n3NZxRHweJCRVlkeITM5hd
ec5kz1b+hjnqm4LNGOHGDuOdZo/kQi0L++ii25y5u9pewlzoaFyWU4IXQam5nSqi2JCgI1zW6aI1
+6G9jNG04S8qWnavVEHeInvOpPboX+JbdSRexuxQoeJo7QwxSQHWfD80hhHjGvmMwQmOrqfYuhKM
83VBhca125n7ecmpn/famohMEpxmVtUfC7L8jJvjXwlkUCYQA/lsjiKvDIjN4FXd61zhL4lXZyLU
ImIZsVniKYoMmc8a1w0lwhtEntQchwKYE5QvdX78a3lVschNc9onBU6QPP5IrJMU1ftIN0pufABI
z84XvzJpJQif9CaHUOpVBee0kR7Au8ZeoOWW/SlIVlwhc46VLNYH6gfhHJsh4hRNRX+toJie7oOt
+3vlbX5voIrcgqTGx1nTvJPkt89OZSVTazpPb/u5SS3AI645dYjMyqPrw3RvA1qUU/IFyIuAloIq
y0v42hOpxggwPkW5Eq9oxbjNtu2OhzecEbcC05Sv4zG/cuMc8mAzWMrfb6LRimI8LMgdTqMa9kZJ
AzFPFY9IwcjtnELhuZaGgkwsFtfKxrnn/NebmJZ1DwNWDlZG4mM9KEi+LyYqaPoxmjcL2cMpB9oi
zRheSCpazIeBQ63BNpz6qq+6Tyof7CW9Dp6pfX6rV/+zeSZu21ejzmyAwIX7++pIxwv9xNKajonX
2gLXv8LxVgh4jpuZAI+ClO6pJ8AneQ8ybU+5CmlgNGx6dgGxpf3rgmsn97s+s+dK33vMcwH2LLoi
7YMx34JDC/+JBXCCLwk17U8XMmf8chlbaV7yrX5N9fMLYZ6Yd+JcFqX81EjL1f+Jm5cwfIy2VmTJ
M2VzuFyfX3eeFPrZiOsvdJcIw5tiBFZLFPoZoDaoCRMDsUN78Y9ZkxkrzAo73SJt1jJpypIgByER
4NL8EG2MPQIW/GY/aivYeGSpdWj2C4sJR2DJ9iW8pebEIzLdqIiMiRThKfVs/TEGHnJsIK9GH9Ev
4lYZyJ/1PPArLlGQL6omaruwrNX4C6MW5Xttg16v/13AkgeCfVdjuNOhkaiSZ7402E24fIf/vry7
U/VUVHEy096aeFEzHZL3hBf5Wvx0y2CuOcKsaWjcetH7fKSBBED/D9z6sgzMKEOhDZS659OCZW+H
cNSeL7PC0Ala28s72nBdJUe3HdpF1ZTEkHAbRVtlTUyMTrtHcvIW9IkN81lDe6OIM6I/mB02R+Kc
iBGagDgarf4hbrrOfXv2Xyj+4fyrQn1OngK9+HU+Ay3UmqIRMuucovp60KVzXNbLhaPKynWaRyM/
YnWH9oKNa7XM+BYQjSnRU2Dm0DeQGZHrltnCuCbz+72TVYTLhUT7cdL98rTDtNbeMbwb0vkFDzl+
bkb+0mrXRTFrojaxDDu0ISZLQP+IjiLl0hncOpKaahckOIt0LZJLkoKBpk5tXeDYumyJq3IEUnrZ
RWOXMV7p8p6huxdOcs3bhd0wssagxA455GiSa+Y2ARzQ7wfed0c05rK7yAg/eMgnKNTy8PPJlGP+
1PUWpZTclbkm77YMFLzaXgrRvXwb1CXDkh71PMc9D4JJoeVp3aaHBRDRjK8LhRAbJKU1PWKw08dJ
fenDdsQp2atC5g5vHodGUupFK/3jnu2w+a9Fnh872H6rQxX7wavHt3R6BirVocG4Nq9khekYLI6h
g5U5tkKUMnVpLPJiyLlGf26hOuc5kpKSU+DEMnD9IPfoGcOgFgxuOL5N6VZvBMepytuOKeOddENq
I0ivlXekSFgI4OmMTiWwg+k4U2FeWtAPZZdJXiiCXJbDDzqJ/94TrRAAb6fbTwvFkmn6aw6BpU4n
u95yI2SYSYFAiRbCxSaMe/NFiQti+xqNDhZsFwLB13BgYIWpmDEJDDTb8i6We1TfwIjJY1+TEl9r
ac9PK06OtqI6WTigyctlGOtNDBHJDQHgLuZ8oosZUrby+/i9mQoU2JehInUL8BAOgQ2WGlskamIh
8aArbD0j9R2kDvvBcVJxT6XJHD7f7LFpbEcbpDS8xNogFpPUXA2szw1MibuTV9AzYjcMAQJF4inB
1sODqirwHJReCjSgIErgvSBt5291YbtVZnqvpx6Wgw9+z/DUbgCezzNcXUysd+wQkxK4kGuQtyVr
iV+j83eEt0R+XOk18zp2kahq4lU1yYaiQ+BegrrDPQIgSOTzmQ1HIs9gjPEGrIxn/JEPuO4tMagy
7rig03vsOE+JPvaj2niXFepAGYUceJTR9964rkVD5u8wBgKJFmcO2Hg6lJeFsEIGWHdVkaX5gTc3
SLKFA84yGjyO/I4Pj2lgmDGhiQVlpWO4SaSkeX7XwHJJVrTxghcXsEKkDRvNn76dHuZMJa0HIJTL
h7ZUJoCFMRHS2Ndb1hkIryuVfw7kw8Z+MQHrppUhT+/OIEyfMEHE3WnKrEtL/f5HoALuYqwkWDq/
vfXmj0p4VJ/iUeIUgLAcUTmeUFgiF/kAB7RRm2V8SFi3G1uqSPtSuvcSowRNxm33paJ1zFscdRth
Khn6vidjvyOvTHwb6Aj3wI5ZkdMyIZF8fe+tpCv49k/ZL2K586d7ehWrC8fm71Nkgl1xQPAGDuAY
OvIEwjAiyxv3xzgBwLe9x2S8cNgalH+CNdm4in9xapf4vT7k+BEW8J+8I+tVKTwYYtsH6bJ9+dp5
sWiQvxBQHu98b/yf16BaGUvff0WtpMX2izqwkj8SDygnNEhPUdTuyQJ792QygPfRjjmyw+mHzwIE
Jc0R3NgUXZEfVVY5lQicc86eJXZN41GIoNSLOxXMi45DBhBMop5M4rawkUbeoWq1+2unmj6TN2XC
lBgQa0l7jEWLCP2M0ilfCn5DJufaSWFGlLOZCOLXxHI8PgIeI/E+4xqBTrAWE48GV1aMpnTdVyXl
1Njj39Kxyj/WwQ9Lszn8tJa5Ptp53564rFLRj6E4pX1H18u/X67na+cS155rbTaI7RJzsIZZgGmK
LmieO1KMivmPgYzXdU9T87JH2kDfPmyiNlTojaC/WG0LK0ztKkErlNFVp0itUAEucoFjWx73JarR
DChszdDmzmdbJU+F5wj1ra0RAG9nMItsyLKZWCwyOrgrDNZHdsrKHvRWvyL5loARDicl33SP3z2F
L8CIiyajBEzjIGPgcGvvkCWV7WA3uTy0YGn4bnBGYVosnklS47iEU4sZoqlZ9Jf2vQjM4r3v108u
7rGLgUxO6+c/zISQlf91yBk9EGW1k/8yHgFEza/zJOQdgNzQIVhNfWk6yBSUy6KBUb+wwv26ba1w
YczT7vjCrCSlRJ/v+q2/bsmnZxfHR0t/KQf5gAcO9Fpyy9/HdobLOm83vUWRh86MBUgFSbh4BzFy
75WPXGdvd2uim9/+pBuMIxm+s/JrHI+mCpGbAS4v/43PgSNaCk9WTag3NxkzseYD+ow5tp09Q0VQ
qJ1X6IanxlKknkG+xI47EoclzdB6mbQTNgOunxQm+gRYpBORiMXU2hDn/q1jw0vicN10opT9tFVJ
AHoGstewGHIUwQVZZc78HGbVDNwcxMeMx0fW0RgfGfDWr9G2WpSESqjez9mu8jgJA5rxl3nE1+uf
qSSdgpLUBrGJIi04ACg6dcX8KarQkQObQq9IKg41E9TMEZo4tWZyb78Zzsf0ryMF2Lj3wg5AWnyB
3kIEVhGnTrDtVmy7EBQk7w1udOEhzrYlJuKhNz7a+jfcFcMk+0E5MqNrVzeLvJZ2XH/p7V7Uo4LU
h6YctqCYDGVI0tv5p+/9lXu1oUYeBBaSOqhP5dObzU4z5P/+Jmx3Mb64dG3nUGKk45m96cnTDElo
D2eW4G6VjK5v2n4wSP9EH5H5GItB/IHeliDX9WLZA7y/r9+9DuIAX48ehh+8GWnnpSuSmA6xeS9Z
lMFDa5goVWZchwNK4WZWi2UPM+8wiqq3aoad0UQF3F6pgczqGSmmNCEcr5SpN6pVt8yO7MO6C6pC
6zyiAEPo9hJAqd1wUx0NVK7Jvypk1HjG9nLwQyFWbAhz5COXCMMVqZcRP4GDqHzdsCDlUhZ1m4He
QhmdO/xoNCyCctPDZ8RbGGwDek2byvwkbVEYLBCQn7TSILtP/Pm5e3jL5flM7aKmAJoz81zpdg3D
nwf+n0bwttgbUul+HpEeNNOGFjqzFh+8TMsHHjZ7WCwsDzk/8P4zGDfasiwAwtohGrWuyZIPVFNP
jKin22x9oUeSoV8hrBR1vlta93JImNEdUkQ2qWSpV7eBC5i7ZJHWP95z9jeUK2VtY1mgNwImZtdZ
lbw71Rk6+c76WDF7rgn27qaiFO1PKV8FQIFX+Ut8LSjntu8clmrhvBj+Bw/d8Xi3xJWNThFxIFl8
PMJVEIZoQUW1LH9r5lAB1UV2z/JYp9s4HACqpuQojzIcc7LDbk81oKVu2eeEmHH4aBI+1ohZWgy7
UgmixuxX9GuZ9Ge9nbyiun6ssUcWjZ+AuECgn16i+W4guxcRMUcNEVjKXSH8gMb1b++q1sGvN3Of
aBLq6LBkSjrod4NPGuP3q4WlSDvkHsQIYKYhyO2vX2YToCLqIHWSSq3kqD4BI01vexexEuTX1Hdh
9tOJ3CfSFO0g1wRWIf0qOzT+23X152AFlh8kwx5YHfCTRRkdr3FUYhx+EOZ5eQcvUYtA4/G9/gZU
3grZmhoKO2n+W9JEOdLfRHWzb0qO7vqAaJf3rkj6yIpcPcylk6ryorSYxwimf1N//AGQOFcanFTy
bDj3dXjYJao+qjB92dGZDLJY6eqCOQluk0NR0IZLZLsi+5C5AFqjaXtozPwZynHfRUrAiq2XNunv
jWwzUJetI89w2FKY5DxvCYCaIXhki//njNI4RppVdOGdeVFr+5RWa0Qk5wQ+7s4pZnLUkhTveA6e
V2LRXdK3cdnnmsXsx7Xgda8kRl5WrcKmS7dQFIh7PRNRrINhqZJteZzFGZx4hXYKGMdLokLdjtpH
7zejSPZvUjMi/Al5Me+Qs1M92AgC1ie/BvySDIJC/9ZdXwnaD1Ts7NGZvp5Sjq02T7lTiYLopQfn
iqfJPVGVteGpH3NFSmRHBzv9lrQSVvl1Xzol+g0IryVFaeOvBgqUydKJUDeBMN0ZTah7ELPqo4It
IX4Ch4E8F+UhwPu3lhDt/MrI7VjpqJ4RcOQw1hKMjCCS09LMKaiLIRPfTujv1zIrCb3njaLKfRBp
aoBIzWCsvZ96rJ5qLAtnnv86tXhjaTPF8GXzzULSrA2Rr2AcSDBzQ3sv/uXNtTxS6YZF5WrlXoLU
k4c4m0ux0ZW+ikTTRxN4jhOanVs818uoB91FYBlPHi7oUy31BRyQw/ReGpQEqdcJ5mP3Az7Rz7wT
FmFCAw3d5PVTfCTbYzYzD/aKCsNJx8tfT1vQHAg6FM8Oo2OiylYHklY2SJ6jdXYjrRSaJAzNW8sL
Ut+CeFrqwKYYoVTdErhv28+oHDlt7OSsrRksvFx4hN7esFsU7YjU9W9tCK4p+Yo4lTGQUW+c4YTX
26iegcYgEUO0LUW78yElt/mTLB7JJJAMGtbCgmLCph51FwIGOye9JnPG42P3OQTvMeGhVnqHVuhx
nKsr/0MRhj34NUDdBwFcBLIaKsWGYm3H5EE4E2LL/0VGBwk3frN4M/YeJNq7rV8lc5omxhI81nEN
qnejuylpw9pmyY+7pKl+mXIH5iBEOaCJXL2utP1Is8sdXllUV3mjPI38P22A40cC7Yzvic7tj3zB
Ew3LduTk/Gns+sFdUTPkTdm9Bj3UhyYAjXNlp1GCC7+B2Pn+G4c+gM+O9B1pwCwjeO0zF+5qPZ0u
VLBwlkAWzJ+NZHOsgN2jg+zTR347OeC4hyI5/sTy5P/GiTe5UfssiD+jzAxmPMkZsNP5P5mozIxM
/nBnNx2GT2afWR12puOHL1xtwXqW03xstKJknPwh0wemIk5GQqLzyHb8cUbYZzAX4Dk34HhkjyaJ
XBrvn7AX8gWrD6u+B5eeD9hbi+GS3f7gaftKLJJXeK+lZ6c3uVE/2EjkeFEKZhV8KcokXblHVElE
NPVCQxlz1zkxXD42O0a2aThlZp6xSGCVWsguicFJscEjkSZuVtxBYU6QT4SoETfyE7bm2LcsKKp/
A2dKjPwCkYO543nP7fOYTFZwcjf0i1waR1En5en4qXHZuIQ9JFxERDHeUrB4zDtkFYguNC9zLCeF
kyfiUA/Yok97m0va0j5EMhr7Jyw7Quds3S05IwprHLp4nXACS8sx5x3k1Fy9EGFweLG3DfboT1KQ
TFIANbzhI67/xPveqCN1uYnfSTkST4ib4C9ni5eS0hRGtXIuQiPwYxA+W6n7WT/4xYCssdI/XYz0
yJe0wZcT8AGW/nUHMvtMoDop1GY4jg1eFiCz4yxdGdF8gHrsfqlBM718DbMPorOekYrWRe2l+d/p
Z1ytRDgfsFx4I8+/eLbP9w7rcZG1y31ejRlTMIqDX6qsvvfBncG1uL3HKn3+EBDqYMB6H+aFcvEh
ms3MXviMerKuXOnTNzS9EYPl1sCk2YUtSOes6ZUTWQx9Y02aoVJp7m3DRuLgWNgqpR9zjPBfZgQ9
dFf8/PV175t/EGUxaMnR8cyeOBxXqG/B1ZWUgmhk6i0JEScmft/sJ4R51GkWfUuXsw6S/L8eJQmt
gqNrd+imdpYsN6qtyup7SQi1LX510Ny4U35mTj0oasSfnPTPGEfmYkr72fSoL1E8lrIYJCF8yhb7
I3BDt0z46PLT9nSBMw/+u6HrlaG2fwCp2CSjfPZPeeDxvBUNyVFSAaJXUkd4CwBZgyMrTzf2giPC
1WoEBZwgphUz+17YKrggoqxBUQVD3QPSJIQaZ7WtZLRLL49jDsOY53OegesvRwCJ+gn7iILl9VRJ
ew8bIvfCkk/Irz2o+p50ki7mL7HPvWHy9A8hSdmvT7MPLl1ajGVyoK1mVSfJOAxByPoHvQbFNf+0
hZovVQb/rOY8jNfgOSS2ebbaJLHkq6hfBHkCRbuwbCCBsQ8TTnR60USP7RPo7xGgDfXiJLYyz4UW
337QhwSJkePYG5iepG2+23/MywBjMZ5WsOCYP/hthtpLdyNjhEL3EUkZJuQ0/Lus+26dh8LUg8zr
2VBebaaQ4PbBW47t1L/mmWMoqrhgoqveySk+78CaM8Fn0brI+T8CZve30OrC34CtD+WAzZsw3V8w
FQRPS6HTQtFlCbWsthAmt4ZhgqM5AFzO4H+O7XE1Tb4yXViE9GoM+QiKuDqiRyOIzOri0UbrXtQO
RcYbTpHGBg5FgwWyppKMNlyBeOlUwuI5pHXq9/h7GuLOTuIpKoGDjlunZSXjWKAcwdcbR1+/TzDS
1pJn4yFn4RP820/+EreUAMheDMcxan534p11Tgf6X/ki/x4x/wFrHxlcoiIt1WExq+CN/tdjvAlB
gRfmoNOLLzNQ0Fmq/LFYs+qnFGL7hOvOUHEsFGHS2WGbJGOBKHODTjP/ZhDd4LJ1JPaaIKZZEaH5
dNiwtmu7ZSeIPrr2czxMnNyXOLCMACD6+AiRfMbpPQzuYbCmWW4YvdGV3CCcUISJY4S/YKP2ozgJ
toWiZCAF46QiMIFd8KCekMK11AVWxGcfX0rPkXam6ja1sXJU2uN02xawEQGGFJK7Hrt7Z0Y5KkbP
OKJeccdDwLULT8eEbi3Dah46mRLeSrSSQKZ9Y/6se8Z3/Wg9G4NogrvatI+Ca8mCZffCODqGkgG/
bDFOvYBoeM+tT5ZcF8Zgl7WMJfd4tpun62mhQimIgK9UkY9YpCiJBU/NzaB2hPUcPQtf+B7vacb7
Bnq1E3OsmJBRLEHAkI7BiIR+AR2cOHjrzWVnn1Rs+HiD8bjQLpwtTZ1sbaot4ApPaYwicY5KIFbs
qEBtUUS0qcjIArMtKHDEXhRzqeKd9QJoGVz86R3x6E9Rs3w298VFW9wqVqyoIm6FxYP1qpFSBIEB
lS71EmKlyYfJJ2k+wMDwz8PZCrpm1jwYS6bFaZZJ0LxDYsARkidJvQ/bH5+GelNmYvwmmtuWTboe
ie0iObXSIAkubXP9jVTXCjVcfr6R2b4vOmm++SYxAqrTR3tNsGYZSOL+gApYiDnAjxqai+tWjpfQ
/1RFG6c4aJWUAJHE2js4eggepDerXZDjROUe7s2IUL4px0KrWxQMgbcddkiziZvmdT/6Rc89dL4U
PH8x7Jak5zxc11TRPjc8D57/H+lS6EcLXw69CGGzc3AlzIbJt/7nYkE/fIazYS8vC9mT9hdNQBjK
d6h3SfOzqmKCZCWmhi/sZ/cTe0+ePnkPoGafVmQRQtyTWHyjtg98egDo6Xr6eefdUU4Qq2lqqu8A
w/pTw/FkHHUdagS0KkTEXJZ5OIWy+Hfo4uAXLxPeJ79/rp5jpGW6kj1v5ocRjXG1SyezwtnnX865
LbjRNEOkE+RjUPx37pERL8IMDS7vZBPWJnMi4hgPFIuplB3o3LHT9tLvaQfvc2bpPq4VpIYCr4sW
rgLVpPM5uMV5J7iaEJTUjC9G8PpXllXElEdOVR2C402bVBIpIegjgsBqSv3VW3+u1EwzsAq5rYCI
eBgyoS2d+VQCIP9KblHJs0FWUBz0ReywzwoMr/8/vt7266iD9kwuTfPqH34J/uL3rhPy+M+zqakC
dxbvok1Poepps5cdGY/f/gTEuCgkq7jwDqvFtt3q1lqkV3/zJcvKEvDm04cGGF93AjWaCnVfMumf
uVYRme05n/+4pLVMy0efJl6XEyAXbZSbqAHNX5LFv+osaOeG7N7fWc31pa2aTH/wLasaYlt8b9+y
70Hge26N2Yxf6OPlIZ3nzeaYobLe42/wXp6Srj9SUPefRLthw/vZ7Et3vi584XeYWcebaxRHiVvC
KWYhENEMSVEvz6THQoitEdCeeLkQfJ6eemcnEGRTWlAKvkkLEnf/hWfgS5GiTbtPYLvfjMrtKuXX
BPjtXN/ywz0OlFAXVuS8/gMVj2UuDNJn8iWKvsmRFMaeCRNkcwgIIsLD7oyBDfvKRHjazPeZ57K6
91l1O6wJtYYFy3LbyR+JBTc4r2bhAFXlnOR633K4KQ2QXf1za3koGNJW/0VSGJuQGBTPjqSigQ8s
G1a7ku8QJ9kwKq3L4V5M3i9VqN5mqEyj/j7vTiECpoMoU8PEJ3CE28G2YMlYXccnASBGtTY8pOTl
n5qxFsJlnKrB0mfkl1AOQ2do3R7sOF4XFNklXXppQ5IjRVP1/SX1yo35uOqr8Y6A+lWKi4mqycoJ
DypcFEFoe3VoIQFBf1xquxvRj03WGlvJu76eDpWTL+Q0UmnNNjhfBiMja5k3ni+OclWBVj8HmRi2
MGPwwARLkbf1Cg7B1KmwHDnMsuvtFQakEC/PJ18+CoxHa4lt8dyUnmVbX1syu8YNCnBCI4Mr1h9t
nn32sBnWHOoE4MN/Bp4tQZZ4uK7GAooe9ZcQquYnmek7g9brO04bNC0YZCBcCgy30ih1M7Lgy4oE
uXoXanrNx055FGiqqomOZDNK2KGHu2m+cZOnZDmX0sbuG4IOewG0oWp2guAZ2BFAo3sPJSr765p1
W7jN3BAgyPSSxfc/jUh5dm75VLTF4MePmZwMOmO/LQ+zrd0DfEte8lED2iRghWO7btmiwoyafHUo
eKAB7aEwH5XiId4jh36i1eRl3FPvXci1/nGr7rZUeibfx4HxsNxgxBlULB+qmTghAAEeolMtYQbv
VkjCnBivJ2fbY3/7uvBQbyF0rYSO5FPbUAoG8WcvHDDn8azv+PI/MzVdCOOn+pDXd5bxiHSqDXUj
8YouIyP3Y5mGvIvCxwHE05UjrD7XtOfgYQrIxkUNi+qzIuF8R9SY9f0N9ktVxf5MTLHmkaMtttnQ
DlBnNJnXa9JYClm7wOAIGynNlCJU/x9qwXLMQhT59oYb2pyej8SIPeHqHdW49+T7ZxUosUiOt8H0
vrRqfvms8tpMVOSMexx0xBizGyqRqMc5jUFs4KNJ7tNAbtjXrRpbHKzVngHQaEGOniA/jD0w+yHF
NL+su+KJ9qag99I3n4s4rR3PnF+bUbaBhxhU7XXSLvBPgtpSkCmQY8luhixCBaXK6X88Uy7aHC/r
rEzWQ/SkgTxcCoZjN8Ugyuj1TSzW+wddX/BbA7WF9B1utE3hgLUjQgOy++6JuL6Fs+xkRC3XFFq+
CUv7Vh2GczkKrYgNTnejdrN+JvYY6q7A1XQPKatzKKM7VsuxKo69426r+SkDqSRaIK7n65NdtUGV
0SyP8crYHLsEx4997dFCA5y0MTEBYOO2zcgthUdOTUzOJQw0MtWkCnCu9v1rcsrFCwsEKKRIQqnk
R/k8mVebJY/wT5+xCeiWEtTzOupWNTWaXFCH5D7+YHp2uPw5OTnB6pH+JsAFe1ARmVOEOSt1RB2Q
B13bVfsnXuAuY3I6XK1TWhuYsOOudtSUW083QRlgt3N1CiL9vNE8Am14yNZ4KkxRHx+0YKe26B6v
lNozmnMShVG6kOU7Vr95eaJ4UxK+I4KxEvi3a8YMGRIV1dcVcBHBmE1jkq3ROkZdEK5JYZPtgvZZ
MYxAUrrJVPll3vVAkJ+8V+0oiWaDYPTY6wKPlPXnOdH1xWqL+GST9oyL+EaIA3IIpb4Z609LmSHW
cuB+n6GQvYu7gSN5/nyJP+u5pbtO+4XARQ/x2Xcv8tyeIwd6juvFxBpxQCJyG/K5IlSHqLlYmZEM
1KzcihtxKk/YK1fmOapr8/5lpNCi8Tsrz/U/PWgkoFtG7Nl4B3JFsvv4bx1r920X91sf8WymDCIb
9m0Wrdr3hnJI8xMgGLIQ0N+nTpjExK3JrOrQVlt826aUzAGLey3MzfObLNkcrpul+mug1oVXEdtL
7d8KChFEfC5ixxnHt4+0ksndKb8VEZTzLM+6WnLjKeeiLi1sNuQFIOMaJ7syVBs5Eh50oGXCHcvU
J4kWCnFbbqD1tV1z3nexVNlGO54E+RkrccrIXISASAmmMHksqsvY8ay3ybnHNa3YVSHH9CcJclQs
zqBtUwrxI3G7LcpqO1sBJX/ZnPO632Gq1tYvDVqjZp3MBtWGplRkG4hvF9E6SqK6d5VrfZytQaIH
Hn5daVyBjHA9ZbBa4P4IIvNllPG0Cje9Ueps14o9nw0rlGSWeW3bj2131YLjeHmcCUxJXZLF1K6U
DmU4wjFDXuIll+yqkJzAYWBPTWjvUKr0byFcoOvPCEMowItc31DtxZvQBk29xZMG27HHGpNdBJ7f
rf5PZhDrqxbZnpj0C6X+Jqm4JgP9+03v22HR27/2wYhoKAV3nbrd76NFu7M1lmxqfyEb5EcWuhFC
eymvdDb/SyU5w9Es/Ff74UzvIMniXqhZj4DVuTvNY5Hpw6TxlTMr9vnpByRB/n01qxai/aCCvA6E
xCal7vHSVO4he62O/PQDYByzq/IkY4rgcgOp5ERsrWEMNGbV2BLxkLCFrDbExGZHFgBFUkdfo1pX
1lSIwfe2v8dO/xwGSKiGa9bhPi8YQy3jXlweeEbjCryohAD7YGyL1kFcQEGNBaUgM8adGMkJIwdF
Ri3GVE9XtysfjMClWQhW76e861aGmyRFherp8D2OBcuLucf64+nYBPfV0nV5oHQcEj7gs2Qr7IBW
X1DcgdNT2d4hofeYRAu3pL+KmQdfQSNydu1+gO2WXU99AoPKsGPBsOWR0rhE/jA+mRnPYKQA7yaY
OdyyMI/+tmFhkIk7YuPY7mwQ9VB4iJgcXPE7u/hAQ7EppPe9PKTawX55L1GtMlfILpgy+YDWh/M9
6EclsVxbWOhUVZIlNDNRNhjhCp5itKu66RPpCAVPNwjITKk5is9w9/7G0QCsVawn0O5/Mp9hn63N
hvWLQxDXq8WBPTFuz05QWkZ2zpREuZ0fGYUvz4xk6sUDl1lWjsHWWgV124jeU10rczaeX6iOn84H
5xgzk2weI9RKTCeCqfKW5uu3KL/EGK9se0s1Rbg/y1FmdYa0Wg/MdTrPwBLDle9hbbHqf55IWA7+
NKq1GJfDWHsF5qzMpKVaqck2njvUn5KtE2MKGZt5p8q7tVJCLp4AVW5yHJPpnIekhGUdANJOc/6N
hRdNAdGzv2LAMqqr8gey1iKSoNs/vaU3kd0MyFsv2v+rG5GRdJIuBKo9ARunbD+hq3km/Rsow08r
kyVjoosxozp2n5pBmVEkACE/ekfqycqlsCXsjb3Iy/zVWRgvy+J3CPRL0V9bOPJo9ghL0kKeNsCO
OnpqnC0l3fCEo2Kmef77BIJvOftsBB8aicZzSeI7SZcqtCnZN6ZZYFZXLgbdYGYwO9mHEBoRhJaq
i215yGVr3z6QfihnsdJ21I+wsdZq89YAIFEHpMgM9Nro0vr5VJreD4dkcdS9vUEFlm0sTwwhddvU
EOVy0mOpIXbiOkmPIMDd2N5Hi5VBH4/g++H1Q/j58AyPNKYjbEMSmVYR9UtsCE4BsS8CcsbDjGLd
cqS4T817VVDfKbnO7kK1dM4pMk01zfh31or7aIdjYRxi2QOxMH7qfEYSOOuP3QSCtx4hAh8x3Als
XSDfDp4WALHUYgpDxRwh2LF5yiPWKhn/fwXrn2F6tyAlFe/BgXEh0qhc6iqKyviRGEw3RTiqA/uC
9SUWiAaRb2aBsK/zOyXeKy0chbwXluPEOfmJGhXc/jQR74ESmK9P738GopCigvpgjd/v1QaVsmLK
n+AgvV31Bhs2pO0fCfUzclk2TZuIJUC9CFCLdGFfctPZmreEwJ9cXIU4V28M8eJBEc38kqcCts65
AIukJIZ+bFbb0FglYDfsaOLfZ2E5g9VC8bQJ2hmgEMr99QOrK3reHlET6Xm5EFCremmOP+oUjWdH
dAe9mIWidM1HYBRMfd0FHoju55mpW8NzxvR0Be8OhOmNbf55p5Nsig3rY4dJ2pdLwkIPki+vSQLr
CvTaWZL03acVQi4/u3Qt799/l4sFIUGb90bFHk3QTRMZIiCPAXJlNCQ4HAwgz2//Qw9RMpu63evH
s5Y86HB7EdVPPgFUnoz1YsWf2KNXZuhg3uThX6iT3MLxx07go18wG6zzd+Pcjs21CO17+ToRTLb/
QSlJKfAG7jLY39WIKrdG5aA0Ue0VBFflysHFU5gVFuWL5iB8slcKoA8zxco8Y+KMT5odZ2FYm0IB
wfdx0cMCemU+UlwbbUF6kxKh89aYqqqkqngRTq5h42oqeAIYdJi/gytzUX4psjGBv280cZIE6fHu
1Far2xjNeEWDwV/HWhQiU8t1zIb/GvJJXD4XQiSNYcP1FymwLhdHmrn5DmseCK7VdDwyGdud7kxp
78oCUws6KXIu4hE9jZIvnGYcEEwrflRzGHWoe+om4meHHvywyoZE2wKLRx7F+TEhA1x3W3wXjykm
xXhyUCi/wPtPk3yD/39PuTQPzcZqPN9sgpQ3o5O8zn2J5RRADfTBFC0QKWxopZq6DgX+4aCB+kzo
Dv+2a5nrCkAsWgfPkDY9GAz32X+L7szcWN2eNz1F+Hi23qECiPhgKcRKu/BoQr1r004QTmMo4xNj
MwKQcbuFiJRLRkjiJoRTI4XXre3uX4MDyMg+Y4na2QXbFrv6XfQdhaRSipCGyKcizOzFYeMcbasj
WOaDpFyPeU40QezpnixgP6yucXIj/Azko310Qw019h3dRu00pX5yfJn560R4lc3GBSZOTNpkh4Ur
wd5xQG2vb+HCkKGrvF6HpQ6NcTIC+zmfXrIHE3MfCFHAGJW+EXmd96+v4Ih87U6SQZMeTvBVKERq
24hE28Lg3Emfk4RDUu8GNHlNzExRra3GixA+4USOoncQgmeCI6BLvYSyiH5IRuatSv7I7bxUpYXL
KbNddk2f6w7i9DuvK0nOwBDnbrcNx50yRHAgAnU6b5OqmkpugTmchbBKp0LBzXGvzcHP7vrK0lRT
mKUySDqpPL9+GywMxDL97R58vN/p4B5vfW/AKEzsk3zzQuyzVg3Dd3u0mn6fX/XjuN1pN6YuGkeh
ACzyNb/2Y2/7RcLd60NjNHK4hnCYe1FYk4w/v4Uw7kpBswErLo+kvdb5ckz7utq8BmLJN++OLqUh
SHWiiNYdLj+Mnm3lid1ECk0iazpM9qVZIqEjILla8KUkOBA5F0v3tBWA+cZdSIrUUwj6qlSSsILW
DcNT+WWAPCkc1/tsw7Sg5P8YQrGdUnG2B/+ifKJvONNLjwtP/Vw6rN53N7shq1UUIc+hiW8oQccJ
BugM0rykg8eg+DV5ZGPYfvInDGhZ9sDPhkAKGVZD0xR/IlHPedgsGJfu9iHmXKh9nCfINU8o/Lhb
K7J7Z13T+Dm54mnCYXB+BgG+5xv+QzOYSc+WUdI9S6XKFc7rkR6XbWre1wszUgrsC/tidPzwl0cU
wYogldJM03PpUi6GzVmYyLro4acvKjmBG8WdfztFJuM4LaJGnhAltzDp28d5uO6J/SMMyoH2N62R
9U1PUKjC318QaluRgbZ2MnN5WbvUuMnmacl9FylUOL8gQ5/2UHTt8DIzoPWCa4PefefKQT22aQHK
4W3xZD+X0OveUyjic/xIi6hADSiKeoqjim5lF8CiTWw7eZY2Jm/dcU4cmfSnUinOo+vAfkvMnXTU
2BckJVf3O8ZmZafJD64Vh+1XLJ2X7gJoVXQ+Y6APslMsyB/FjSyVAyhC4gH64uaUb1wpvGhW+orP
o8vfTHpEytIvvzgXKT1R4LU0noL1XqZosywtcK7Bw5MUT1byTufFhbxb+AWeawMWQxnYPMV69/CE
ADze5VeSQtxZuqNIRDSku2H/HIwiVbLVMD6a8FjmdoUSa9nPq1sFTNm3YCrwTIj9Aaeekuoghm21
MHYBeoTIXjvzMG8zSmS4IO5DKM/CpW1tVkMlnI0k0sHltE53fDvJ0gytUATVHPL9wzzrWnPF5jGq
L/AVANFqnmZstSApHrwXgZFbaerEHfAjryJVxN1tQSYbHfJuEDT9ndO860L+rBaKhuEqJ4PMY8AG
1AjujnDWwQnLp9gq+eiTtFW7BLA+OEbRS5YxQkr8o7qppXvrzlmGZWcFian/bk/6DKQQxXyVhgAv
U2A7DSCEigOq7h1Wyfutbb/QmuXGu71jFH1bo9lFMxzRJ5RvI1M1SyQXK20UoB1XrYEef2tqM+AU
DEydZMhe7VSjAMEiAKnrcKIXkHa1D2JkA7Ixp/0PKIpkBmk2F9it3VFKtF8Zy8Vl82A4dHp55dj3
B2MPNszRIRxTy+lKPy/WK2gUSVANvarXJtX6qi6s6KLUt2rPFuK59JSx4unNDGHuaP7MuvNRWVHs
vWRJmD3QTzAM1N+oL9Tjyuc7m/1hpeisEGuikkVh5eRgK7rmzKrkmNLy8VOwhzSFOkJi3v3krGFA
k5vj5d+5jVU2WugsEIja9gWh1NPVvPjj3hQoct6ogarpCTKNSkuZNen99n8Tzg4a3oovLePraozW
MEEqLa2KGij5DTeaqBktm6Ltlip3JJ0DfNs5FvRMIGbk50NAqYAaCArjlPs41dCjFSy27QPzPhYb
lF4Qjv5odeDwllbBI0EkZ5bnx9201PWzeCpqB8jQTbdNR5j5+vMr/nKOgrAMhJkUxbf5fvMqQoOF
yAJHY9jw/d9DA7wz0nBZJGI2KcltfEzdgXxEyy4etmhn4lZG/cLxKPbEEV5S5mpNu3pkXwAQz/qz
hjkoJOg2KPlj9qZSaOuHUFIZy0RrVmAlrq6w4xRQaIyvBeW/VfmirKq2gVw/uYEKQWLRAHWRsj7O
2MoNjWcsRcEeeFbjy8A0Bte0+39hokmPwnTFFKNrkCLjwctQ+v2jH9GnBXgbEI5rywd5Q/a1gC5b
BSrJwdaT6PFW6uWq4q1veDsJm9Jb+JfCbCJzGz2LvoNLoTz+bus+uDc9FcNEx3MR7UTLNARhm0+c
wa5UsjoXdKnEJlo+wriyd+bmXDIlaCS+WdSIi8oJfPqj9+EnkHGvbSu4+ehizLC+C37zaisibLl5
Dp9s/TZ2fVtgf0IkNTnprE7aT8xYGSHTHDHvLNhUWrYPs9qmIdn3edjfDu7koOr7KpFc0L9/7PfW
yKxIrmZiX0Gq1opbMJzYrQmPbKvOS5qqaCRmdrWOHrFPY6wbWib7kzJONyvQsqijE9hJnNcg0Mpj
zsgJMKkSN/rZKUOCz3im5f7nRWpq8xwHN/LQraJT3E9aincx4mlOl/chdPd2MQhYw/W6A+mKo+5v
ib1n5+9Tpcy+NesHI6Jv3kD/xNoxXIko5oF+NXPNaMwAtB+UzrvWaPf69NxmH9Hecs5aPJrOSMzB
zQ36807WnfTQb2I+HaKrO4fi+jjYxewtc9mrdI7JHdLU3X10NJP6Hp5Ccii9Jbl/wfn+w07YTYxQ
dVaDrO1+UxN5J2DFToB9zgWs9JPZPXcS95TfUMU0A6Wx/VjHs0pmUUbUgU+8FfFUQt/sv0KeA1a/
8uv2KZu5x3ww/70jWkVfSSzmV/1lXVs+AszWPoU2QTOeJG6CnPVu8nQDJIiD5WpnpwB5BggD9D97
wvsyYOsbVeKigkgpVq5pDU/3VDG/APrXSFkzIkFwh3wYPCkRneAwf9dQmA7CRXuPw8iCdFhRu2vl
GBPTmmyiGodwHDg/lWPFDyDJnZzI69Bnz4wm+CLLXWLsfc9PQc0q2YIkevTtxAQN547vv8typPPt
eQXS8lc5BShzCnhXY4uL9MdKOj19BhyldiupDVHQIn5mCjGAsbYl8ry0XXI+DCSLE9Gb/Hb0HXDU
7e8QTJHLgoQJk0Eho3cOmQb4a9z/JDn1Q3aLezUqwg4Z7irpt9M2WK0aHkGhGt9iAb2A97JL28O9
cK4e2JNurnJ+tnmeHHZJ3MyoFkuT6+aM4HdfbFBPvzmFTlcWg6YmYzYXvmwI2n0PB+vc3/5h1kPA
n+TvXq/MFce4KNRU07b3vyl1s+gksiw4hCQrkHxJmlQKDRCEpMZbGsLvuB47ntga40WW34/rKBYM
K4RFcKOGsjxFDTE+YgD10Rz+ugnls9O4ziii6FojOCWufSkDK9F8n95ZMWm9RrKwnOk9c7NjS4s4
fdRqwACQGdzw7OPdCGc75YojUkjyst2ispXTDlAuSgcmS5ZgcKQ91+vJMV83Z7OaMRHME+c2vsIq
rgq4uPdh/iZVycA5uY1ty3JhosuYyTs/YKpwysGEcEruRLs53+2df96T4+wUwtmryAxDn5UT1NQ5
fz6YdHVfFfJB3T4C4fNuZx20AB2piRWnli7rioyIg/Ww3yiyG3keayOnvFaDLJjHsL8MAJFE4U9b
W7ctcgxPA+VH4HJBy3oLk9SLfzixPFK06cv2BzjQUCJohQV5lYTyJVuYZBpiLmDLSzOBDDs7AWcS
2WVWU4tTq+KLelyhGXtfz9RG33CkvHA3JGH26Ls1fHnThXbi7W5AO9TUjN6iMElv1rA8Vc17zX/l
s/vchmf7/W0NnP4uHaTnL37klO86jpmYSNDHayaHOl/vDZb0J7sC/rDIeV534S1Y3LzOZzy7SLNL
dc3ypKY6t1/NoI/LtZvcd4qq2aVNgc4XH4yenEvPt5zfYmje1cbXtfb9ztr8Rir+IQVKli+eLgWe
4BKrXsJcd5Qt+RI10Xmsqb59Jq8x0YOFarXd03jpHin9piVZ9is6lwqbytmCuojv496/wgaG01F1
YxxNsaRzfaiH+ZC4kktg0dB8DY3mGqFbojb0Svrpv5PmVYIurkR9sLCGONVBHSD8hdXng1UkmU6F
+rkESZZPBKfXscdL6DmbJKorRuK0iQsuMfGUF/nTxG4ZpFFKv8ysLqpzINvihXZhEqfYTYRGO7gq
2t/8aIPTA8dAv1CNKYuY5kQLj2ciKoaO/7p8Hfe6aYJAJ9C0VFA4w2vWnh8ojQzRbtpfmcntNVFR
gO0um7QonDwvd19cGtCdWBsPfU7HUhzSGrp7T+RvcdbtwldSHarepzX5lnhU2kBn7xuZ1M9hhRjM
8KrHoxOybWtmpHsNvL6murRuMWIryLr7exzF2MPxQHzI+t7yXkHodDR/CTaJ8KTEbpS9XUhaqzCh
KdgFc0lIfL7jmw7py4xkos/jFvZaMEJZydf3llXrOrvhT9jS2aQqKQAyJ+aJC3mlOFXRX0shoTc8
tPmLysuQBVNORfoNNEXeMrnv3vhDv/dNiK0feA4LMdOGnISTTEJ0DW1RtgK44tkePEDh+X/tnVia
QUaQv+E4arV7ti/jfqMTPg+yf3j6HCKupIMBTOBzFmwruD+SBUBz2Nt+jZ8V447Sw6etE3R1MOS4
Z5xV+nbKrhdpg/9mIN70QQvtYcuR1/Ub9zIcrIXvV+U7EvxxPUAB00He7pdGvhIdi6pXnXs0Qlis
EN3DkUj2ARSumeT+8GdVWJus+dTp759bTxpIK9dzHDm7iPuRJKSHWxUCbksVfF5BgHS7L7d8XKsF
YmfnS50BOQRq1FniIt4WAUl2u1DrkTNLUiS4kGZN1JRAo13bgF/Wlxg+2BNGT+8U9m+IYcVSWu2c
f1c9kFAJti3EOMcaCWcMAodCJBtcsUsSvXAH4KAzoeJUtG4B9s9gG7Ac6wLn0vl1D8m+jvQL6Iwf
1C8wvMwZ22yhB3V9iG0AI/hJ/EkqrX/JJZpNv9XCdCTB6cQV6ZgDj2sBBWzfL2arySp7wvBhQQGY
Ja+v3tP1RYM2Zdq9cwaVHIhWQlSvt67ynHIiJFpML1mZAzLPPun+NHSgNHFNcHlPPixoFBVPjpYb
afIGmQlYECB9nidhJdb7JkTcyv4ADy2fL4cLDvu+NWNUbPj0Tv4x2A6jIrBca2Othjvr/gq0AasB
gMWMPKOYRo1sjBEbJl+kHLLs3mJUc942ufUfgxVILzlUrdEvuHWBMV9/ao1VXCp5OCfUSE2KCBjK
Zde5LyXFxoLVbpJ+FAblV9xdbCsXwLLw5cfIpTdLIn0sPhQ+XAxO8+yR1zToHdr7lAi1B+KhsRnE
zRkV9paTaSPg6REyP4rWyXS8iuve/UfTpkmQolacGwThZTRQ+1PZm+KvAu1FkElJ2llkGk0TGPIK
zbfhg0ArkplD5+wIzHg+pnUKcswh7tEAgw7HtOC8zYLwrhYCHLDP/47VNKqlHJ/2+5ZjiOvB8IoA
hzpBudamKrR9iHjUBM8Nwkgm82UNZG5l+kSjB0VZw7PT92Bv/gB/gS0x2qjJg7DI+vGIpM7XBZ0Q
BSMxFSw0oDPB9O2F2JObExyE/qxvYKa4vMBr3s7gkEEOcCB5PiUqb+i0F7JsOi071XSjJ4oS6e/W
uXtxRvW5qgs6W7yn1y+9C6wlbaWUwlxVxnWjSUN3g9+oBlRkNliUm95mF+3fVnH69qdjZEqzrKIE
W5ypAvKPJ8R4DpbhgtvRe4Q6mBUp4ke2wC1UykvSiHzhrkRyUVZLt2tuuCYVj8fS3PThBtQ87Rvp
B+b3UV8TFeLi+HvU27FCLQ7fFCMPA18cYqKxjHWteMyBW5DV6ao+FJmpuYg/a5iXTwVHz7knQpSP
yiLfWfohSZCJRA95PAO/Tn7zWu2M8hpD1GAuZnmW8Q9e5V9GWVvGOmqIrLgE5i+T3koLt3x224KM
YG9/FU3Vq8q0N91V4PUBz0HoYAlhnz6rNyk6dqAmpHx8kbsoZA0o443jehG/sZ87EjeHZYrE6LGK
m0AmDvL6uyYaSXPEWqOv2yP3a883IqZR2SIqDmrmQCPR0H1QcZX89xpYZ86URgNXFLgqVKYp//or
fYd0KBDA92WBa6iAsPblKey46TRjvwIv02EmZu6Gwn2cUixPQP2fXML01PKKiy0+ImQAIdx7aBYy
ruEhItAp7WoOvbImOxa6HO+lQjjXRmGxsvPrkVQDUV9fPmzFBcXSVUX1/6NcDw+lghw2v08TwKuS
5WMBJvAsYrP1T4b+wD3rmUVIUDdp5IKbX0NUFuER+d3zww4vRUMvRKUDFSpwmgl0UXhsOcvu95pn
NMiCyy6pSsC+IdM0XTuHxd0oeXIh8Twgf0tVA/ohuJlXBZvqgGZAjx3WjrFU0tXnTxii2bXsQhmj
tfvkN6RuQtsq8uCaJUHrrx8RmIz3bI5oKypHmiR6lMo2CnhiBthuGIzcu6lUlCS79IfMpFu4e9NP
nDlO//Yw0QuX8eQgzjPBhk8yKI7lCEAjshcSrv0bl4mxX4msjxAR6u3owvV+q8nvO/O8RJqf1Eg8
+wxsxNqfFGaAaSiVIwW+W4/JOSYpwQ9p24QBB/Wz5Ms8kDk5MSKp9nAtL9KFg/xKxvXXZZZglFm6
mqC9zyIXHWeSjnrZudr9bKEtGBWFoHF3d6pJ4TuaeWXxKqDY6GW2xpTgm+gfL+cRaxQcPP9PdkGq
Oepvw/hCEEAwJxB/EExylIgevU8RAf9mhy161RgGLYHWj16fDaAE8GLwuTyNbpO4xNJ8pX03b4oB
C1HbjPQDXG3WO3nB5m78DKlSyjZJRRuNOcWiFHrvxly8oL/XWxXJxTe+2C0HU7SAEjIgrcoPNnVd
9HKH9NCClSX+ap4mPqNAGNDNAr2duJQD9lgG2Vo5H6sQDnxJKyIXt2i18ErQiUBkCZO0kWY+rqUk
tUwXYTMzpPzIFRTdMD/zkC/8S+Nq6++e+LJGNLt8xbKQw6kSaZB+Sn1JQSXKRcNB6+GBIpnhC75I
zLg5kJHzYzL+5NkFgOYBLAj60XvbbfAuEu8FbnLkSrGLTJvdMay6MZBo9vMAdHShaZoTp+dvB9Sl
bLaPYwvEW2tE1I6RnviCaBmg/w9/W/duRjHwa29puhM3l7vjjAeKHcWtImbIbJXrP3EwZY7M7eWO
9afYhLDW28WSS1Bk/wzn6rdJpKf5buqhxJIQJLOoiYTb3GkGYUdXKQnyB2fdfMhYcGtZBBBGH4d3
x+TI9torje3ynetOneWwxoBfa6Mcw6NkVrRdG8zyCkqyuhRbylmze/Mkt5iCnnX0MD3E+A1MteEy
IyBha2ifIycxejXx2JuBn2K7mZvkD7uUk34ZrNVUgPQZcqktekvOVnz53uUOiwHV3z4Huo7ri0yA
/oi9zoaPFSlUZr1QYeqf5IuZjmvQjihviyIIsZfWxka7KDWosYxdh95pq4zpp3Eu3CMC+c1n+eML
a4de6SlaNV6NMhU8MJ8v3lh+myA14+xco9u9Fn0cOOWrHrs/KFX6A0dz5w54qiCNPww2bMIqyR9G
sQJDCrOIuzywxk4IlanNnfPjO5fdsOO0LXttUkUim/d4j882kr13pK/XfAVQEZScHaUVeOn71t1j
3/4y4HeAusFWXh3hig5xA4QmEQ55oBDdCsz6YZo1QTLMXIihoapJqKwzMAplyhudjafdBhBDbalg
MhsgMIriQjW0Ekil2rsgGdsC0RajrFA8imNYoxn8/uO0g6LqSphFUVCSlFUEQf4n+Zqdz/7dKM2+
tXcEy6Rf8yuPO+7ay8e4ide41SXilqOetTw41/o1bEs4lmaXTMQ/KzsJ7hKInzio1VlOxtCYG7QB
li6alfJGWQRceA3s0xHspRfHhsv/Kl6kNhjuoTlKBsD0kMup4xEgI4SNjdMRUI/EgplHpmkafDgo
UWzdkRP1Uy9LhO1jBgPwFvq/wL3oPeBH7shUt/NR4NSEhAJ4MQBd1LR34gYSCwZ7JWX4uNvg81tE
z3wyLrzj3GWLjEejBKvL2IGAx5BwZwaKegOpvzGcHWgI+NICjANQMvZHD0NCYFmpCFwkYRRuk88t
c1Ed2agv5t5HSpEw7sLMGiiAHuQCphh0BNFdlXX1Fh9QtgQUjyJy2HYQAda2avGlpHM5T0SB9OT9
IKC5PGvMuchZhwsiB14kMcPWTsMnPALCa7Z+xX2gIAZk6Yp1naMEqNlzzmeBoFIvrXTqu9+L81lZ
bencW4Of47oZGbBCuak+ANFmwRczCVsfM/ahfOZLDT9NxTf3GOIDutRXFaGriPxYfrgLVmpeMrxG
7GUu2pmo22VD6uYmPii46hvHr5G9rK5nzIaYu4nItAL/cY2HOFnqqBvI4F/uieQaiFYOnBCK+O3q
37AhiSrJAkFqedo/GGWv0b/w6KDoaIF2jdkGtXozQ9nIou8obG2l/y4CfDB1BZB76FvldGbmP9iT
l01rPXTApaZRTRq5YsRytUgRgCmEDVXUUolSvj5ibGrepUtlXI4iqL4+GSJxEs4mrW6eqnFHrhO0
WKKLbEBsjwnpbFLki3hRhJ+eW+/qq8fXhkTGDeaNf/ziGs1qqU90ljcP5rDQz9XTFa0TR7vtS1bu
vdhccMLYM8WqOv1IZxgGVmCkcKqsp17+t1BNyozNGPvBmEKrPc0kCOcv77pgPgxJ74arfsSpIKKw
GonpvoJ2kEIRjY40AG5N8NG9JHRW6IqJFddteYXRky3fQDBNBjMChlMsOJgNi31X81dQWrxATGXY
09Fcnddw9Oj3UPY+LYAyeDVj8UqjqROKDfgC570ZHIgaqNRQZPe8eRnQHPpsDoKJg+O4Y5kGry08
ODbZ53J5oOQZBjVPlu+WijmZ0poD8fhu/3aNXhFj6eiPMCyUhz9udoO6wlqQT3IJCrmSAX6E1OtJ
q033Vp4rdhGiqsoHNQ8QnkkmtzAoYWMZRJbn+vJjEXukmvL3XJE+TaW6ibZpstBGjrUN9LR78bgq
paYpx6+VlCf2SjYP2akL6hoNun1L6lBH/co3j3JeVK2PKI1c7MgiPeTHzTDQrQfLGNaawL3gRe6U
RImRVwYYfU58wjaD+JldVVRVDGZHADTV4sEA/AH/siZq+ZHDBEBoJfuQqFVzI/el6v9UJO0zQsj7
qel2Xcn2U0weWV8WgY9siakDFnvIfo0wShb0atsjtrr5rMEne2WGco010UZpsWOyigF4zEhzHXjf
2PHdXweos3q/jEAKiR3hErhC6u5W7bZltSXfJMl/3iy8vvWP74fRgfWHHl4Xa7jXsfCYjFdyEnek
A9dUBQMD+DcVpbMpZ/3f1d4rxXJyZ0Hn/1xbceG4EZelzZ7fNbYUS2OLIX/nv/lGBihdQbRQIbeP
v6xecBRLhD7ntPK04vQIDTCg0KpNmw7WsjgWvSb8XE4l5ieCAzxzENtKyAPnLgebA8xZR8b4vhhy
zi3s2wGk3P18Qk0r5Ke0nBPo+BhuzlX3u//kAbubonxPgGE5D0p1AmH6qMDo6GYfcUG3g+au1sBk
plBv7fgB8LgmItI5syzxQuXqpIVYEemsgQpzVzqOjCfiWIiBn2HnI8kIJzE48VzMUx4VmqbP2qlT
7hXRx/vjb8aikWCzBFrDYrCTfQNTpfq7T9jObbCUb82WnX0CsfmcHMbSYXjamdfIf/XpQFZLvAxa
YrL5jFMzmhoRGKT5orvNqWG46uAe9lvsOwUWBZo2/zGbnNueMmJXZy3zito0W394qNfkuYrlTuSM
XDukhydwFd9mkQohEFbPBwjaT2v3SPJgl3vtA0v8QG0dTLNDB5eo4cuXfvzh98Cyv9y9VjBmnY+m
t+DreJEgyvD1gWCNo1x7hsnk1zf3PzByemR3XljtrQLzq0QCQEkIGSm6LlS1KuELWTlwjwPRxnB1
YxfACLSMW+VAZ/V8Q2dXQpRP+JdLaC4Wculn/a0Iph2ecBM9ye094e3irX7raT5gwrCR8cNuGWh6
1DBF38g+JHEeJ3kZfoebL6UeUX1Y5QXrIidNze2hXFBGccbunjwHDdW7NlWhH+aTiTOHYylnBYSR
n1uEA+7TEOjyjnkacofDIUfM0jIoImvq/aWa3bL3zpWHMG+xbxhO06N6KYXcSt9uk//x0qRSEuwU
AF5aMvr7nsOztfyY+ArEcQxXKNsNGkBYXRSLNWoUpkH6tTUy2KAvAUPhF9zUiZQyVtSUtGIy5K+w
0oeAbEO1R+AivzSqt4MNnszCHtas2/Kbz0VCVjvX1oS61xPzK8fi7MXJO5OI9m5EHs0hbTeG46lV
h/OHawV1q98U6W8+43b8FoxjjAsx0nz6UML/fsAFlJ7wvjiCiJltJ0HgOulBHOrO3rSdmXD/AeuG
M53LfPWY2efNCm4DApg41+8LhH422s37Qx7+mwQsftUwYSzdPAMQWE9k+S/zf5QMJ97z9xv4Hd7e
9BwUt2B7+0EwdwZKh1nqBC3sMfOkNwG66TTHL7BfDZLkfRRygW3YrWVRk53ci1aI5o4JLdrzKlF4
uXT+49wvPa9hL54yxOjZTTDwBalQb/Vey9tVvVPYF/tsYTHumDReLlod48DyZdzFB2MP0YdB4NG8
N/pIttoEXPmmlt1Qv7VyQd1X2H60qILXJhokxR2iQ+ifeLly4ZZRPqZzMcnOap5aBK2yMOonMiQb
y1HBHqLng5cWl5FOfLiVzBPqGevYcMmYVqo/CPX0vSVlE30KzKgX9OhJvF5+gajwYSkJbCEG6J27
rEHvZBWlNTkmZGjvdulHjxR+eXlvGxDkk5m4lmYDlylYcl50rTnkE7xoMjyHIJufgvUlaaNQUvG8
zcpdHaiUfwp4jJKKWuTi6CjzMMqm9fMJxlHqTK/eIZQbJJJIQjljrm4Xcbd9Ih+Pp2Q8aSP2S5jC
yUqK5WZXZ9aK+EV5kgq3/PkA3j8pGbJe2Hz8euO29FASHCJjzYxB1gZYi1f/stViZpXMhESxoXrE
BzHr0W6pqv0ouxZZ/C1FbcGqMtv8xduqhJXCzUqOqmc9cG37XWbgLzcKXiUy5m2/wZT99ghOuOrI
wfWAHvPKvPLrZyw2hS7BWTnjkNQpQVsHdYpUIFTPbPrGFaBQ2VRKciOD1CdhBrtkMdbTpnsxK5Sd
3X5xuOiITQo8frB5a9Ue2XzH3V1r9VkNaJDuoPiib48FkuL23MWifj1ggN3XXaD4HrvpBxbITy7g
NjcbCE8TUTZ1+GMgDrHahrsmI6Vhgy3sv0S1BZn+536xKy1jzmf3yeW27Azbk2zAF0xLE0uWVNCH
Lc+5N2+8VtjU5gKth1j5cJrFaV+rZ33YfzKjsVotp6a79wxWxf29tY21U6xm1rWJZb4yJ0Vk0Vqo
5ELbSDwU7xNpfXP4SCtUK+RQVs22ToWOauseJh/xGCUnKYt8DBtJxpPPBArziM0OmngMoPGW0r1o
6vQ//JgL0OiNNW8IDSomNATfdLoojpZieqrC4dSSV/kvMWkD0CesvNYeqXfd/8XaxlHddp4UM3fP
fiveG//o1Se38k77YSTk0S3qUiSK5+fybt/K5l5Woty2wBB9yP/XRQ5epVn/9A6MyWWDla4gKgA3
qtf5jUvhZ+tCWkHpFWY2PUpPJov+kP8+Q8iaB4BH3xz9RlCNCBskWXPguxqMAwbE81n638gqByaS
Ssu+dmsCyS7qgO82ZOYi0JKypykJv+aYXdYRS570TTirQH1pbGKd2eLPXRGMTGtgjqMifU12Fc4k
BPVbdGwed+HHXaIO92H2+wl9am2i4Xog7nQjQhZ/7bdVDBcDtfvtvpRs27jziPdUj2MAgqC6PHVy
GAoWd+GOZIMMqoHBl6GjSlDhwYAoNe9i22GLf0yq7fscGbAE9Ydh08vnQywPE0xqhd8fFlp7djN2
nKcTX4JDV1DNCoTfgmP8R5bBpT+qR/8YM6reTEP6B5oN4uIX2PhpcxDXUXGMcjWwRpUDAQP555dg
+m1vvnKBGwaIUtSq6C2Xb4PnZK8vt3Y6UJhvOGGJe7E72XBxTsAlbBy587FcdDHRUATPXGLPuKlS
XkEKBQC2PhCSgR1TMPa22rtGEkG9uP+Aab7JYQUTqzTqPMmz7t1fjWpCwZLlxySTQOBr+UHNERDH
cneN03KnNQqG3m9R0ni5p2VIhiWlEP8MF/FA37HfMpVtvkoRK1H1iZEYxnIWPqjjYlpTyZQ7dJrG
6f2wiBlRyK35Pghjw6il8+Og6r4rbrYGn2/I13AF+gcKYvrT2OSkmm2bGceTsxwJykjF+sKGHTiQ
Dfxjzj79E3LjfiyBpL2sbTGAvFUsK4fBVXWFn1lkrcYhmEvCU/s2+IGMDi9ZCv8JtA4MwVCsB5bJ
jmOzwX72rPfvBfDhQBemfoYk6HwgxEFC0/NArHmqsXWldStuuWEvjaLIbpwGuGqIGJenSnzxKoJN
NydwsBK6GejMCXKPN6AHzaKPuQXXa2IM8sy950/vOSr4TveYJWoFI21yx/Lz2z3B7XYaFpoi/3Hh
7l3xkf/rIs6NKSQT7OUStk2LDSq2HBjUJ/kRYeQLbQqrFb08WJ0WRzw6HRKdNHIdOPiGKOWOdFx9
P90PuCKTEdw3R8k2wZ6RNB38ZlUdJvb6r7bep4XPiWEtgJZEB0YE1tE4gvHqaiwMbgIXMQigBsDB
ZlCyiDtCjurK9/GGlk7i4bSNgvUInIcN40IYmVYPw+i2VMJw47vbp+h+tQr4GrfA04h65kyvpXL4
MF9OazGfLuxeLTsz2brRbEYK/jfVVP5HPc1VMYyz31RW7AOeWhBJGkW9dccVmDTJP84pWzIfRVh/
Kz9xVa2wjgo9yggl43R55j/xhCUHcjPP4bS98pYJ+T3LjOZyrRaIpZCYbyXcGM6YJTl5RMWFqL7W
2VZ7yWY0krvGpe+zU5Z6jZeUhfmhTdx8ERZaUkVdB2ghyhBKsFJGJqA7qyUcWKN/uowJ1qM7o1UL
yp2maRUIj2ZdhGTnc9Fic1n7+1BHjzxoNFKf282YWjBpj3iGp0SkcguaeKdvR/x0I4+zO/HNP61U
C/NCvOZErpavox6uGmHIvuwPpjtXaBJng5cNeXIrgonZnROyUwDlLY04vfP+AgxGBrx/tLQX7G6r
Zx0kfupZs1kRlbdMl8f08HkabJolJBwUz41BdvAFqWdkP6nKb4SArLr/R5h0i1GI86ocsRnxOmze
2Jcu8DAXdu1HgZ3E5wd0NPNTnU0yocJUy4avZg0ulbu/c1zHmS3/Vub0wl9cu1Se04pc1E+b9btY
yN+2cKMFIoWaDA10XyTqr13SdIJsWlZvRAbQgRPz4ByLNEkxriha2LOLn9NrYw3sZBeejUGiTxst
B53hzKiV7zO7CR0UsxLWJAA7dxOM146cmiJmN4ITRUtgLh5gUO47HXBl3otnHB3EnCfu/I2MT/ma
PJDuKhTPQMzi0XLVJCCQqTk2GIKs8rxt8lEc+KY+mCng76GVHIlvhqZjG3GeUsp1/X1XJ+DVk0ug
0fFv/GvCGAqzAlCTH1wMicGkqRsE9kRa4Nh0DPqBUSRYoMRKeMnVpEufB1aOkQMe6eGXR7UxBZhX
IvjQrt9HZ761wx5uK6f4A4YabFHFxTjMfpQ5cY4VRJTXSA0zL1SURonl6PGbYmyEtsiGO9cjpLDE
WN4cu1ANuJGNNS/6qSGGpoJQcXbd7KzzoQMaLtWgS4cOZKrnSnFAwBEgO0pOLzO1D7IP9o4odX+F
cjBaQDXZRMq8TfzfShTvKdLCzg8VzKdin7K+BHAPSrLb1P4+3vaQAOYH1yU+SZjAfBQKnfxpd3Zf
JJXGl9Bps9pCn6iBZ8SEtGW1po/p4kT1EdqVffYTYVsVku/KrStXRm7Win6WtNVr/7tMTon3H02/
Miy6NlQFlnvdzva/h2g8Vtq02edZYw/H5ZcZ1EqlbmDDMRtFFZv5EW3s+8tQEKt7WTznqibpu/uh
NjISx5Y7blIHYcsfNj6jav0rfTqGtu3vGsdegfXEa+CEHr7CUMoE/m+houqMgVut88K5vkmt3VdL
9VS375mDwGtZD4StF95z2hwhFrKnRKSJ5eAxOXWscWGJhLT7wQPFl8dJNq5uJaGjex3rHetNbSZs
L3dLiIP3ZJlpvQfRtw6fWUkxNQxC511Z7+4osjQ2vJwxJawL5qlxAXCG1sakPMqqVBGaNdiFujkI
IgFhNL/gBXLmMuH/2oaTz4+UH/RiROnTPuZ18lnT6L2JGfbAI7ZAzgslSZV5J9UZ3ai6uh7vJv4J
N0vqg8/Q6OdCMP9NzsGcZKoQeH5CBhxlQ9JZqHw8GJjS8MYQkQLfX9yr+YSo3m7tg1W5RoMLb4kM
ZpQ2mbNnrR+kQKoGfCRQDJR1n6dmx5nuVxmqYF2MMd85b+RZYBg8R9Tu7iuaBqAoe5NJtBK9MGmM
DjVtahBGKWsxL5Jz1y1+qgaGmt2FE4zdko67rRdmoN6FvyhfqdGLTK04fMl7dvvWuGRSAHyv23Pk
H149lt0hWqqHty2KGQDsHRrDD9VMYUeIWyqnOPPHLGwv3Yt2BwwQW47DNOK5JPcdTMZsUUBBXJu8
S80ek57blWPFtrF7zAqXts3Fn5z/UuAJ/n5tnICNYCA8jckciaRtjUCeMEbvnfyXS+SdCRCrncwG
SezCXRnCfvIrGnmo3fW1KP72KzLoQHMAArtwJipN74oo42Cst8volPNES98PvUxEzc7yOE6WCuHe
AHiHmKT8sM+hBc0oGLjDuCdF2sPldPS7glfb0/+/E1D9WhsjK1Qma8XFusXlt4YDeSm2jr1LMg7z
PSQgBrsaisngW75WqFNinfoomfipcxRMHdsaoXLdyqXXjqZ7kLwSz1K7ZK+cHw4Kv0NKq8PBZ9xe
ZPglEMPRyx9PQkBCNqohe8/7Ld4ZQWxB9QEBcN788kuZZsYBKLCICs6biLuYdF+SXBUq6y/6HeM6
J4R1me+MislSjEixIsli1QuFVwRiDDgZa1umVjL4xF4HO37KtJKPN/9j2rqsuXtA2pCLzZbkhoHj
eDyiSobOlPSEdn1nOl7fBWSwV1CgjDSB/a9esGYXSELYkccl9ztLbvXdGHZIIv4lcoX3ZsY+kNHw
kd2JZZZctQfMnTrmUP4/ow2sl3So/jZHucRTPVh37fRIO+mEVUBJ3PJjbU9ME3Ta/shiXY33gkON
0AZ72EXK7pLFFVGGingSisVcP2jNCIQZkG42OwRL2nZiUQ6nMBngLPndIrX8JCSZAo2Mnd3vcAz/
NadDMWukasYP+negOJ/z38Ri6qrtSfvRPSaQ14RRnL8aqMCmSd16/O6q14K8a7rb1i0iUX2ey32M
hcnYZzGJ8d68vSycNmplD8xEoDhZuE7MxxrHMTVhNpSI6Cn8jeo1XLLVJ2etQX063CFebWdcBqZS
FwNHqlXmcUIj6XBZfgpXTZud9A64mDdIvup0KdHQNzXa2sbXy1St1egRB5V2eoPmboliGRcDjO5g
YLFvjYXtPZ3APqYyZS/pMF/LyDiYX5QlO5QIjyV8ABux05sOYr/TK246GfQ9yFjQG9+rAJ0Nl2T5
aU8sooa1plK7M2s6he0Rqcwp1vuaAal8F8IShd+zPtfaTrKnFNE3897brrS5SDbBXRjbO43QpNEv
tvnENvTAu8xISRTB49EYj0Bw29GD6PZt+y24RpZ4KLxXcyFGmrjW5ajG32fAK5wsZ2BcMs1ayM+7
9M//gjF3edFs707mVo7/pdi263OriDxQXIQwZf5IDy8qGNMdAJnTrIV/bY/ImCys51MkuYC7P74/
scxxPmpFBqf6tXhPx/DZzIlYetFCcIJUKvY6gnsb23c4y0w5O73HT5pytBqkeKSXzvM3Xyykxaid
MLbhF5tAJLCtP0wNIsaafBtg9Q6liEjVItHV46Kw5VBBIKVm/JC7BEEtcGj3IUhGkJ84uLx9J2ZZ
0HvU9wLcFV94kf/UP0Aa60p/Ze64iHP8+/wO2VUf+9lNFcCxiTzyL0PxvwfbIkKUOhEbWQasAMMq
jVr0zuR5TCOdaHtPI5jVeniUQph815Ai4GzY9zSkQjxuRKW83Ks6cnSSCVUu5vkhBR86yISBthWY
HolT3ZjUHaxzQLrHTtHGLSsWejquEiTK9D4z9k62Leuam6HbYQ6Fq+6vuiTsBltSx2MIA/W8rAVe
lW8siFDrhwAFYEYlVCw9P/gZJ+TIJ1haUuTcRCNWFDufL70WKTxf/RAQlyzmp2wHgl6K0cjUpcSI
JrDp/xqRZhJxZ/fRx5ImBsfdc86ilQhkWp1aB5hffFRF0TpLCf80yhAPJ2Iq1RlB8PLNuRyBFlDf
YpxljbE2UIXAnqFeolwHewEz+GY/4NlSXrIQYIW58lnpbUs2PJPPCJvEoPF+t8qsUrxRhZHyLiqp
5Pf76KMGFFWoYg7gVCB2NRu45iBK8gGn25Cxu99wM3Q5wyCYKkNQ8rjM8Jwbpmi5IS6IjyzziX+q
pVtbVbUTUCH6awQlU551/YphCtuSD4+LioSUZsndxH9rHT8BEHrYuUdOsPRjZfVQxcW7yLqDR4Vh
pDW5dyujWFNspJTEM7y2TVoJfVomF32BpM/oj+yh4/ray1yTLotrz2uga7YHi1Z5AZXkegGDaSM4
96CjU5/UAcxQ0lMRKriKPVvWp5ew8bQVIsCI+2BcM+Kdc5AkjeNjDFMN/VAORlnILwfl/YVrose9
lJu4ek7pJ1nmVry95jV1QwE2F9GDh76gBrB6ZcypSBhp7LF/h/4PMcSZ0XPUqY4DDy//LvMyOlur
Ecw3AA9v/aEj1alVOhIWP1gCdZR+wrwJu9O8T64NKbZs5fRCfUghyAos7lsxZr1bhLb9opC56hxw
VVl6gaeh1CVplj/WFQVpHXBYkwLYX1NKytyEm+doOgr9osmFJ//5INvuBV5BANjGA/SUgvimgrTQ
Km4By81lHiundGrLpoNEXBxmX521QSo619MHz3NdvDStSQuVp42/OUP/kq4IWZ22IfGSmrNmG/uW
+VeWfrPBlIpXyZRdQMcZ9t+HJgNo8MU6k+EhQDFjF+TNzdEYxEsUJCliHTk+PmkgMu/3E+oWbLzk
iBNFPGpEYYFkuJ4A0Qj5l1A5eYL45xTrHMgKq87JEULjdGOYltu2mnvKu6J7CjBnzgRNZ5I8Dcb4
6qNPa8hBRV6382ICr9HeIfcFZX3uscgTchxybBj9uXpMWNbsphYDpuzypkLDlhIwvNBoZIl90fXV
DXY/ck8GRvRAjOTPmApHW8NUU4AjPpbrkVk0bi2uzlGx80j87+gBqH2thCC1ptl7dPciUGpPHi9j
DI7g6tsuRccmk1oVptqS+0lqEX+87MurUFKXDu1iofYb8O1cPsnZZmPRrmiytiVgUpQP8vsRnHuJ
05M0KSYJXA5FbUHLp7ZLJO4pJpW1IMvAGBTZtK04yRfyERRc0we1TlltJVHwoca0mnAFDmY+SZGt
xAYjePzEvF0BkQg916IEHIKH3tDlcbPtu1k9E63fRd0EJQh+67EEQyHBboacxVZHuWNoUPKNv2xh
i7WNQYV8yGDpQZ5i4KSQEdEs4aGlg+dvPl1lgvTd7Cs1TsWeB54o1IzQHpQ5ALfyIOgNODNE1+jT
tWsSVgwpqgpRH8x/ilTqNFQmNDTf3qqQTd1z3S0yRF1TtjuElnGRtTM1EOwCSZ6/aC/jKjAQ8jFR
o3V9ikMFuBgys6wGNDc/ceJIIrcSnhH3WDSEDWI60fwwXCPXACDUT+o1jlID0UflUGUu2LOKHh6p
badOTTCnZ8i7UeYbapc83gYik9sfnVz3pTQf0ozF5/QvrSt4zoa7A3QYgRtv7xX6z8CMMBZwczf6
qXJ0WbRph6SBUQOGUkDPzLpqIAoNXCrwovurub8BCWbrd2HxfzZ93UB/3XYYs+fkedg2vpRZyKqp
FBAS+UT219U6V7aCggd9vO1Tc93x7URHcsrgY3aek8lTIHiHergGgSt7hibhPzUksGZC1Gfm5Foi
CPk5LXjvJRBoudIxC0k6bBKdmPE0aSDY7HKNztPf0ev6JerTwNTwytA4Iu9Em3vWA+NdlyYQCCAj
G0CRfxWxlCY6px2lgxLTByjCXTvVpNEQEPCEo6rBjer8nk3n6wu28kEjmQ1z0XA525Qc9hrC2LBG
+6tv1K8FXzkVZOkQbu3recEj97yMPaXp3jFT+aeRi2h6hUdmlCjBmQd5tg6byJX5ayNeRaa7h4ja
RjivVh8W9mJfIu7W4toA6HyC/cnqOrpYPE0edFEawrVSUWpPJLnNoKZgrnWHfs5cSiM0WAAnaijy
GgO/ghbdg58vrkrGhhMJ+cE+3y+tMXumubd+fsH9hyoLzgz9xXE0YXgXXGkyDYoy7G52ACioxff0
l/X2D8xLEK68s4Dk155lveCDI8cLhFRFtdcnUPsGMk2Wtm55XX+BogoWJ7YQ9XndYmWG9Sw8fLIA
sUF7ufwtvafoWZXVBEaclkncepFVbbAn7NAYskimY8I940OWberO8qYQeC3tz7SNXFyYwMDDFeRr
Ewl8OiOGE7JRvT+0ut/vpt7d/VO0jxZjL/Zr3SpFCYsNABOF9LZXfdh09QKn7cfj1yYRwVFg6CJ5
PgAQS/Hn2zlOOMUAczyjqR6DQ96UUBZ2vzmYV1L0MyuDUyu40KI8sP/Pjw+WnL6afqcwr6PwH8hQ
y9DdF73MyyJxMlxC6P21GREhHZT6+YLIQvpcVsUlJDxC75A3R/QEZmbbQWS1WDzNUvcldrenDHMx
7q4VXV30VKp5omrszD9DypT0feeOeQQdLvldC0NUxJxfRNUuCRGcVVcbPm1aQcjApQfa1JLlGex6
XCfOc21qmn6Qz2FETAhRaYu2TEiWJU6DMbSYydnD94+7Omk/pHh1xtz0qnib7GDIj9YvnFG/gCCG
gnClf5pi7OesW8yMIYwz9qMLW5U/6W4LuL8IxsLl1m6LpeS7hgmlOqKibYuNEPX1DxH0PoXF3SPd
dK/hi0uphJnBdSKDg8YUs5jxlhIsCal9oBt4QOUorVkAzbiZyT6Pe5Czngs5iXvHjBcyIebh6v5f
PGQLp01XRTNG/1OMFjUgHwtc3EOLW3gHJ8O+68CerzUIfEOwkXsiklVDgn18cXC9cj76pfRny7UE
m91Nnm7ovs5lvSZF0h6xHpR30fHZWqZWKU6RSX7gWvXyZoT0vln0KFwh0/Kc2BiohNEEo/HtRhW+
gd75B66v9OaMEhjXcgOI5nsE2t/0w0NEzxC6/M6uC7BcdLAWslp7TmzJBoC5UKhlf/zqBLWDPnLl
owjXNHnV8ny/cX48qOiOyIKUSVRcVflp6fcYHRyCPcFa4Hu8Kysk/WPpZAdmCI6cHWBOfoXgbXDR
u5vuhnA/svSoB3nO8Tvmm/VRs0kTXcU3F7OXzhVOQeBxV+tgutAQKjfLfZOe0kgumNo0NyiZtyQ6
qmwTKpaAnbwWq7u/yasoCngOjkeHZXconpTlfRij7B7aDhgaVT+9x68JXkGXiGKa4evRkKrzD9iy
uj4AbKQM86CIIxV30yIU0xDhB8llsTmDqUfnp0TsMHrNrXVKqG2A8JC93IyDDQg4edo3N2lX42vD
eoP8i6azKJt/7p5+AXDDoQHivdsSn7q7rgV31OqaPkDajaq90CuTr47ARqH4pPVaPrFypQJLxU/P
cKm4FnSjMNEHDhR6Oqvn1fsaP0rxxFkut2gGmeAU3fIgB4BU9Lu6w3KOi06pRNw94viHRfx7p2hz
IlkJbr7cgZUQkBko3Ef8oOOXFNAJfPSCUC61MmJgIawrg1yBdd9HreTbrRSPH59ZrSXEsIhUR0uc
g+RZ2z+olKnGll6fdD5CyTBpgWVi38Yvtp+52dfLFb98AHtIJ5B91I9/LylYRhAiSTwnn4INHmAE
WhPIErnly/HIt4Un5kdxgtZ96PyysJAkIjJoaJGsohkasFq6dz3jXeAsUJWhxZt4fFeTI9aVHKP5
T8iYNoT2u8SBp0UK7xbNbZFbBVRuF24EzT7D30eb+I+Ci9MRphcxjyoJcaIo8TbzcZGsd89YYrNf
hzH9K3ff1h0eGm+K5qwa7WqyOoxWpCjMqxdMtZpWAb6p10AaavbSfaiTT5Li/iQcaEnUT+foX2pp
LLljnRoeiIEbKtQNTiuL5n+lYDvFzX6x3ii+mm1Tefzcyft5wVoU65M4v8qDQOuAeMdL6O0QTmqw
I0ucO7yctEFYQYJd0Nf4f2ppA8KywBYAB4f6xmKutp6MktPMJWfzeM8xnbpbrwItAnh1AQX9yvuW
co4X2wWvyo8rsMe+E1MrschtiVPmW8wts+NRLOJ6SFMlDxk9vWtzRZtOc2HaN5djF0TvnYolvVh4
AlouGtmEgGX3qrDMUKFuJYJaPCwP7Z34MaJhfrw39b91g79WLp8IT/PY+F380orBeEK6SuVF0HP9
GanVK6tJj193MfDd2iuSvXgoJy/VbZfkvsdKJT8lEs59kF20aCjiOdNhZ6Pw/AgqNL2JwGq49ncw
2P3hkbaF9VH1GsJtVgD7VTtivRCn8PiPqU850EvQ/OFog8KY1PvOS8YrmqKcGD1AO8Xm4nYjbUW0
/B3p+nHu1w/IXZPUCOr+yd9/NR5DLDNEuuJa4BGXJXSL+X61g7px9FGOBSjNSLxPKOCUT5o9toEF
5kyg4w80IfbuRhujRYDHMDRQxfCsvfk4BnQlmpx2uyDL5i0CUUbJIRzU96MdSw5czc+v6ryO0TXl
sUv0BQMAARqSIlzgf9e/0cJlOivFYuWxkz65E1pgRhnadYHdCSWmazKVBKPQxxPqN/v4ng17hZ8N
7juO0Ma6MKMPfsHq4siqMJsUN39uccFXDTenlheDsJO4RodDxgJsEagKI3Psm8dRnkGknN+ntb3E
+fjH2JEZPH5u7k3scOLRXNK9SJBtMipCGYyv/oBVtdqu2PBn532AYXzgPGoY5jH6rAvFIMpVTz9H
yTZWbnHqDlmhFQrd06cBaJO/p19VsfV63te8okER1SZBTK0ksT/YYW/nDldrov7cDh2CFbGJPeGI
JAUAW+A+WwsaBYdR+JpteJaRzvlBOUUR4GNODOtJlaxC0rkMGL8TdkwUolrs59mS2q4b3NzES6vO
U65CMdLMGNOI1FarWqIVi2NYsOwlKFub8YLkXi94pLeWT75xHha5LeWxSwUO1IQVeXsbgpyJyo5Z
nxdIK1RwOodi/cS1wkdllNl7BN4tAYfD5SWNzbnUrXsPHZYy8pP01SIYBodot77rK+wpJl4U++X5
f8MkbIUo8qdsACzlBfKxidApHqhN18JN9beUPh/YaIoJCKW0F41HoiOnxiJSkeBCjIXbXy9R2m2r
QPVXZcBdq6voDJUkM8RFQ6q8wN71setH9ZB7YwvnXudHBtgqKBveUrsaIRIcLluoYqJPhG4Km6Qa
oRRr7TvgerLqe4xSZlPvXMl5lG+efVS5/Vk1SwSssaoyNfBbuprg4Ko+HDtQ1F1BJeHNCDbXQI1p
BpEYkmSDWI7ZFYQ0JnxaSFPcrpxzXNEAAxdVt7TgTGuFR8cwYlVkilB3fk95MtW/bWmRq7J33MwC
joYECrDMLcF+eCrtUJryT8uGOezd6UxfuAqNG0Ss1g/r9hdzioiHz8y+DOK2gyceD25gurC4J/z8
O7o3f7ZDsJbJzQb41r0mBnyMl83nUmCjEiombpR6qm12/Ce9BgU2YRQv1dsnMMvwSFKehLDABXyf
bjSwQlGhW1X8/fKkBRlbJeUPMj78h8xck5biJfZE0WJBk3zfw0m/+NaCP2ro4VgivQO4IZy8Kxkl
AHv+mZ4fDG7HrIIEdWL1V0eSt23DlMUXZOOrePXbLl4dleDM9GvAS6kSICoIl5EX+QHyFDf+BXSF
pXDq//ghrIfi0QBKy7P2CYLLduezqSuzyRxg/TdaP8fpK9Fz7lIrv8jhYP3ECQ7RqtUqKXtYP8uu
81zIU5jk0iHc/F91aTleLiAd+Jq3tS9BQdeXXE5lG2KTDYnMBXjn4ggLkDnwYwljkTjLy8spNddM
WniNWVUhdtUQZ1YdIRD+MTObtcgpDNOJoX5ZLHU08PBILXxy2Dfvq5KbwK7HYH9Pz8i8Bqk2F8eV
gj4yVl+VMH44H7FF85z2fIbWUUatZMGUkEM4jkkcmoq5WFiKV+WGL5ZJ0kKHzJ1CcDKRaH9k5cqY
MJeyWZD9SPvsVHmhkDwQiG7rq4HaIBHYww6XQ/eQ/YseyOEjeK6//ybyqFQi0KdmG2Ihc1nXT3Yj
3o4tce45I+Frd9t3konMxY5ttq3XedOKMIbXtTnB+3ZqRfMRj/hK2lmxlZsZBIzHD/xgLd7EUtc/
LVEY6HraxehR7qeJZUAsSx5CPGb3fO+z/ut3TjwWzrv+wjrAasw1T2u54kDBZ66ziO2GU/4K9U/S
QIZZ4v3+s1mXpyflzAmjSf19+3SVQFAbzzP9cYqX+YH/rldttTVCYUpThUEKntiCEqbN98K2oBxw
8MMVgxm1ML+zDGFRoREOPItmzKTRkvMdXtHHfBJYmkpWIvW5ypxTSGVwH6/PnA2/Yy1+5U9wygQI
c07+MbaYTda3XkIPeKJ81zi1SyfcH6CweIuyfHXDmJiknP19VClrkeH4Prn7LIxEUcXMq5/XkAD/
+h1s+apMBbY1pwW04suyl7hrU3dhl5ZteDQ1N2hIfM5uDv3Hi+p7TPvA7ScjEoho+9UQO9hbs3EQ
lsMYDW8r5Cn7PS47vMkuOojz27XlXTAFkikh4KqaHaxPpmUY8F1PTGGhxYZb3G/2ZxzbXMxVbk26
NAIcs9aG2CVvHNWz//jw7EW5RVuPKAHAUtFiuo13iflaE9GSV+ssCpLBj763egXMtVI9IvCcqqsW
dPA2wGijCaKjFX0zBGWX6tvKsL6gno/mCNQd/h4UEhsceP+9LVEsSiFJwCiO8N1UxZXa2mvRL4r8
sDiGrB1kOVO9If2orhOm9TG1D1cq2rJaaJzq4wJeolXbD/0J0oDeQ+v6Tm154CnFSxNaRaPtO9Gs
j7WJWK9eNPkPNmHbCebIR4BtUAB65UL8uXUpue/GehEMj4k9GqUSsLdqKEd/RL3OGcxALLsXyddC
uI7sXdkdWhu4wEZvsOIvoebjW3I1HNr2xWiBq7FRtz87cs0K3DJkddCI75IK+2VZ4Xe5KAWGXl9b
luEkA0FEB8eF79rpLQ8eEZqXxGnD8350Ykwfb7WT+/oeVD6lM5CdRtRwIOTmhVRqf2Pqs2TxMxFO
dss3gmbQllDL4UNzjNHCscfzJTud41NQeS2uVKIqw61mjJTYAilB8W+ZBUuTxPMXomGToQ4g5/WI
GkLKPIAVMDO3RYXA90snEeOBiR4L3uYeZCf9RtYdBS6frkgyK4MUt0i+OUa9cO77AipszHI4ACO0
cVqBXUdigrX7Hre306bf0NmnoejetuH87U0PW7A6x8CX/rvWB7K7vYKPw7gI/NLk0qheBk6QeiJB
z/HnDRxcTgZSpQX2sz/kSdzjm4ao72jOGqFpqrgtmjEM3q4AogmJtQOLZ1aPQs5CEmbFjt0lUZCa
RlWfUZqXjQi92eQx83a0PuFsMiz0BGGVUdl8Hf5iaxuFdT+WUtpN5VisuHdtOVbjyvp7IsztQSyk
CW0LJ3koZE6YK9DsMP6wp9dBaE/Y5klAxE1+fq9oYbpjAmMXJo6bjp0EXFKIjelTCzeYxSdw1u2K
kWr+ZwNwbKcySJvxQ5UpT+rXjQPmShFpuMoyD/Q6vruS0DTRIpWrg7VXDjovTTBlPJKrRuDjLmB1
G4SDcczZ2GaGn4bc51BiW4MmltBzDsz2yjMHyMN3i1RwlKkxtmvNwL8fE7ndr6qAKKNqNdKWpR42
2YYRWVR+qLJudLlFOMwngT/fIWLw9WHJ6ydU7eQtrvmfHzyU1j4WDko+Z0jrZRgmgaVplhmY0r1H
o6ECjc82NyT84maXakexYWKOB+33h9o345ck+Zy9wIrYHzltf4P7pgMt+y38N6dCJewqHrzKw+oS
hmggCRXuHSNB6a4PcoMgQQzzk8cKFyXlZIVong2r+yZ3E1h5ILqjJsvoAdG592WjZGa9VPN7nX8+
QeXbpZXV/361yT/bTPmV0cY9zn6ifXOx8qfrqn09lH7Ks41OOy7NzNfPFcRlN+A9qjeUhXu6KSVP
plxQBIK6uGhGFESxSAlRjjl6Dy6TaPeEY43cSBCtkcddjvc61FkanD7WKsjCpY2hd3VrA0Gz6hwJ
eB0J0kmntFv0DunyD/Cq/uE7R6HGaaf37EPZn5ameO3EqISZSF6M5mccx4A2Mpz5iQqyKC3lMj6O
TZzaOGxemsQHluWGxQeiSmYhDF8QuTqzBXH7likc8O+5dMqnd0cx+kUu5D7hGy5FrqnwyF7EWnUl
3JusSo2WRuAAMqcWnjcafiWlc6qjYTrFddS5q/CGbjBImvXpzsFxLdf7JKJPue7wBGB5StfuEXE2
b1FUr9hA6Dy/B1HJ4Yj+xvPUFfy1Jw3VaaeY7mPoDTtsCGhulLVeoWqAOFagB8qwbwvr/+d4MRiI
ZVVjoLknKVAtrxtT9nr59zkbroZ1tLATrUuYhVk6XrNZSvor+vE2vhZMEUhIoLLTGZRqvHmQ7hsu
8BHy2Ky8FlED1Jk7Xxnt1LfppnkdYWuVNJelPYODQkWNknR3SV7IUaErNvAzadfsuBRu35XCyQ9H
EG2377Rp1LSdH9UZSrt4o7+nJZdwDzq8bNtY6Z/evhUzurzrvAd7U5X3wJP0nzn9f5E/Si95cMGW
Hkoh3h5Z7Ca2Cfc9TnOtwEOnbubG97ktocu2q/pf4D8l3/tOS4fMluWLQe3QR9nXS0dUcQrG5cM/
hqsqeAX+f5qucfplakmYNZZ3svlO/D7WLmgPrB+MG3YIsyC0VEwB58A4ztDxc/QJXbg3eMWfQpuF
YLxyp+QfOnNUyBHQvMfpLbaES/GXpPjsUAPs2XHSvHOXYuPGwSvMZJCXjPEuWoDCG7dx3pvkZPSr
innj88962FB4gRzsgsT8ZFOm6SGOTEcAQqJtVr+0fJKdyynIbhmdLyk70ZFbWgB9kx/mHZcjOW4q
Du9qr7Ez5KIVph8+uUf+sISFOk57Za0syPYsROkSRvR6aRM7E4xDFIGstt1tzVC79u6ynYqQ2ZCV
CC7fcQbk1PtOO8BKkCuaN0LEqI0SEOwaFMFqYK9FIyXM5qGxqToNfvpB8R7Uvzl9KUnNFLraHuoq
6/G4ri4Fe2GHR/TTFKfziLuWT8+TLTseMvFsw8nMVMenC2JPyDm6Cr7X9NS7tCFjfhuc468XCdOe
ZuVt3g2Ls+KEuRpszx2RI1pPKxR+/eWn0nRR/T0mzukeLrTcoHT+KddUKWhlrcXgH7tbGUha93lj
m00gMrltHkFgVh12brn8YVdq53v/zDL9PBc/TVex9NsxptPOHXaoQNbS+Rzhi9TojGokJOwu+vnS
MWEa6+y6wj0w9kiZ+JZ0EmXRSqbUTo/Y14lLiiVNsX4EMFbmV8UVoT3aka8jt7Uu51Kb8ttnco+D
f9UCDeSXpWuxbmfcSkoe5XncWYn0k271bvGpKcjfz0JNBQ/h7S/qwgvRxDzhzytwRseJZgRZQKxF
e/hgEqnaXhVTyFzWiMhMm3L1reHHrW/zX2Aq8S1KDk2Ew0LooV5el28ZSJMs46opozyA7bMtwMhH
c+Ek6Eo80FEXL0uN4hUP4gk3j+8yo1SW4qc9oVN3W48Q89PrMr5myWrFGPP5dB683VagIIDwt7bD
EGT9AV6Bw3ACufF1NkPCfOPS9oEDjZ7qPuQyS2VwIRjPSQiemK/l2eXqLBoZswTqQ+xO6AtEVJWL
tLJY3s+nl+qgLKpruTsHk1L0waFDtp/hcgo6ZwrNgl6ACpfldAOURj3OauZEvr1c27FiZVpAZCM6
XkVbRZkbFkHW+vLWL8Gqni2vXoNUv3dgXCry1zpy8T6PxKhv25Xp4tQCwyqt+j6zsM9PXDE+OZX5
oXHwdHV0BwXM4vCKweEmqajClYW3kyyIc0+/+TYEbMGuFUgXCfYl2DwtCsBPRfzgTL6PPdF6vPK2
tYmkaobG2vc61m8GSwMvLdBfO/uODrkvK1vfP3FS6MWVOYSUome9L2E/QzapHbk8euzLOe9lzmVp
t89Kqf0qFv4zXZZ7MSJO1Uz9vRA26zOEUxF8jBLgkSpH0BA7UmdRGOlMohvAsSpo4xjmoGJFvi65
8s/rWIqgWcFX8T+jDZAMEUYjwPxh6PN1GMrnTN6ctqaRPfhZRcflxgwYPIyrhnHgmzz/OZOb7AKq
B53KQ4f23RpOTeV7bbqDOeaVV7KwzcLMPdRebmKDAP0CoL+73iaVGxESXWwUb/CKHyYkWJWwR2lV
2GdVDsIUqXNv4qzMq0Mow/im3WSN8A7NZFLWxFRtdJDeRndm+I+xsc1h4e4Dhlcqdsy5o8SIKsdd
984Gj7mUAx+QupAIz20d+8ij2APPyYS4IajENz0DlRjoPSLlzBb0mZS6I7yXnCESt8QDs2LFXaG5
xH0XS7/VYipp3hL/7BWm8Et/a4TM9/vT5gu+HlOjmAqM+wKCdcwos3khm1a+a4YbB0AqdlM+MaH/
cUVLznFwKHkhgUG5z/F20khuznZRzZ7Vnat6qcySR1DnhyjPEV1BDQFRoQ2QZ8eMNKFUtxrPv2JS
jKpSeB86shLX6eBokPGAxoZLGKOBluwdDKnQwn1rREqsepkpPHwa+UxmKTsvzPf7nX5j34elayTW
J/Tm1JVLmKX8qOglWBvdN+au4Y+zDa9Pbmn1Uk+39uSu1/y5rC1Jh4wtqwmgxClaD9s3OFd4l4fJ
AjHmAFzxrQ39ehcLz9iJG/NDEsv7S5X7lywmsQIiJwgtyLzm1e1CYg2b51xDnpGFcbTsJTeHa0oF
tFXS2cv2/7qeJ830gwUP0oitbCYOB9NZP2wGeen4asTrdG3917G+Mbt5PvBhrk1AD307BlUQYvJ0
N9fsCjpAJQI0JhUiRntC94FNZrrALOrOV13OS3dI08h2loHhO48QikMQuc3o9Hk1Nt6Nj7Krta4g
1ACLApZGB0c9y9ZjbnFaflsG33hO6Dht+1E0N0v2JgUn0p6FjXXfGq3OGfDUrE2eUuTTauXzBe3O
hGKvZDJozNGqJPu+ACwNUWykmHVRKQ8fTy0Lw5lCK4KgQoME60D0l3wsuxIYJxpS+r5eV+q47J+G
tCBSdwnwC09GrkvfJDV2qYFLCQ3KV5c5YkNWg5YRKYwie5ii6VtEskCZoz2ieYakX/fqOnxR7igR
zgDXSG+RDs18YNbez0oCUsUIwhVHM7aAgSQ6Tn5qRP0mrdqAJKjJ8/TeqwsSKEvhtIHdEdOn1mvN
zCDZca6aFHD0vPJIXgnB4NhZc85R1L/TfrsIVZHcqn9fk0mH2/mRzCtn61VCH0JgsLMH2gcyhOkk
PAQ5pcSCxNS6TfS63OyVbwCQQpndClmmGNZiuKIli3ywEWPkMUT3FpdPKRuo6LMgWwEAvT6sj8EF
0fB8+36Gl3GGS5wrszSXtymMk9tRaRkqfglO8cMPpyVD/XZqBQ9hBW8PM4tdMfcXFJchoRn3NCUu
4ZmZ0mEol7G+KQ4JXvwZCebhPr+QHar9t7u0OVIznT/Bfxbk9mapQ+PRR7UrhtEoRUk+dK0TTsGi
ibILcKXzOJ83hMOwHihFUujz88p+uvXNQ34xE+b6UhFY/ih2UQCxiZr9xb4j8ca+8O8a0DbJ5jO4
nzv+LSYqkdM62DR7U8WQcIwaBv+Y0I4Hs4AzS+NwfUKFxQPh2XLC/3DxXGmmI47M+KAxk9MJbfZV
4+rvgVf0rJassJr6+JVQsWCy0vhyr0MzCpY5yzQctWUn3Er99zwh5TTNapvVXl6wnxpCZTPRbMfE
+JIH8Oa/yr49PAYP9NLMAqZYNOpsIU4jfweBXCvoEMWORozXvBfvFuJpCD7yMh59Rlc5LtDh7o/J
0UUf7uGkX38bxbwuRJEMWdz6n+idJpH8a+2ZQTl4owOjH+7q2I1o68zBdA7fx4QZPTP8bGyaH99Y
nFfMY3g28Z0c3h1NhBeSqmL7+0b9SE/SIO4j/8k4dabcw7DXh7Oicm2TpM58/bQUOQRY7SHhm+ru
zA1dyzP1BSQP5tDlgGRsZpFxa7f8mGQIjvpisfplLb5P+ayXtCZ2S9AarCH0F0UQ5VddQIYD0GJJ
vKpEIxWGAERWTss7AEFI8WeGok9AYTxSVS940m/gyfpw/HaI9gzGDWB0lFATTT8SsvyHfe7NFRHr
vknBkh+ESPYfVED5VoZjTxuGLJdWOOsL1za21YuJdVFABxvP7VQhNq6IJZra5P440P3pzvu29zdi
ia7BIdCY6poSOg3HHWg/rdkvlbrPKMxmlnNKIG7WuUh3sihRsk1E6dZnWlG85sX+T1fGGJC807KZ
qeTsHSt3UOyO3qwV3/VmqhA3Fy3u8iYH5isHH9mC5SaE8KFkun5+5motDZeHm3e/zInk7ALe0gwp
b4c78GPgHeQ/Hg4nqBJ3BU6yzrVG7z9o+2qpYNIyXNinNfF/8FRrBUFVLcvlTYQo/pvnwtg8u4Ri
MEHLwZtlzLQPM4waQS3841qpAQCNfppdB2pPO9XD5f8IP0cEn4cHLh04QdupqkQbu+8pDdqT3SR4
d2Yx4zGf1yVkH6XKP7Tqhko0eeaVma1rT1M3cte4p/EIbC9j9yAdOvJfGsCTvNP85EUa94OMj5+M
pPg6TY2grAipiQ67GqvO88GiqeUCP1mSUlbpZdGhfeI1yiu+ksTBPls+GWKzLmP0kqNarAz+O3x8
4h4/g1ze3uIwvKn0OPirr3W+Djyj8sNbenZ/CVAI9Pt7UVFBzW1zuOFOHWaqi/3K1g8wjQga6CCP
Yz5417Vc7AWdTyiFzby30mqtiFF9JtZr/9hat15CDg/gecJ/zxu3GUj+ZbcfcQPT8awXXZlmTtPN
oRj+PnkuudYYCRAbjG0/0JzUITgcVtf01NmkbG3tjYIq8lhWwqF7JtmPzkp/TLGjA6C/60flgWVb
a8stLb2jRMG8nYIDjZ47WE7M5wruYiymK4vHzaWuRIxcJYvFvKlJc9RL2tbEjdc2DEb9gNQ1QXcm
1P2kviD8qy60gu2R2xLNmLEOIiOKLM87O14YLoMp4piBkyaFgsH4xPPe1B52Jeg0gpH+DAxnePXa
bJil18hmWWs8+HnJcBbMlAU/CzSV/h+MCCuKJn4ciVKrchJv4jQ8nnLmIAcUYntW3WWgxSGkyNxF
Lfo8DChUgyiG3UDrsHEg8xHNsgVSnE/bnHzS9yZE9e/GFAsUuODPiBm2CwlwIpFJlglFrFl8xTaK
IFQvS8vQThrcRcN2zKdf9JExYudYIemvWPYE3RNVZUNkA7E3AudSsIGwR4RtiFuz4NomSs4UfK+Q
DLB435zVN3IwPvraGEhwfGAu4tAhs3lAPVARJSBYZxnI7nTZq4MHj6+fc9ynRVy+8Y5nrHJhJKze
EzoRQzpKL8u0tZHyrtE8okMH0ySc7vEXM5r3injswjCFL+EJydghqTuKADJ/hB5jChc6BB3XjOvK
0l2nAqAeYmV9RjG6AO6RZNEggT3pdyj51756OlyKQCsKc/FsHdll7GEimkwU4P7/PCaOGYoYxXUv
eeGhKHIouvoL3fQcNu9o9ExkAjgRGfO5fLNGO49K+vAsJQJ1Hrzirvcrt8A/7ZNKKLev77mD7n56
jJQK4JYV82es8pZZq+It5pE7MKo4SUwDkB/zPnmxzjCxsqPoZ+jBBK6oU6rNynuTXvJG56bR6J2P
L8ykTRL/U3m9koNYEeFxzxOQOiBHqk3cJ8Rxs9Na2wA3kSzkGFFPJL5IELUn3BA7QuEtujamk7I8
C2hT12MF1q//mb3Z0JbB4B6uxmkjQjw4Az6qikgm2z1NjO0MmTevGGB35w4UNVNf9mKXyQAaR+Kk
RdyJp3zi6uYOpJUhtVV3zcKlSBk/FA8wg1lH3CFF/FVuAORYhGxOd77vBX60Bkg9Zil9vtvOmMEt
kLQgmedbnLY4aPevRC2dpRwJaDRLh/a5PCehUdizFtPWnAEN0BeBLs4upTr469SFEqUSva9X42Mt
mjKkDRNb+qRIMsmT/SKmCUgPvGZsGUvrBt21DICd732kbhF0RE4sYI03nQI2wClfHM0zBn74s04X
re9DpgeelcNafdHQKIBcS88T+1hO0TnU6l4IAw8Xpdj1+jzV4pzCQIFe1AAksgAGs6xDKQq7qZJk
woSnap742oMOfudNu5XopzlzMD6mY4asX7JpT+o1/i6mCmmZt8eJ+Jx5oCuO8a8o1rzkpENw+Wrf
OaUGITQLWKir7XvE8ij/1BrR7Zv2sCx1HP1wZx8shpcgsjyAGJEv/+e11tblteq24DNEdwYUcHKE
0rywCevpGvzajyqLDgz0RR9in+upkX/m2aXTRy1ZLssNlLaWSPY6IGyl567x/qSGeN5BJz9EdL81
6hy2RntJaojcdJqTQf5b1VABctYRy89CLGZSVnF52hq2bIvFFJYT19KzmYd4k0rUOHBdeC+eKKJU
cddFS2okRydxWkIJ6UlvFidBtw/eURuogsAjrQ3BCc9NTXNoWPCjw85El2jZfvkpiK9sCc0DlPT2
mwD2c1pxn3yfFap+fWznbv7g90eQdiu3HRcom0zmAiOtHHha6Nzm0GBBLyfXxbrLNuMz+rRzUrud
Y1ye4M//iyfkUTqGZFiyxPB/RgugqZFbyCDFJ1MZ8cU65U4BTkFZG+jZpgGWgvOHB4nCLvX7bomg
aFowJaYYFIYKZhV6CMO8bzcVEUjLg5iA+QwfnCl6N/BYXOAGfogJ++YYan2/egzcxeHqXMpOJg94
JDg5gFhxd58oo+EC4e+fE23IlIqR/EmlR3V9LQvCvci7FPln5tVPIdonzVWQKj1lj9ZS3ckG0nV6
DgxN+/ebXCbqbgBVvZ96tgx34bip4NFugHjgCTn3yIxgBwBHtX7jCFHTxT3ytCePUTSZqKr2Y92/
thI2vFQZQebxR737OdTIlO6lvDqGYuzvelZQAro+cOu65BFLzJbA+Fqlt52gYmD6uh3EMc0fv0TG
TkXfSGnRxGac5EVuADJphdq5VmrC+FVZPOLwu7gvrdw9YkzaBN2kOrkieIcYOIUVtuEQVy22d8hb
PnHSJi294+6g4e86270joi6eGHs/G/iYuqNp2XzEw302pqy3tR5LaOjqmQLIs8oEcgJEhR1EZDiu
FjYh3Tzl6Es6oWt28im7J1uF4qDDQawO2ZjVizoMkYes17qQMXkQdNuGkXVI9tdMvIom1G2t71t0
Ybu58I10DHSo1j/ftutfJWzkWcqBcaYgLhUkI8XO7snBJy20qPiMli9YwyNDbvA/jIZVjwjgX3OL
wxnOTHKu22SLd2ql1YdAnEn9N0zfn0oZkbf+28XQ4H3fmK0ltth1oF/8KbgQl/xCH+e/fZ5ixjOm
EMYbIygFcHeqAwYx09llp0NiXl7nDxugKmS7eDmCkreWvVOOrJ/TZOf2PMLf4H5hwq9yYGJQ8BO8
+QMYyuZEpqi+qrFrDLsTkqzQVHOwwn7rO2UWyGd3KOgmejiKcPzkOe2xN4o1SxKmezEjJLm+VSTe
0J3APlnGZiPs9BS7kqTVat2iX+JmbOXWXufCE3MWjkNnS3tW0JctCeqSjw/6zP7yPjA1L3w6OtiX
o/8OZfusfNX1/JhzILbPuDDJSOMbblHxQ0tmMTUbGODDIEK9yNX0DLZsvLo0ZHa2UxpvBu3GWOtL
MplIZrtqni51whDuk54Xf24b/7nLA8Q1Lq7ennt7ZFHg1WN+qBqNpQNu1Dl+sGNirICe+TIM0qSI
+Ylsx4daKX02w2l/mkQipoEYVE3c68JAxAAnrBos/Sur4omexkgqs+aSyZnu87iC04R//Rjo/zrR
yo5m/9I2YP5J3+pjJZXDlnn+P4U8SNIqpE+KVs/x30gQGIvQRNQnMkgOXtPBf35DElm3a4X8rcz2
b0B8adTRNtSGyJ9SQ1aQInzPFvp+OCP+jw62E02s4PPKRFirU9uUcL8H8tLjdv5a3g23m3sLHHZn
Fn9DbH8UJDrMj19NUaSq2NRLgdTwaU3O7RjeK3f6VNMxh/n77bKcBq4n0UmrortPpbLLNBasjjVz
0I614LR5/P0eHbjWrNfIHNUTkmEdGATw18GMcASLVGEy6qJ9Vpuhis0a4QFtRBHjStNEsWt6gmyL
/8LiI8JqcWS4HGNiybisCt35cwhIsJDP05a3fJOZivlAcUZznBliym4lWZdQZ9epz1q/2UZRNgwF
5Ec4htbLY1dbfizOXgi1wt/Grru7K2S1NQzlaQ8l45fyQJ6WE5Eh/VRgp4sx+fnL4fjOTSXrxX9G
24E2zyUkOYGc+Y7HYLMJvKeWU1nr54YqfaqUe8B1uA1E8M4rx6OBnySc2ckWpVLyIr2E39Ge0cAN
jswi6kmPGd0QOFGy+VXQSjy/1b4TGmSGhCTkT7GI9l5tryF5ZdS4fx9tQkTDl14hqYKekCUKd6sX
1BtAsSwdwAhb8jxq8g8Zh8CD9SoydM2DP1UPrQefBp3RQYDLQBh5gjtvXR4kgFNZQRjO3FHMBPro
E8jkAO2BKitkt8qMdQPRiByobjvlXcdAcbG36Iw5dCum2tOcz/2nmfp6uT6KOVefVBKuSgo/6llP
CjqhfJykxcNzgtgWRLBqYrQJX/MgToU/52mG8G2Q8hVHNkXBVK55fnofRUKeoOxLPa7ssiyjuq9+
giTMMJEnuoXD0cErDIG22tm6wcyjgTIq6oOLnB+RjgQVqHf0SSPygVqLrovm3h34v66rvP4laj/Y
29F464TKfH5UN77VwPFZcPUA4TzwAqFsL5yHOsIoX1KkOBxLV3IpwOr8WDuwaKN50vX+qOMJA4r8
MESodbd0A6cRL8o+Cwl4MlXrIvMMTHR1w0mdpYMVeuv5JIUTpGwzGJbORS5ncwRm5h8Rf15W0Q55
SJmPQPhb6Nz8Y58Stvd0XFa/TT1wyohqy/B1zJTY+GE/O543hNcpu+PSQsysg3YfnLzYZMgkadQv
3t2CvEweUHgaHz/DAoXB0HbGhRvwqFBiXPSCCJr0+y1S/LxztKK22nxFHJReyxAyHxGxN/ihwXez
6H+pp7zzwIo5mARbjCPZooBpEfOiBaeL4Dhc45eNGMKu3pczT3VCtuhbedwT9K3OfAi78QQumqIT
GrX7wRuw273MlsPiMP0x+cYueM1N3MnrrPRSk5cBpE4u5SjNGJliFjmymMmgfH+cMfMYzG88zb3N
e+LtfSTlsgvEBSWx0wMSYLgeMEebvI8Q5cTRQFUOJcQOhx8Qzr1TOowSwyjjsFDJ+1w7iJoXH1Sm
T+TKKyKc762DLZRPAGJZ/0QqTN87ZdUPRby++deK4AtS0lJkGcQ5H0Yqhfpq4e0YmpHnmqEAX5Pz
N5Gip3igSQd6IkUzDDeFrgwIcDC+yQ+PqShXlwFz4IlCW9ehHUsPLNLd9b7MQ3V/GoMNOj8aBeyq
FBJb83wWVHVtoke6Ye1ox1MEsREJkXToPA8H5IhtYO5ZNwE4X15WTHRxfVVQS0ernniQM8orWzvg
9C7Qn3j1gbQkL+oW4INZZJOuxtemjifn/4aj3fu0wmqlbE63TTzH9QOVvullMgltWYN8UfUNDH3c
1kyO2TmsGrBLt4Zoljv6OWhzvTfo9W0d8ntLI+c4TPA4vWoH4fZKUQOoUqrxYDthkU/s6etX7i5D
ign8S9EG3X+zaSglcN/6FHqm7tn4b585ZW2C9AOvTAmW+CHAwb2OppFqcSZce40lGFlp5ckTxfJV
DawGjT9U4zHOPPn8ixcWIVk18H85lLUKfK9I7miZbe0x+SugI1E5Sjt04p0iuQE1CqnwV1KwMlhH
DAA/M8ftZqznUtVuQAw7hL7Rn5ckBoyrhabAbXmwkSyF0td3pU4GHL/Gn/UspM1eEC2YrzH946vk
ji8yZzTl4QSPefZToQCWSV6ZCnm3AE+eOMBkVmYDXiE0ZO2+jjdLZ0kW1r01/o9I42pSrwEVzsYL
sFaJuDFB1Uf8CixGKSrKmYGNrYhUaFy7JiWurDgqFHCiTKbCdCNnAWUlfD6RJLgN5BuCP9BSTA6o
9vPjdgn5J9LrvrehvkCWckB7P48Y9eIZuKZkc/pyvyWUUkRoWyyAh7aTov1kVUIh3XXv+PhUWDCe
qwUwcEivTV/l6UOqVII7pMtr1KdsQbueo29oYq1Um1o/+3rC0emnAyE/POCYH5/TrR8Xf9JzfW1g
OObIHk0kNOWBGPyMi4JbPNKQ7e5N1BagOw+GlcDJ8SC+C4pCtDGqKJAURNE+ZwLdgI/FWu3sO7Qv
yJOz+KYzxIUz7EX1Q/I01U9Y54dLXvrEnVaT9TwcRVO1T1jZQvZGe74fcwKAD2daOmY5/Z9kjRFN
xBGCPTfS4ntkqoMFEnFbtR86OWGXHoF/GAA7waIV2fD0CRDjEztPa+sCQrE8OzRNPDMsTG5RsmHL
DkZtNbWwbUWRsO9UD83b1fXUPNaDzWBKjRJuFtPCx/LKjxWq95ACbAowaEiqf5h44uRAoIMQlGwc
0drxy7hvq9syHOwgOyRe1Ygl++euGUj9QCeIdGcp9ZJntjdAHQ1Uth7hY4w6ZyVjPoelhizLNg3s
owQ2UGpOQAIZEKOKuqdkonFiFt2ZGXKFqVuPaH/LytbH2/+N6hEyGZJpKHF4aUMz1WDZBzU+mThb
iWtST4gOzUuubvjJNHI5hZW2Lezbh7QRgqwhLfo5jhZ6z62FABdK4XzF90rZ0mYTBV4Q4UlauvG8
0grl7pwMphfaZ81qTus28nMpf/wH8lUKyn8/6c/0yXjLC8cx+qU66HowRsdGbCGJnQo8iMyXlFEw
NO3ZNa8T/HyBfO2pKFZHJyDs8oSBXkvIbnPZ8Te2Ki4Mej/ytJym4toaC8Aq778Gc2h8MLoTgi5G
7svrqmhKykL25xSspX6BAjT0yErojRWmH8szwV8tUIMoenLxHfvCtqH1QnFfcpp+nBLmdqLU9B/Q
UizOmRmRhliou58ErVCgNTDSU9e+HlDVEA1vSLsBoVzuNf9q097vQHNwH3IrVqNgwq0LozTDEZUO
gIKQTpT/SAUNyuji7af/xcyz6ugIF4+0MT+WfyRXtMa6HsNjYERJ1q5raI7XbDst6V3yN8jb2a1U
L5W/thnAA/7SqC8wfpmrf+FSdWWLsyfNztI8IPZJMJ2+a1zi+A4No1uoXfjpVEmaSC+UFflDHb2d
3FK9rcIhuBRJfxUr39TNp/8yXKdw3KIRZxxyYIjucpTz00YZkjoEBgZm5tW5v/GZP6s05QEiUc6m
OouUTzotDFzMAfhXhpRDTZ9sjIGpc8U7XzrcoEq+aET98NUI49LeLvrB0MYa2R6wAZiplP1vWz4U
LYrib54ZQ2ChnX5p9+JJ/KTXk20Y/bBYEnBqvObe+qCa3PKqanum2yKbcmhXdk4e4g6m2/RfuPAE
hTriIzUtvy/+xY1VKGeeRrZtEjep778ADbKWlEL+Q+eEUFwz4mS0/phG7l08BxOOHMaiDxCtrdTy
TAhpO3kRSat8ktPWxDYr9arMLfdiSBRQbTXQt3Q6l5ICXXBR78k8cfpAbOLaGDql6UMJR80W7Xfk
aBXvRVthDxgEgq5syvjAXWP/gVzPk6HyJvKrCQjRiUxSWdtMRlOAtT0VE86UYD7mTvhkttkgxIAm
aMyDErur/6f+D/OgcIP9pySnxW0LmLO04GjnHxAPAiYd9X5xR0aeQNr1eRqgQpv45o7DRETuFuRh
C0XU29YPdYijZjjYd1BzTw5mRN80ukVqpKSzNJmVFNHbbevIMNKX9bbKonKD5KU6A+H6GLbcWROF
ZoM7cCoIuf7f7iGv7VhnzmHlPbgZAS8ZBv2vjt2UJ1WHlhVrUyshORs9hVX89k3DrsP5JraCd2Za
+hKEm9zpMaSkD07NPigrxSuqujP3NEtsw18ti69xjmk9n/lOdrrNPziBpqSonlLaeAbRhWYiKEE1
u7DHfsafqfGv5QH150Zmq4r87QQ18OSZCQWMvcrBMtbftXfnWfbF8xbIiA2n6DRr+7R00MyfO6dn
VgqwGY50wRfW2LA3etPl/NTCrr7ZnC6/C5PMWOPLgXDR/ctzfLlyaUkinyntw8bC7vgDnx7knubK
tqxDIR1X3FrrOGEN69kWbfGFyRGQ8xM/6iUwXBJuDajCWVJIgJIF/2ZCHyN9sfBVtu/k3f8UH5C5
sceRCG8sEkeL+cq/E3gKlSIi2MY13TTbqPc4+CAak3R+qCH7EVR3UMsRD63sjx4yRAPxU56UA+Yf
ihJCYwBtreYpjmQT8yfAmaGsvMWjPTQNnZHH2+yNbNbMm1sgFtWtOJMkIpGhoYb677JIZtrE2xzg
Bf/Z1w0Ux8txpzrcmIpZZWad7f6BJ0T5aUKTC6k+Bp7kIbwpHy6RyPg/9+3hgm5ohWG/7mo4u4nt
g607sRLu/nv1Jte4eAKsGZ0p/zmPyVor8JDhnGQkYAnEnA7bLwHfrESBiA8aOOaBRAt5qaB0yXkK
ch3xutcXZnjQxOpnJ9YeLQeBOvb9VMc0AmTqdzZTUyyPlKpE1wsj7svY0rnHtYZssCTMh3VPhn5W
QJ3cq8/Uhr/9AO9q7pD8W4ddrRpre7lPf/qqwW9ystX/0huNkuaZG02xgrkmLA5wDc+Jhl7AQBHJ
o23I0mvyspUWnKApRhvcccMxl5xGRdfd+vSAWoz8OjDIsXREDtDJJVYUlEPBjHwQIH5Ct+K95Zdw
v7nvF07+YfAr9UzgovfXJn3+Y1Obc77FJMWlfTxIsEsfN29v6nY/Mx1g9hRmacOxxO1U6pOADZ3c
H3SjpjnZ6CN9Awuj9V1l4PSJ1+Sagaxa00mOYdh8GgcRrb5X8eEbwWC+61om3wfXbJRgxNXWmphd
rByCtxZj/boYdYj7I69FK4E5169Jzp2wKGk1s8QKeV0grzW8txYro/qhrHvsUzNOOAFxanM0gbC/
BUZMOIApbbt2Yw7K8dsdswRoR19r7yon3z+n0t8tOIQRrTExDYBkSx0J1bZHFBXrgynvx0ZUoKwJ
684zxezru+3Rz/w4BT+2akLc4rDxJfHDPZz0rcoywIyIHpVpRimvEJJSurtk5nphmfMNKR3+PF1Q
qzs6FKTnDZdpDtzBouUJIYILh9boi+Xu5/7DXxM1A/3BpHLEp7CRw590TBjPRU2zDt/jw/SzEgjp
8yhppDZXO6Bq8LcZRwwnXguYzZqWPK+deO4yKUkMD8Nx8cba3M23xdiBPmcoi74gzLch4XFo5X3S
d7YALmyyzlq/323EQCrOew4aT/nboT46Oo890p880AHBuex4UYhJ9kkrmDD9wINm/LmXPduoww4p
30cUNJV5iERqRXwfknJdyOj+fV1yVrc2pQ15XHsF4bUL0Jslpd2awaurS2MaAqkIODpjW1xo4SKT
KGg0PbZlxicMAWqOrMEokizGMwks5GXaNS1A54mBTxfG/rFFvkbquf9WpUSmHrsqxwBzTEdZO/xW
DRVJvvIi+JOYSOlm/DM7gz5x3NmAQemcIh/PUe4tF/YQlgcck+aD01PkLPMyJsQQqFgEE1BLcgFu
aSf50w7K0tv3X480fTVAA1YRvg4oz32SWK3yfTqBUQ5M0BAz9lb6kAuWVXHD5Ymd1bIWHWZk2VqU
AROHZQajvVK/PKZVpD81wvij8KW/E/c+9/0aws+Ys2UF+BdFfycKUWRRTIa2whBd0JXF/cXMQlmJ
oWT5/xoastuv1cUBDUIQ0oEVozSt7ZxT0G+GzkmDxt8Wdvk8zZw1NABhHSIEdUcssMOOyCl50q4F
L6U6otBQpaigaexyGKZhl2WKZQ5nqmTY+5I/32wywKwjXAM/2O2BeN3uaAbWDIvfhhcfJsMu/Vmt
GgRQPhjINtXTK01gbwVfvVMewqTBV2Qp5Rors5iGkuEY4alKx0m6rPZXhBfyszq4EJKVC/rXDe0b
cKyMjF0Ig4DcjNH4+lQVPNzzGiFBAVNNkEb0LWg6+cTJfECNuxfUXg/3+pq17IV+sqXnd5Ze47vZ
QXWoP4J8w4wTOSZto845dhe6WZrEbhUU/Lamak+KI09tppUdIFCsUIHIAuXS2g4R6WJ9rrl1y3WL
CBJuVlZ/HqDcg2RfsOOTIVk1ClYWZgfzcwp37GM3XChcfcoqOiGNwMLXoJjkKNNEpsgx6DfLv9cj
8H1KB6YVD2bhJA2AW0rErIRbNQlotBechL7/uOC9QSXIc4lG0bxBa9k/gYPPipJlChjH99HRV5fW
D33Kc27NZoGD2HghgKnnP+A5UjXYzs2pz3m0xTWwL3VDoFf4g3UgJxj0P2M7luBJhHdnDYzGTV17
b8PC3pvyyokqMnAERnBBlwRVvfb54gCn08jTOySqCp7NpuLZvpbJ6j8Q+VcZCd/Xg4D0m+sdlkWD
A2RYU59092frma0YNp+s426E0NFysLEw+WmG4yoB9p2WFLYIHdHZWF1ZfhvvJ8NQiUaQ7RqllwhE
he05bujkY+wjqVbrF5iqSoHpRJAv1MDa1dQPYs19Q1qU3LPtmew8zNHy9RWaeuhybqYvbe3N0rbn
Y0UhI1U3dtjdrsrPwt41/mucamSc7ldR8JijQ5AwRP8KtCG1tGvTTogp5VA7QNuft7Yo5P1KwoRs
O1j774SUwH+uwQrdee5cG8BPirhPScnJQ7UNXXrpwnEWZ4XBnFY26cj67YpgpQs8psSKjV6T1pyH
a/YwC5ejUiKkpcgGe0ASQgJI60Gf1lBBkMxH4VdV8WSAmfiCias2nGRlN8cIoMQ6PpOXxlVwpKlK
p2wY1VcymAneewfyaFZF4/hK83QMv823uLjy/GoQMBk6MN/oD6msSWg675eMWPL9KmSiMUhPp1VC
vRM9QQCBdgUwifwFqr3r2rmnIGtfY4EoP6dpuCv28/pZj7qM9RfbzPDKhGB1DakQXeeFYNk7mYrP
oe7XGuEgHP/7OLp7K2gtwkCi0tWmrPRX5WykCYeXXK4YPTVwNLjvMe+VdXYoO4WvTgHCfnjhPqUF
pRvA8aMQAzjclvC3DTJxnpMQRZhB/oNSQ0+XEJxYN6eDtHKaqN0n+NTtIGKGrGNffB0ReVj3Nfl5
WwBGuW1d8zwCrHf/8trEpkhPdel+Z9PdZTH5bauGrFJbQyNBmOBdn+DkjO75krad30QqVp4t/8a+
jz3BF764o6SE0x7b4XlLvNI0X3erBvAdwS+qDK76DkFSyxNfiwTAcHB1lQBtAMRxwWusujAHxtz6
ExR3LodGlf9ucx59z7VlxmFJEHdyJopY2pk9Kn/6ri0dBAfFIDVYqrkguboJEkGgGvGuXZAV61QT
DJWS4J3StKUF8vERJpLoM0MhUlr4owK7ohIxidO2NPchx0aebOu7X11i2GtjsUISssAB9YN0wFpb
H+lWr+IP+vRZ8iKCfiHLvpUy9VcRH5QuZhTvTduPN5XPUD+8Ufk/n9JGBvaJRWWYFbcLCXj5ONad
q9I5jRmpMW0HeDq7S2vEUBIVlp9/afmQrVTQcjxO+/urnPjEc7ebNZC5UEVRRd2it12D989S9VwD
2G2cazSPCNphUVESXARNQxDlyTwPzMtq8QQo5XJGSb7hbuCfTUXEAbcpisP964D857wrSWRQIJtk
UsIJGltvSoq7QHkFf3ntiLhW7I9nPAmDbtAzssexk+DPCF6/JQaIkaX0U+q8yI9bvt1jlSAprttD
Gq3j2rgFOYdrxYYaC6Wyrvpkq9k6VhiZKyJqcMLclgXpof9vwPYYzmVCeEMZjaDYXQR9nqF0TvkX
nal6UurhvaRE8TQYEO3WJvO9OrLiJfi/OtQw8LWj+pxgO0YJwgQpJ31HgT4TAbabcCUew7pv/L3x
jX6RSBDcOMPVqqtPJf5m6iQpt44/xDua4GkDWzMMv03Ec8I6Vst5/hax3kam3CvU+iNzKh1Nglbb
p4U3LInOSJvU37J72MMeC681d9ByqnMVZKKH00xaRw5pMAl/C5uS5ewzLL0o/XyDdzTrxJ8FD7Qo
/wfPerNoGUj1NxRfMTgjFSdPuSEyOeyEYk6hTy482zodPq7U46jN739uUTGMSnMzQxBR7NXp34fz
rCDbXFMe+eQhOkeL7AjwmysRo1pKuGQAIALTRZk973rPW/s6NKrKRinqJE3UgBtqM+w6g4zBOT/j
2aLvR28gQPmnuUp0sjDEmeFs9e0INiccn361lpL27EinmOGRv+JsPgZ8kMI0zoD6x1hxYquOCfse
fpVt/xUYxUk5FtxJOcRSFrjjtc6fX3vsbwzXf2SC43BFSi2/DZ4pMSC8Va1BQOB4+dHGBiCdGi3w
9LctPONBDtCr1yvcIVjvDTRUFPJBQYRKLVQjLgjc1QZ9i6d7a6Pp4gJlxHkOOn8O3VrevZfzrHJf
NLIg87F/FPUQEzlS78ioAWXTAcmtyC3k63k9JPXRFy4ESGFIk4RoNlTV6ePRm/R+XGV7fbgWRnbo
p9GpZzb2nqLOi5lj5F506LKnSiDxV/rAYM8W0f2A60inWWKTSntJJZWbjUyZKeO9mWrQ8XhEngqu
G1AHLuLJ8WzQ7o5YYZxxZ261cVtmPZSXizwA9eRVCTLDx/B7QiQuUijcDwPWHOVIsFr6aJVBABH0
skS3ej89Lc02kaXz+PDoyBOuxY9FwWhDX4bhudOrddfkjkFAexryIdD4se/F0Wc0c23R+ZuImA0b
6o+nBzZyVIllklaGsOODO05LBNpNwzwu875rrbnJo3QrMc3IMxSpKZpuzl7xWBnCHXmtItEI8Jom
wOBMu0hyly13ZFNTkC2reEF2hXTRqrLIkRTrKewk5C0cWFO8SlIc+95Hc2gKCq6YtVGuGuLEBsyK
nCmK/Gsd40vuu9eWDCn4du5c85he95jWZqEjml+V0Ux4VEoft3OJcEw3kxyAx4Cs518Zx4MeHDtP
//ew2FWrUqkxmqxFndRLNzKpVFA43pSA7ICuvvuBC7OaXU74ND2tyQ7eb1Vjq4DuFHiZcRUETxWQ
FBCGDVsAA9N6BS8tR2JzE6VVYm3ixz0PwG9B+iztRPpI3HIkKofGGqB6AQYXFeFpWW3Lwx56uWMc
+qy+1GelmtHxA/kSObVw+01fFGKQzSB8RuWmzQZAz6Y+bKQu7WDxsDMNezRs2DkJxSi6X8uIofRi
4yDNjvbYK5/uhuo3GPtocRkzJEpoadpizecypKA7bklsx/8kg+BpxRWehxmI1xFfnPL46t+fNUo5
3QBt/ELSZUsiy7sR0S7uXdcszk7mNxJoe5yf39BEMZYldJz46ib3AEVpVP25PkeeMsDt21G5e07Y
xgfhWEurGKuZMY8j/NcxlwxPZx82jE6JaT+XFaeEQ8j/GROs9N8ejjTs6UekaCU2q52wgLLuii4n
7YHUpZrvSmebwXQ9YLRZ3aQR1piaEGiShQVkCSgUAI/OweAdERWgKoCXiu98HsY2ffdTiXMnRMfl
LT51HuX/29FQa7a54Pdef9hrfP9nyi4PAhiu2YjoApKsk/1a1Ky2J/oC/p7CuTMG42LGgKS8zXsm
hu3WhpIcuBRIH+52JyfE58MhnqRVZg1PERHp39DybEc8WBjIkT4O/+hBscDNL6R9bjB521WSyU1f
V3TjCAqEFWaGdDzb1kFjnj8r7sXEPdtvRKuaTetlWP9BVyLNWf2jiCUaZp0dQq8JpSMxOJueT+B4
0vs2DTtYuhuEyw/RwROxjjRC7FBqAqcvklzlZeS7JMa3UjRG7pBj0IWspQaQLD3n2kofqLTCajUb
Ohdx7DuszipgMk0Q6hMMFuF88weMcpD8VuW6dGqbwTQtLHhgYFnrzWUuHJ7jfi5OhNluMHDvy9Kd
HDzFHsWT08NlHcDGh2t+tUPEq0agvLUkhgimr5MQS+xsvFHKTLL3aID3cpnqRvUs5CKA3R1b0ToJ
ETrRhG/D52sfLM4i4YIXBP558+PG1YtqepSeAcr8JGQMn1fC4bp/fVmi2lPyDHDWvjEl1a7HF56Z
W2P3HxlYhHCncmDc5Xhz3behf6EEnHR6m6h0lMKhTxCc0Ds2T/L5Y1vZdrkebM4A/06rfLXt2Ixy
v6frcoNkmeU+ksJ+kxz3il/5eREpo9B/bDS47aT2HjpppSbnqollcqEUR0PxBCAUY7pwbgmbk11i
X5FNRHnjf4ObjMcVm7EKr/H62rmwFU3n0y6wol7M6Tv904cQMhJ9AwTpO9u19VQeIZFFbuyJsHax
doEFZ489cvVfWXumLdUEPzV4VXNhc3OmfRQzBiX22J08oO54jwxHa/Qz2e6JFviDlqAD9ItvdWdU
S6DWTAFAFXEaVtXIUJIRMMSXB4fJMr3OgjIaD+A2EQneoYoVHBLBkKjvwE0v4TiE+CJOxLtc0fYs
rbfp1Ad+M0KE90FH/xBqxdFULHJ8RKMw1fumFeFckPhZK8eL8pWsM5uzwXhS25vmBwd37qkS1+SJ
7NfCWzj60rxhn2sQ5/wKvCqAl14NP6+yG5QvPclkyIov8VT2S9v+eAcIuwkjKqcbQK/NS798GEAd
hIii/en6GXk6Aot7R22qBeCv0gb+rA/pWs/Wb7VehS6+EH9mX+d7dqgj++OXxvkfp9uIhy5t58Vg
FTgjB3YNqTOhkx1bv5KxPlscM95oZK6GDRBt7uZOTNOB1R0ygeqPo05WECJJovAajv/QhkTxa2Gi
XOZGCB3X0+0460j+YY+0Nz3fhC3wLSEQ9EeBpww+qF6bXYLDZjdlcJr/YhcpC/3teFerSGo5SXSU
LzvQgGsUVZgZ1XeyS4E5gpnfsQrBUajhGjWEifapXnfBCG6muKpchwaEGmy02eoEBJKvDt0Z4Wk+
9xPNoxh63vd1aj2KOUUu7RYfEkoOK8mp2Khmn1xXeGu70gHUVW8OFpUN5dP+y29mFTpJs7GIGbyZ
KE2+23ufG+GHkQd1NGJutid0Yf1cjJ5uSQ4III3AfnCDuWM56OBxCX7vps+19CLHXH3f8RGm8wjU
wiXvL4+Q5Qb8PZNyj3X7Te9tbkB79PJ5wx6NK58rOkseF5Bjho3urOWpLzTID9o2t5xbHkmVCZXu
1T9fBtlQUg54TMTnOgG5foCc/jzE8AIkGYo0DVM0XKM1lb5mX9nhiz5zdo7zJWvKKPQEO4Ix7xIe
NDP0V1Xqrs8JsxGtBb8ejv52kqoMFaYcpaf9xysBYVhMY/ByK0+tp6UfzK9OCL+TDJSl3j6O9a8x
BD3bUEauysWwxwit62azh5PHqbIANm7KjYf0pUzHzIVIF6PLPeG5rA1ggE8lg+cJiM6nul8jxE+j
fb20GvIt6KJStOg4E3ERWCRqhOOqcnt2TuuNhePKI3dvOlvmd3pGAWUyZ7CGx573DjHfz0qy9AjJ
nj77iNIGfT9kVVTZs5/7nYjQZ4xaBCOkWS4mtYbMV5/oDU/5H7FXT0W4BDHopQYQAt2Z+M5i1ivy
H/fTBT2Efn6Pk2rAB9YK0294t3oGiqdYxw6gHyUHYHEEVbIIyEwQh1P6Zfd5+rwUmzJG0DI6kaXz
AFribRFV2Hbg1YVgINSFJt3/DwlrYhdz1mIxtHlfixFLXNeIfSRYVGYov+9nmWnfyWsaUT4Byzp4
Vki3/fbQRflj7MB42WdGKpsKDud201kJxPyS/qZ96evoG8c4eaP/nFSRUme5+8GgGEM3RFGah93j
+Xr3LZgCecsSJ5ikezIofgJ20pMSsgvgaAXIovLRbQ9e38TZahmqPa2GygNuV6DwGbItMgeqmt+Q
F0g9oHa04Tp8j2zJ1cNnyZHLbXwccvfTFrmtKZ6f/RNEei/RYLoMYpa/YADz8LJvGC7+Oj9sntfr
jfj7qeokZcF3bT8vUHby2cuO6RrHYocK1Rl7idDxiD/0OtJSe2BvHVQIZblyCGoy1tDB1vDkrUDQ
uVOrTWAzVruoaoBKImgD8YH2ttRA2okuv/2qxRXH9HrcTfy4ndN3BhvhDQScfLZQ3qBHeYKKPvWD
WKHmeCw78kySzf38jm3DleSmppomJN5omYcNURVM1Pes+En6XaXAjVt7HLy2dwNV/mIcp11bmqoF
OaEZ78EV3VyznYF6THwme68J4bM+920c8xKAPgap86u3eDP0jIm37GU+iJSX2bSxhcE1L35vb3Du
zrZRtx3pceTNKJ+yfya5aO8Y55IXPI7UuP3DfzR6mgFXLc9FHJGLWlbEnLKUNOMYw+6P2Q66yh/L
Zo07kVdGCyJ0eDGo/HTKAe6uzwtvgRSV98827OyfaLg6fWF/ZaclkF3X+LNQBJsE2ZD8OF1b7AGy
MfZ1yxm/Kzdpjzg605kdfPAv7UKtHNMrOhhW5qBqQwfidMsbmftRUqzT8B4h4zb8gPgEl7EhWp/Z
pNAyqjUtuPmj3aZmEBAk/uNIpQ4zUR7vxNAmRMWHmaO2Ovcri74uB/U6OXAPrx9NhHg+6yYFWNO0
AKt5jlzejWmzujXKuyP9V4od69T4N2xIy8RyuoRWsf/fvPWO77PJ3ZSqDIowieAFfC3yMaza5ki5
NxfUU7sqKS0Sy9+Ze7ga7ZHEd+k6HNjSIkkAnQT9W0oE5Nuh526kDFvBpClnekO7OdRXfAsEUNww
1mm3BnmzAenhDS/JpZ2Q2rRfO3IKSRB91hwPs/WGZq7RBZ3kLf/bFWGoT5lLUheH2B1cfAvEn/S7
JPt6JcVv40QaRuqEByvJAe+zCs/BHfSCaoKXH4N+otBnhVExmYTiLmtuMAI+ifwC1upJb6sxByiN
o919yDhIBqWqCcx8ZX8AkrsNDas3flDZ8lGrYV7jvEByMixBEblfEyibhNCobRgNErkDgPwN/Qe6
RFE6ZsFj6qCwCWlYbi/RA5RcLQSaQ4oTNpa0smDOCRand3359KrEVmVsZiyR1jMDmsVm1PucXaa+
3y4grrqMC91AWp/Vd6ZnteWqkzaexCBWGTSQfzeVI8oqMfDBPGUEGW6QROrnCUU6T+Db4TLIugEP
HIMbX5KaXQoKwxdhxpugMPdE/k58QF0DmcMP06wdskmpylcRYxXHmJ8MB9O0PObRy2PVGuEa/UA/
EEUaK6k7fVgya9eRjAixZeMsxHg2FSM0DVxEdAXU9WQyACXtGnOS394BjGfezEKdrBGXDATxDYOE
3gRYgHI1jHO8o+4IrdBKKbQ2XEJmRabt+xByaqQow7gH0+BSjT8oT2f6SCClODXZdq7Dj/zmNFhE
uD/543Nf4Nvn3QrD/4od+Gfcf9VDrLJdJkXUVRrp3Z/Fx3yAhpGEDn+7xRoz6BFlgjeS9rvpTUKN
KRq3UqtkXou5dNsxMIg8saYFBzR+Vjg2f8NMR7ESfl+dDA7ZntTHP5Kad3tPEyWq9iVf4ptkOWxX
QgfnteB8ajZol7zYRDjaWaDBTiUBIlbDx7tQbtp4oCqbZt9Uq25+O1fWhzhFCAH0Ke/sM1qMYoSY
Y8KEsyDl5drjNi5BbHFjFQ46YW894Uu7ebdrWjrYMPx7y3h7/Fop9HsRqa0261AWgLfI2fdgmG7q
xeHx1a8xtxnS1sck0byDXGpWXm4gUwpJd524sQwzOy37CcDDUcA9d8qB+ysTqIQTrb/wVmu9IpTn
VwSxvwYCSzwAMk2V5Ue5jlsgaIp4GqCTt9dhDeyvzBAhriZXg2BdJOEI3Ts8BQm5nk/hNezIejNU
CkaPmc7tAOHyLR3Pp7M/SNZpHgBI9Ufv/wwP1NExIV07MN5+oZch/rzPlcQwPnQEM7AUOranprCw
E86/ASpg6EnO5fzp9Kl8bosUUBN8HzNY4e8XG16BTe9nkaDL9a6h6oewMEKDLW//9BF7sVhhE1GK
8CoY8IQ9z5tBPmwdnb4wWwr8G9AyL5izl8fwdse6yrL28RI0O1JQFOps+fib0pBeVVN63UtfcMyZ
joXAx7pChWCVt/7Wquq5a4ADmu+Ss78LgIrXmhGMsEtZpWy4GdYoW74b3BwX58swvSK6O31WdCc9
xSwA+GHg5gAa19ojFybj2Dak2mIt6iayH0SEqTanE2lj7O7YBPgeVNHTzbC3jRmj+EgP2Rd4c6tm
D+B+gWJrM4xrMjvSaesdHVH508tlCvU06Oh03BnjbAV0kJrzIOInTJzoSF7AQbhIecd19gJVd0ra
8fAFHWjdc+nTktbCTRgxcUSO0E87YOSzgtKiaIRw/Na3Vj7GMi9zmnJp2rbxOlMLtRpbhGCaOhfF
fLYI/rd2F+IX1Py+Agf7cyk6ZNBKmPIGUNqHQT7l3+pdt7EsAz4gY+pfHjvCteewZ5UFMlAQsm42
oPT64TAPbi1equt29LoZ+KV8vkMGFCRam8yh/qmqgiuxbCiNxJZnnbmglWi7cIrzucXzMsVrpxaY
KIkAwmMVSJWfhYQcHRnPTFU+KXgvIE+DVmmhAvqZX4D5U8ZSyCOGEQuYcBuP5NMDC6QGr+6mIcRs
i86uYv7lZJS6lOkt4lSU/GSWoIzdXXhhiP/Ctg5b5Fud43DPfCOBhb58frl+OSxJ6srcEFa9yulq
5mYfP/HbMdFMgPJu5i0RFMO+Idf0X30RwymuOw16sjSTsUsvHWAYlg7fAkKJUOvG4pppIoGQsPjw
Pqr26odNkSsCqUCN6XOkGsGbsfDrCF5qs6VaC81w0w0XjHABrtNuiwhDdF7Z/Cw0BQUI7fEO1snt
VwqnCyOZJbLZouCgIvc7DiDjPgIBD0MPFmVA5xt7J0Bf6L4MKLQDjBSH4uZtVwhKy+KZc5NKZ4ny
l0OKI4DInDE25brnlQ0XIFI9ZDfjIpACjg5gmFxwX5g1bllee7yLKg+v7cV/cHN0CL7wtkax+FuK
UWaTqp4K6HwJs4zMPC6Knijx9mjlAPNjKmQ/+kRRvreYdiEt/+EkDLsIH6MvhLPj1Jvwz/0x5zQX
bLfSaEP0paAGBAFxLuWhiag3yQ54df5bMagLGkrpMky4k8lOgPxbxQsM8lW43GvfI5Pvp5uQDVkA
NJnJgew9AMvjYqtauHB14RPL9L8H0Z6xwfTefd5H65edttcxZhTs4SvVkQCk1+5RNY07bVqxGzzK
TpWdcu3NQDhb83jNoRrj45YcEmU0BTG8KFp20ginwlGqFiw0grtAk2lhyIH/rvxF61oNJQ8lB2mU
JJrqQ/AnkGxTiVFXroofLZ8+BSX+RJoLu2lFZJWpnkYw/BQPsWcA5V6SCct3WGvFwa0cDRochUfi
23lET1OBWn22x9T2MPcUm5GtT/dU2/S9kw832866mIQwyp3SHLjYA6L8ePkaHAUA2dzF2Alovpwu
e1vO29U3r4FrYnuxOASNA/kz6rV4XmqQtdI3xUi+/BtEWLdhcFloZRGTkZbvi7zuYcptaY8l6jhi
F7wmju/szFU7S1NGTMisT9mnjmrqj9JVCwz8hPdW8oYR9MjAIrgtW6bckWOc+lzVjbDqc/COIPFj
7THLvA2sIvcvhYjzeUfmuJzm0qinDizkLDAClWIs1pNlgZkIqpI9kgQDFndk6kPwx9wrkRM07D0l
BVRWA3cB6XUAWNn8Tyg1Or6uUVZVGNKmlYMxl+KYFKxYPUK7rPaale4Qgnrkxl7ISLk+fgxKPaW1
zBVNzEwpnJzIdHhEwv8n8qhj4uoutsHh68pctSyM5OxNiRkpTb1LENUq9l3IFlCd6CyOEWM4f4y7
3/SsUmjHFr4laD9JsCUlvh7XgkI08ALHl7nQCtMX/lt5+M3PHx2gSUYAAY3oy029u4kPXIDr9pzq
BNUAEAcKZS80v38ryC6+t5iSXMtj2fFMt3HrSl//jt+v4Ke+1W2HXeWrMytenyj/4Hyl7Kb11Jy8
DEx5ItZBC4P3962VM2OKc7PVo9AlMtB0SBQb3HZjFj/brxvIv6/lhIW7tvNo5HgpS2hBeLD9MKpb
YuOCTKfnPqzhrH2pVB0W8shJTU6tfgv2qzEXTyIwc5hrgVmheDsmqlmkFGjeW+pI2MMJ3DTRiC7W
3dNj8a+cUmrHlZoSuRoI9VtewBaTpdig8WFvAFQKQgrHXNJA8jVfCpWs2yDFzcyUkJ/tF7ZQX31z
wnpW7dIZU9uIm5gRe6KaPNqHRAd8s7CX9UoB/JMF1Q9n33qMZKPkWQ4/lJkNOqI2UY1xIgi8W+yd
mHvAPmcxJQ64aEwIP/CJhtPBs1aAleysyj3YrI35EeNR2VEcUlYbIDWUEh5anphmZp5CL8Q8f6Cl
AY+ZabSktB4lFG+c3DXd5AwzqH2SWRVoV0a++LYPZCwF6nBwbL8sKV9UBqrK2Ouy6iYSRuPyfDUe
fuSxmVBRK91X0ui1juq352JFZboy1bWUBuVQ2bQlsAGE53tY49nDln4G3Vu3ILs6Jj2GCwuwfSZy
ff1AxNTfF/Mw+CuYk3gVu/mmvnoj05yR8oGuVwTvf8xvH3hRGiZ/zJLxTsPRUvnoktP5QOwVGjqV
X9eqiwRFdKGD4bsjFwVJrnO5hzkNdIx6+urTT6BELsI5lD9YTU6RzpcWqjeByNMJ2FPeF+5sm44z
icvBUZ952touYAw8Ifn2eINSc0/QayC4u1ZLC+FK884MdrQ4Is1vqZEjscFYI9I4mKSzMAiQfJlq
1g3tOi43ze0X8uQn7tQSFiJh92X6xmCIajg2fGe71tRMnH4Cgi49feTINRQnRdvwnhN647ommUtc
2Gr5nmM30HdbLxQs+zrF7zpB7x3yAksIizzkjLnWVpP3iHfyJ4aDCDH7Tq3rnTU5OVWDVAApTUU7
wg3berQzI/qP1koVDk4QNtExM3GTQlErGo2pOv+4drjlm9756tgbTfoqHPemdzk0KzHk8ZA/4RLs
JEQVyRrlPnXMaTRJbD7Rhfa31juncMGoD0PRCoz2RpxooeCS4oiDO7xMnD6aJxwNqr4pfKK3Xsca
O24tem2d2cS4hnHQcu9Fny5W69do24525CDt6KnRCndaJwVD9JkTvLWvx3R0wf3Um9EL9WZDwzLz
w4gKUrziX4sBeCE7V+AvJ304DkniS94TFqWcORin3aTDxj/c8+f6Jo461e35iVVr8iC1GRRTusH3
UpfOQFCAaw6e6rOCTORGaC78hbS5HyHTT38mZb7Z9MAvLzSjAIryXtcURgfPgT0Ac47XdoPpLgs0
nuIdQ7bNUM242PY3vVk5l2veCD7XbDYWudZ04ep5MRKjiznib8oXOYi95KmN48GHYL7O1AZxV7+O
IHXYVzMgq23OTGZveyVfGtUOrV4M4EZfjB08tiBWeigOhN0kdRIFj7zx6O88Gn5NkZLl2hHeN3/X
iNBK31gGsgTnByEdmcWn9wz90vTa9Vuav5gRUvfudq78OBtI8yxKgj88dlPcOoMW4Vq0IR5O7Vh9
fwvWzSD9ovnUJQ2l062t22v6ti0Xvw4KyQeF2EA3xdeW3tStY47B/Hi44CbiVbxEZIWZOQY8rLro
ZWwIswhi2HOkArz1YOTqdaBIXWviiyuSK9Tnl6WTRNluMyn6uXYgmonpBG68BF+opcWnrQ985QsD
k15FvvCKCD8chzqNltckMkxt+G/W7HvXfBnQgWl7xqQtd5eA7mVqpW7ugKhBib3qVUeyjr7oIeMT
TM9yk3ePzAl62C0z+QCS0QNo9fUikVk1m822lkdv/LocEcM9ELzZybHFzMizCd1Q7AraQ2pzPyBz
asdh+SRDXHp6Us1du2pE40FxgQ9rLkR3fxDPiRDk0okYvZzy8pXYOqJI8FosqgthFyuNMzD/HL7G
RgVS1n4tu2sMYK0zN9Q4QK8slUUdfv13nJvKdz6K6ip7+yks55VNkoTyqkrHD78ylF7DNVpwx4Cr
R54vFpNlhHRKlDbplXPBo8Y0BvjDZp3Qx61q6d2T66BAQ3dxWWck8VB4TvOJ0kS3irLL5/a7qXO+
RR3xLCMMZD5Xb4Biz2LOAei5qGO1oDTDQ2fFwTOSimO4UtRkFT0qBrd5M1008USBjlY9RwBx7jNR
rUYuwn0AamGx1dQrwdPvHLLXjxfoedkuReJyb2ARhBmrk7HdKXv8bsoy97vBDj7UHpYn2CtEke/0
L3BsvYN/E5N2CrXlyOpybVlpG2luplEsef+CQSuijc6/JXuh6k3cegbYspbP/c7oFz+GgrVatAPh
Tv5f5oeZF3Hxw6JJxnqrhTTyUmL/x0hQqm0nOdlb5QmqcxV/nUKvgiGnBMwJTFfSenKU/Aqr8MzA
L1IuB1mCbMfwKxFthtu/fsR+tdpuq4q45wqb4hzsVx4dVxc8/ZuadS7hgs3GyypkCrvITxPzXTyY
7p8rxz65b+rbnAQWshltfZN3uCFwmjga+Qri980q8aNdlj1xrEwa4lI4eXW5qEX4hsdz5W6h+H04
5S3IqG5kNyewikWfxdLbDPZfODo1nVE7Uce8gItWBxkO+EeArbFHdeMSFMLUB4H/QfhJURJ7AQUt
hSlVxg4iFCmyPznXRnsYJ3mwgwZ5vJzOSkrbPwo+pVM/9PmEqvQPgEkgMvW0e/xLz2diylu6z7Nk
BJXE+yzKoBnitCEURncFoCFE5URUfq7hS7uQ5atRx46FZTuJwq6SF1a1//KexkIHYrgSmKxmfQDw
zgh0qQgnyLdZdY2JMrUvUH9vyD9NbZvVuuyGxvN5iHz0lUw1z8ujbSraAz18EZeqwGijHiVOGuww
5x01qfLHjUKcRRs+dISXK88LcDoQiXOTU6la+Be8uhihdDv4ZqAjG0qNxisU46ayw4tIR1X56srE
aXMF8IcCkJaVsL0hhdI2dtp414/hghEuZ4u04OFHayG8/esCT5vtuVRRqvYBKYupCXkaQxLLMScI
SKbd7Fxq0RSdjfMI50HyvfJ290e8sqAHMsVTnXYeqAWhwXHNzvKt7caYnBRoIojPSVlO0Z0aIDbF
pNmVLnbIcQbrG18tlHLkn3p2KFg5lCzIg+TvHy2p+4URQIHoOZY8t2i15HcxCBu2TggQgVHTryu2
33Tx/9QXo8MM1Z9qTN8qtuTD/tOVux3u8p3ugj7I8vDozg16ZCRBS5qfKncori5OaE3o0CoSheqL
/6KOlrKBY4FSGTYqMjSEVlFv1jWDboqiD5lwZcf/uY2LO4Z5wS8WhSjCuyfWQXv/uNomr5+gY+CS
Cm/NNABXeGVuOn1FaL9e6KqikiRdDd4ylqfivLUzgH926hP2UWS2tnnBoPmypZ5jagFUBHhdUvbf
gyaF+44eZ3Sk18rCu6Ygf/2xokr1pYNley4IDNyUTW9Ib4uUYFp+vm3vZgFwvFZPAIHZWkB1xmjY
65Q9y4juRDvuEbvedSgJtiiPE/NOIn+lT338ygAluIcnaoJ1Mt9h9BjSz+k3Wg++EvNJQPVxMY/t
Afgr+9fGX1iqZYBsR5Jr84G/af+vWjwacLFoJaIjERC+olIT+C4ldcZraFXWH68qh/8atvTuJtem
ae58GPbetEY08ZqIC/vwr1ZWJ505CVGqFhPIcrQM8ZrliXw+e96Jsm4mgJ90mngtV5ZZMmRc5aeW
YLazGyKWF0EJUgcNZ/394d/OnKYtRGCM2q8yAtIaHs1PoAmCkVrqQ948qdri4Hn1AzE0W1iuw21C
n50NpEP1VuXF0pf81/1DJKdCYMNgDh0cv9zTBIVXQr9KEbbzyn2lbepq3wjNHmhvYObzOx9w0WR5
iE5Nv0Xp1s/oiw5k3HsgG56AJ5LkLxys9Z+h9J3H9SumU7CePFjoaSgqCgWDDEo2J3LcxkGZPzE8
cdM7PK1O5O9qvDHsYBCZIuULZkS07g1jmwj+B4OWhY9L7lTWGhgE2i6l/8I0HWXRB2zoksBq7Fzz
Sj/EA6U+/uMiVpfNMaCNGJQCfnxaVC/wkBpDYkOJVKFwZR9GAhH/+lQ+bgDKmA/nxAORW2TlgpWn
8BrpdQ5igd7SinHKIxvUoFZ+8czy0EwjFvYmn4V6IAmB6Q0fQqTFnN+UwoBny+uyFtoV0FObKEo3
yH2s2NeTaMzHWynNoAHwlTg6NfZaZO7eHRhDQAxVU368dl+uAEAD2LqQAaw7ieeAH4/s4FkXiSH+
FYCCOX+OZTfdFOkVInNwMiBdZ6o57oBHvmyHKC9ebjtJQcsOXjJIs+tMj5XxEWa/JJp3kP+JCjxx
R9Y1KjSzKfbIDKGv9YNaguCC+qoRgAYnxcrnnrk6KRoEdk7GZQOnfJ+qAJvkyzTrzpt+CxWV0eqU
iWTbnONI4H1bSviJCGXPjFEFLbTD0IOUjXJHzayoeoUenn0ge/StcVMkgxcFzkSMzKl928bP4IEB
z4dfowXkRiQOwRqBC2wxPskdaKVqbM5evOHTKG+eHt6wKgcF0dtQkc0hrFlXoUyt5g1Vv20YUMj4
lPdjwWdyhZmPIY5lJcFw4nsTBa3tWhbdpz3kDapuYVXAO/q1z62tugaKaoLFkgP4+zSRhBk+Pav5
pRpspaN9pVum1wd4Nr/GB4cGDjTiOVplBkMtVBk/c3+u7Lskfi3o0gG+XJlBeTir36jc5musRuSf
5fJIIEyf+xnOXSmWuYoL4d9GfD64k0aLxyedR3J4ImrbAudR5Qls2dVMXYOgpx8g5d4xoEI6RSNJ
9xRxyeEq8WpcaF2OiaujdH5CmU0pLEUmAQKUriCU84mt11P409MCEkLqW0hcN+5ztICW3ufwv3v+
xzpEmx+Kqop2V/NQtME9kIeEF5Q5fkHRqn4d03zG8wWFL9/a3Lk3zsQav/fC34Lk6pSGLkq9aXEP
Gq8xtL0+tFGMAzBfkKQ+ar0NlslcSRpxyZ5wTmtPCymnE43GsujYzowJJiyFEQC3D2rqnZVMYZge
tVPOCYdvGZkKbvREq8p2yOIM/nj1PuAiZItOyjWAmnTKo3MLPLUciQhwgTu1EQseTJsON3nG/XQA
ZrouYH8ZKyijtL2+uFzfsawoy+ZIyMkIvBRoeKR35e2xLpmhkwHuJMdlhhG2Ue7rj9d7anOpFXJO
gWTw9Sqc9Ry63MbD51rZtn9VJhxBaKjvPchMCvuVYXDY9E5HRraxCQP3ADRKgWMXiZo2omdsMfVP
LDls6bnB06AEMYmMW6ZWr5UZ4+RjzSPI/xzVBilohd03bSxa+zjFrqC38OZheDNxMKebDVFbyaTp
wzgwniYtm9BU+WGNVXvHVTlKpdHOFLM37lxttuZNreNYZvpEcwBXPBgpfGCAy1JVEco2RbXd4sgz
a6VwC8ZEmqUPEYRrgBfdpFK2E6lqjukp/tW/iBrvJYtwE4bzVJjjHxSi2jMf3UtbEh4w7K6Qjkdb
3ouHETVBKy2BzHdkcFl3nUVOLei9jU/CDuZnN2y5jS13LH0INpnStoIejvfKv7LJ6/tZjo0D9dVt
fRCMDmjVufbpR2cEg0kSeFORdrPJcnG3O3/83roeTEJRdlWQ1xoFdkZhtVxUCxjus/MBN7CNLOPm
QCnIgu6Ov5NP4NOBTKGzI1iaWt2d51ceO6k/o7jRBuRsp9CYkxZPj/ke5I4zf9gxIqsA90H6hiCa
wY6rWv62513r2wGx9/5/mJjEehn/fHNGcNvdPN50ocs5syfdgxv3H4n0P/Zs9kVsyiUkPGvt3Hvk
bOuQhpUSQV/8lKqXG8GR7JcKW0acNSAUPEkUqgLSkr/hAJUKOsfGdk4ss+5N8hzvWGDuhuYCIxOJ
QwGXrA4iHZjaDGZX9ak/sPayWaj9mckLtUBeTSc84HYWa5RFO6f5gswnMbkc934PdpjeFlJEO5QN
LJZ1g8NlZ/SKBLocLQlvo5JK48Oo6zFmL0OWg//4ZuV/lIs+ANwwxl4c3Rm/IKbhBShqlHeCX8yi
PV5ru2nlFcNlsySjWeqEyg3oQMcQ+9u+xDFZu4RTJGbQUN36Z/RJtRjkRBB/CAQ6yhxrUDjhnNSu
WVUJNX5z9Wbbpv38LsBl9AkbJyQrQ/J3bgTI2TSfEksabMQQB42PvQiP66b7SBgLzyiCF105ypEo
NxqH1ERTSjb6pu294qQIcgJS3XE+McgrRf6ssI6hy2KpbNTRy514N1thKuwSDq/MwGMmMnEyB+YP
L5bGUtwQP7YFoKgoL7vS76Gww5JSM9+LC1sbh/lfbpuNgMOhpsUEtbKENNpNbzHCOO5IqYPvHhaf
GMk2sE0PJf4IH/4YT1KItUMwmwUkJAhhzoO2DoI3MKllPHaeJOnTBfs5XM01TUs4KVOFNc34huvR
aTDHI1+8qlTJXP2992wZq1wxiQX3rtjbU2PrAf9vazUscAG08GiobUj9RpKgt9hvqRaY3VcLl3YN
uTPS9NB7AXVYyQm4tHCcxPFcUb8Oebk74zA15Jp5E3ZEgMWGyjzZkMyABIERues1albwDu6hOGxs
bhnUKOj/sNYsqpJJxiLKaj4ayQbGjRR2od1s4yJHuOKMnwvNUqGdtjjueaEdxL7O6ZWsjGgSwCtT
UBWn6eAowvRrvEJVo0b6QkjFtBqOPFulmFp79vyHO5THq4knftciLApaEr28Sc6TPmKKXB+NAuoF
d00N/71hr51hU8Y+1y9Py4fikddwIpPq7hrQ0GIiICW2gD92N94nypOdj9KhYliGsLp+zVO7a2TR
cnNjzU2VPecw29wZR7zrL5lah/a6xkOdsXv+l2OxEcJ8jOHZn5fr7cD+rSsoM+10V5EN7CfQ35Lg
zaD68NkGf8zCJVF4QZrpFQnML2MfwJq5Up5jBa7kw08abtJbm2e2//EixBlLncAPMuAsWeFUCaRG
K+7CryRmu2UNUTcoQu4Zni5XLlLyaU23w0tD4HJSnRsFeGhSp86QPxztkY1Yi1BtKHitcWalx9Oa
FI6LPnPuF7Ztx+gM80s2rOoYMmqnThIlWfTb9RRVniOhAnl8cxLwJxyQofCz8d9ZteDjyBRy7YGV
OavZ9sgL7vwuoi/tVNpCtP5QhVnvnzv7dUCAnR3O15NMHE/qjE6HLGQ1wnh7mt8MHIV0Kzg03o5l
nnjbCOCBkMBZ2Xu7if9eXaX9wmGc9FIGLU9PHBhySR5rfAdgdFlTcmGIP7kIyxsgBiShXBeY0Y2m
0CZUd68Y4vf8pTF21q3VaUPV68reZ6h+t/7fZrtoVDiSbPvYIL1Oxi6jQxD0G/WS6LzNRRBmgdaE
htTUALtWTlYiPkAA0Dcz1bSPhPh2RZHXum9VfK+6JM46irIUCY7cpdYcTiWgaPKU6s7yyWgEsPXl
5/Decu6vUWCU6iVbmurKliLIWt3DMGkVl6JkQmTWnAjqk9oAO/3ftygXyANDaHtmN0p0FfOUbH/T
+LqfAfyDej2b7+vnA9QgCi1Qtz1T/EiMoF6YvDZt5/DRHv8vz1aP8TOyShYGCcho4IjFG5J7i3Y4
DoShCYcfiEbkEpt1yNhLgUwYCukNdDQflJIP6qZTU8N9cFC0/jk0EvdgB0oW4ewjpKxOYd42hDg4
1sfDcjIPl1u4DY1B1/QYnajLlQ83fD6YaMSMgsm02YnP3h2qKZCUYfOBg3TjTrffZaY0PYJ8aWU5
TV1XidLnLv4Y8LNyvFqov0xSN7Pcbh4dtqoRBnQ886D+X+zpyvo42bA0j/J+2zc/MR5BTaIMCnFc
l2FVXJJ1pD5cSL0X1LM2pHcgw4626zLvBiu+ERtxuqQQWyjDcDqOHKAs1wWFyxl5lu/YDkC4OhJk
WgVZQ6w1FRJiWipKP7+szGDVeaaOMvTWkor7O+IcOA1mU9UvOSPkwQcyEhYtIWJ9k0/ZsFpJdlRS
zi9hinQl9lOgJ+lBuxoUS97cltrUdrXZ3frRprgTpEcO1BXx0spG7xGvR0wvWw85X2PTY9Khyg2B
Ua/SC497YOmY/DiUvbezJOUaDnoSVbP0cTw5yLcd2Xm5eNkqW5IOvPpJYnSQ/xt9lLtAf7kDxFFX
AVzWrp5ltTmEADpRDhysoLyky1DPbAlpkDmnDwHfVlzE7NYTWAvyS30YjM8Ri8A0QDhGuqHsWyXb
YnwKDpoS3yuck/D/A6leqz5LK0QrkbFdhqbJvfeOL3Tsoakq2RXJ4F2ycV8NwqiAtn5udJ/vwj9b
7r1k/iIzF/V8zcQU4UzSPJneulJOLHfv9xTGddSVawoBVA33FfkH0NcOkKra6NcwEaLCGQxZr/FG
XITOBVpx5DmOXgVCytQYJR3qQr5omH+WC4RHUvUNkkbxkIgD+1z4/UGH0ljA0lw4zShg3/RwGPzc
q+ZijJgPisf7V7BDV+YdjHznUWXCfO3erdw91ThhLZ08/Zkws5VXWlbNg6UdrsB+Lyy3I4AdeKgm
wS7eo3nykkVux4zS3hJw8p+C524EMM1kBsFzk+wzTUbz7ZSucmBbfFFKyPQh5BGPs+Wyrs4NT5c9
A8lCpn+jwQ1aiXrKQqsrYbew2xkxRgjwF7vdmXMytcLuvJxIhhAZ1BXdfpmpeDsrIlMqDULlrAXK
cvRFIWsyM4Ztw6zYqd4ZilThUKEm2JmQWKURGDnJTtzMgrKezjKq3phFDyDMsIWyvAB97Nn1x6ai
24wKZVYP3QoUTSZ0ONsVgwFnvexsoY5TMJvUaVkGaCDO23rXeE16ybHx92AxztbHuzqe4wfP58bW
kGkDwE/ak34MfDCk88sKt/bzQjLxR/dtu1ep6vduV+/1gfv4sl19XfgeKUNMcAXmCAU1C6A/90cI
/1HFXwR6piD0z04I4WC68wodv810XF4xojf+8u/CZ3t9LWLObwnpGDJ7huH8ymiSXrVSfDntgdXu
yB0oKmiQeA+A4PsQ3lMEaXXdgCZO/xPdW6v0h+BR97m6aE/b+KYFjSlKiTADr5pusUt9bdOl+HUC
PUb0ovk9axjsY6DqqsZOKbOEuyXdx+/vXSavxhx3mwel9Uwi08NjCFGEyS+iqlr0LrubV7iN6c/9
iqcl+vLqtFEilC1f/eu158/+45cw9CoD4Q5SsF2716t4lfe/STe5vSJeZ614LCUwVUJNH+OpPc5j
CPIaYM8BGoC4JMEsNCtsTs6jrBHgLfZ7SxTKazcgdZtIRYsa37zkwfunlTm9w0ZFJcVlD3Lze7of
NY+zffOqdjzynYGH4ho+PkSVdkK21j2nisV88im/opRTnNoUgpVjqSANAFCo2uED5CJY0/Ortngh
eXUeNPj/MxDSoJPWprqafW2BaOCr7KTAurFkccGwbHkn+Jrj5wudxr8Aah+RJLfOH3/6YQsxqoh/
Vn8+V9njYNYEaDdSxlEvcL/sLHnYtxWAixxxZOD2NipIKgREoUFJBAkVvvVBf4HDq38bC7X8UEVP
e7h4vaeZDILX1VQZBoKImP3PN3jwGBIWkZCozVoLn2AG86yxEpeGaP6rcimBK8SZReqa5FqHVAg7
Lxczq16kNUfKvxnX3lE0yUtF2xAApQ/tl24BQ1NL421r+ZlkatmNOIyCkBXauC8VdpV9ciYtVM+d
RszkBUWTuZ5HkBecyj/FNer5e6Vipw6Tn/i8ZTfSYKHTfhl36ejmIxugialXjn6UnfXm1ncvZ24S
a6LziNWoXVDK/PKPnBsycko3Hvjkz7af4nZnCcKIEKEEDsoLNOsB9GTjnirxlRRmJla72q96Ifb+
90d4SGEYhFR74dYl8pigozd0YY6Bz69/AJ9PUkA3hF+3kivkxjuRg+Yc/SlFvn68JF6nVALMXetu
zYcqbftcXj/+bQI8Om9OiyhnG3No9L1RI3EzENh+TL59/5MA0nigg4kO6ebkabDqLzXYxT27CkMZ
k/0TY5Bjxi5A4kIDUWoL8KrNd940iZweO8AiwnJKNKQN3nYH4ceCj4I/zHwGoR2q1Mkd1Fn+7d1M
GSoGkxDscdAF7K6+eQJC4DFt6ZpcwfGZEdCmBQHOGzd+/80dUnrfto8Qtt9SOE19rNXUIYoQmzv2
j1bU2ywVouNJULXN3l6qwq/blyyBqInOpEwwFtKbBCx62zxsWa81WLjrC+GFhlZ7FjJdsTu4LSew
9k4WyvTxPHlcpodeza0AiLyTMvRLyX8SQJOsJs/DoKiuEx0W4mRIN2wCIA/rrGGEc5+l6DfHdhHt
mA2XrdyTj7q6mMhXvTGis01+72hl1AJyRWrJ+m4L6VWu/qpMpJ477BLgdjwJ/UfqWrIfcAz2zwPH
aGd+dYYZemLaDSRzqh2WQesqlxGABi8vUn64ywFHjdrsWLRiVNoRQdbsWFud1ni1gvMsy86tbW90
vmcjSjHUGFeUBGWnGGl5mKVzL0b+vhSe7j9BQioEoAoaVYIMx+7z1IyWqu+ssaikPwFE1nxRWVnv
5/366wi6U6lmDT4GBkFLfxMz29YfDAuEpC5u/ocx2cwnIjyuDw6H0c5rTPzEI7jLDXNX5re4DO5c
QgxH4h1USulwkkCfHE5L+r/IJxaLyZV14r9suS+O5NtctrdAQcRwKj6CwXnMoN65AoN6+H2B1Iv2
ddpohlWEn2XSLOVTqNckxEi8WsngUKokfp3vGLY436sNh2hlY5ULqrn04Q5ND9tsnBXQKUFv7wUK
lv0XKdyVU2S143/2u+u+gOzrVtFBt77AUfujv1MPAk4zjBiT6auG83kTs4wybwwcJgf02GZl2mVY
lih92cVMCJ/F5bwa8y4bkktsG5H65AaGVN+eaGVNWNN+H7OVHEfy/cS2gTWfVWAyvraStQIbmw9Z
C/An6+7D3zHQevkg7eW5W7aiUL6rQ6onrCgfl/56gaFXQ0pYYOHUgd/zQSOtqnd4tpuuACIZuQEn
O7MoeLIlELmk2jArlNcbVjPQm68IP9lVhbe8DTJnAoZTNOy5rPXrYfcAVEZiyKVY2kRI7LXghZTa
FLBiIYL1vNvQ4LZ5HJQThacxSYm6HAAg5RIboKg0fgiBazTPELT1a6NJoQWTww+29N4ggP3CcflW
GgvaM+3PJ37DdsluirYeKEKMSK6yJEStGEVZIybva7UJyvzDygYYYRDrlZkglCJQ8Wek2le+jkBI
8hezPz/Xcrqo03b9GQwByITSYtY+CO88JMWjjTt83RF9GRIt2KH9NbPCaE/sQ9O8j/BRJ1fXHpTJ
toLV7DEetvN5sB2jXREHnAnon2nEt8NuEs6KRaNfZr3LWOWb9Iuh54vmgfm6cImryjXcFODZK4dz
VVrFCRHZ89yRDXYeyQR04YRJU1DjQ2uLkCrTt1gpMMm0ZY/YFUZ25L/Hhkr66ivRaftN7+3i8Qkt
M11IbcmDhiVlQ1O1OQTR0ubD7XfOg6O3VIWCBO9GawK6FEQ0q/Jz+JdeIu8I2lrXfAQMtVKhaplf
Lxk1diE7hYNR8UkydDL1WDceIwMtRJ/EXmuCx49zdg9cD2EKj+WSBZDhoAvtKmWPV9TcTj2eqy9B
RAllp/4FEG1p660BX29fdnRs0jmS8GOBdhNQyDpGAX6URbXmVR7eVdMzNL3EJnfiFoH89jheYcW+
3MooV6LmsmeeUenAEv1pnVXNeMOWawq94GTQDiDEwThO2ytUDWAXUqN8JNUY05c+RKc4EQkWSz86
bu8s3JCcDekf4/cMP941TFVMBFCFOcdfOciXg/d9K7HOXM1T/X3Z4bJj+wJ1fkoyixmJiqrI5m9D
TyAh9v6N2IB4IsqEQlPthrUCmtlZ+AGaZmJKqY4WoqSFAb47y7DE/uD+G9IEOw35F6+7ZkfqZXGl
NJOnegwWg4bsbGch6zAiDBPNzvifn4oH20ON31BlKAdV8p30NfuGqXGjtZyWbrqWwpTPkx+yCgHC
j7Ac0NEkP4uOvPyohLG6WyJck+hE0DV3uWghLg0i/fPJsppMZ2nEZz2h0J6IzjMbkk+R10LOQcwS
RIDIMoYbhJrp8Bc+ppYqrtPRdD91mMdZSqUJaFmtowBJ9Vtv/vSROx+TUL5r2la9OC8RuqbHVfnf
9q10hGnb01cpuVn0ksT28Ps72W6pDcAJdYmeqDLaaTbDEvplZEs4HysTYG9AVnVHIGS0UN4xgqW1
HCJzidJhMB5w/5sbMxtljZGHKkLjXNdk8hMRbgK/LokuzVXBHu736vQDF0dKwQBIIrVrHfMu5y3d
zdpRvp49v7k9j/i54gZfLjg89mJm5BDwsQTfN0FRQsqaXpfZvpc38+JAsFr44yR0NkQKSPVUs82O
ZDqAbeXeo+SNcj2soUf486/yg8FEl5uaMqWAysK2YF3IVnAQGR1dhTgfpgrBL7u8+VCUH1PX1hub
OZjqDYZjCbX3/pbmoBlTELEz4MWPgc6zMbMp7afTWuwsqznv5pjWW7/CWHYZjZb1hdMOH0CI1Ont
5j5psVuPbgl7ZZBmpsnUwJEtrXuSB/ODogaxswD0hiZitt22ubIXoOtnFGr9Q7n5eJ1+BGTDMYbH
QmOoXFzP8ahfQvF172qiQasM7npVKFIAlzRn9rTx7xReWbl2P1qqyUeXOgVc+aZir4IYTrCQx22/
+xK8V4MgvZQj9XroHsI+SK4qfI65dYDL0QQbqDMSbraeryg1mt4ySRAhEyDaGmVXTdkzwMeHm8/P
Vl0x635QFmLb91IseaBKgpKtKu2dpMz+hiozHBwUm1QRCFlZuaPvPJvLgw5TLMRm9qYwo5kCuwZ9
Mcz8mQdEJjrSljENvtVMfUoRbPtNol1neaPxgVHhGfLMaiKYZnSaxtLYxQWWfghcNMvOsNZLjDFy
sLLdm1VoVm/IurzsLJH82LCu3P+pQ5WGf3RWCiRxVXPPCBLL/N7kyMYgMHX9y2D8QTuGX4PwmsWi
T45cKtOQbyhlWuKGf2KFb40WYBR73Lpa0dehOyiofe8/FI7dEuj6P5sY74Adtyp/2gdYFr2xEMAN
5Df/d6Cmhd2Skn8Kdo2B77nIWBqHBOrdCHCK8zyrex5leswy+2YBhQSEzpZARQ8W9eMmLb0I8y5F
U+UK9h4Q+xdSntPKM6GuCItkwis25WCeVJFLCa/jgQ/ythR860OQ6DTTTv83JrWsDckOlh3xEm6J
lmf/uufyu8HHdbjWDsfshXB5rQN8ukzz8eQ7INclsYfJs6kTEMyQPtux/AZLs9e4XPplD2VByNkY
dKH5QPefWxeQCAaWAK364rTniU+OZ41FU65DCmlwcwOe19Y+2Pbz21fVvwku0RimELYGfrWSkh39
2lTdNiksbTyAzS4+jMV+zx8BBeeEn64qhEnPEwjpinfjI6oCkjnenkljd3ZrafP/L6B65yq1O81b
jvIHzy2IaAdhzBfnF1ujeZTIXF8i8IJJpwepy5f+HnkQVTixf324hInZtUWRnAZVMkBt9cC4nm8v
n7Q3jKWljt8RxUmGAvYzfxWXHvupgtJ1d4x9R/hXnnlVVloYkkdB/+MnjmA05hdy8HTuXluxjuCJ
Qsc1L5RW5EgFsVnytKFfIVghbJCbf0wQesPB+7oFqANN4TRWcwBTsk5UEZpO/rRYUTtaUbXdeM5h
dulNnGSQ7y3Lesl0/Ibn3TymAhv8Cf2tzm+HaRLSQ+KpNI6aw2Ohpvbgdj598haFwaXrnmYSL2fw
0hBwVxhEEPYLdPXfRouOKfYyViZbagF6uMsdh8bMeumP/4IhsqvfC884p9VHr2kO9mltHrutH9mS
1FJHWJ+85WgF5Db7tcIFftHPzUhOzu5wV8zEwZvKkTJUVvRelYX+VAKTPEZUm2DPvYPkMQFz/CYg
Wb2+H6rlXkYyptJvTpp92R87Foo25Luf69D4NEk8ne4r5Ot1G802f8yhlEUI1G3H3NhW7DfyZWmG
b6FJJH7BcjuplScDFiLiKVWii7AeIpS2yj6BbleOleOAQKwmSUCnpPdHZbOjhdALHtxs50tczscM
ABG5KtMw2lJiU2TVK63zIv0O2QrcTp6n8QB3cN1QW2Wf3jRqpOgJBx45liJX4qc39R1a1AHzHc6S
XV6YnOSeu/4ew8T1YR4zoB3tHi7SoO7S1OmSVhNl26Xk9+V9iwZezMpPd8UhyAjMhuWRaIBsapBF
xdj463xdQPzHvXNyqjBdYNlSJWvPZLS6rKHHg1oTIxvy7PX9Z0mm9sDlOUb/RpIz6XlHAEZdHpT+
NwW6f0BS1WxqZHFAHNAnY/pEj4VaoUOx/j/ZCiYsqQ5f5EJd4T0TXWSRPcFFraiaMQQqHjBVf9my
NGegqf3/ACVMLAxBC0wvs29kYdJ0kpRvB9Icn4IzGJxT6tuxrDCCWfpgK0wrW7UN2TCiG9gpt5z/
/NMYe95fwJGRqoU0cquXchx73+Z4uZwLfS9AhWkQjRfRwLoW81R66iITOVkP76r52q7aSNrMuVVJ
KS9SspjHn2gRknFbLcOwC8SPAiTIJm0/Ej127IEgEiKU8mrfdlEzfji7StleFDX8a91ApefeuxEO
Bshwa7+DqtPm69pt37GGH0FMg8pIjixbE/DNNBqj5Vj5hLtV5BDjRkS6NuRjYejL0WpDFGvoBL5f
Sefwcm+yCVubfaZDME+1IW1g84g5e37Xwgx+4XIuH+aVA/C/77GVJXTJdDJfrDS6dhRllpeZAg3S
ZIFBCqGBer9Mnffir6HqYJK9ZWoXTy0j7hoIUMRuG4z/h0WsJiSTWBy8T6oJMiIygcVOM3tRsihj
buRIWOhwO9vcL7gH1ehvbQhU4DYCwy3A1lFv7NhFvHixtCHT0I8OIr2sfWVmIwdk5z2ew02fnthL
cc+ggi7TFG0D8ncLtI0zgCBc8sFvdLzBiEsZXK1nP9Vq8jKp/9VX9s7KcBtg5qVgKARfTRAzE5TL
zj4d6bDr5JZmX7nW3HUbL+X+aVZFidxZEglfILrB4M6oyXTX9l0y9rXpDUrVXItUUq4/VAvhrCgT
HYee668ITyReEa8Xgzn5rsjm7BOspbonKp8jU8mqi1IN9CF4nnQbj1FJK4szT/q6wzGtXZ8vnkkh
dYuJ0DAFs0oJvlRmHjyuAvZOpJvP2HK/6gI4b6H6eXmf7DnJ/BERyCBz+4iGT7hP098CKm6uWOU9
LXVogh6SFUbxZzurub0PWOqFExyGfa9ozV4IlRpPUl2aGvF+fA06FAFZrByo/jVrd+/B+TziQOa4
mtFJ36fhtmCxCNa+X+LSHIEFblve1JzcCv+W1/3MklgzEO17f1ulOnAGCve+RM2GQIY71iaeVZzu
/eoDrjAp++l0K1OHVWjEXyYe5ZnBgIWbV3UJ7qZdi7o5o5MZBUlvXx8WJxNODUMzrgUPFEuYSPar
oZhLOejDn9sD1QEqKajktTZD/YpOc4DWyCl1Zyh0icGQA+6Cpm71i8IHdkdzEBC8vjiQNaFv7a7n
ZOObwTXEgwvRG5oDcoWWcfxt1B81Fl9cb+x9YEr3k4p9uYSrWDuIhPm8/pdedP/8F6g7OsBlJi+v
C70onn/lRX3oYHajy4XC88l9bmFaFXsHAFiPVSIjgji1eoorbzZ6lAm8pMab5Yho/QrHTUq9OcjA
3HHR50xg66DVx2+b4CiWKb/pAoVJYXbga4x7oNYO+T9KBXa2FNL1NASx6Lio5oI4eJrQ2/b/TNF0
0ytlRYPD5nI91mmCoxFQ+H6I5OFbizw6FnxTME66OuxQMNlNYkNaundKFGDgPFmUf34X821+xMDI
pVdWkqPzW+pfID34dDIzCh66WmAm1D5TvmB7ByMW4wuzjuXecq6DauPZyc0PUrziaa9yNwyDcUE9
xI/wxxQSaz24xCg+X4HIz9/0LndLyE2uE2nRYEGqs47VOrGuG+FvaCmmlnO61aBnYv38bg5vayUG
5RPEsN/D06mO/BDxYsdKpZJkevCQsjGqZAR7A4vS/s+jQUqovxd8mlq0OVvvXCnkDcQrMWUzOpbg
rnlaotcY2ssETqSsteTx0Q1HHTdjYc1eGq5VUpgme9HJF35QuytDHpg3qlD3HAIabxqqqOmXd+sz
rYS/N43BoaGXwNC8KeBKChQOBrBTUgELhTkgTj/IRUEErr6oluz5eXwE+ZARoRviFxUA0AO+F4bT
NX54EUqVzdX+KNvqVI/j+1iws4WhJSL98pPCYIYBNCb0w6dT+z5Av910+x04GkuzWyeKng+FlMju
WG4Lrey8zABWDtLjjyFsDKSCwI7iyyyVSDoVjOvlI+K5vVTKjrzygXPOSIVtkJs6cXA7GOUbdPl7
DVqHj0dG/Lq7XQ3DFSIxwhIvY/njlZYEbs8c5muLd1Tbg7Qi0kOhEcKm5vdbcvrGop3n3sHtpDYS
dFSpXdhRTtP25e917I6F+i9jlRnSW5DOltgxpAZwxsGkBD8n7MOzigQ4OlJZ0NlGFOhZ0K3rmZ5j
ZQa1yxZbBhBe0qqNUTzSoLAIIcN3xg+NGyY1T95F+/PMqlcpnEaUseM0vlj8iwiBlh9dpHmv9+z1
ZssUW8x/ttSMH+LxpFFLNFH6Gk4TgX/7TI4+njutCtGGpWUkor3yqqmgfoSH0Fk/PY538tCRd2I8
qcxGkeuD+fA2GdHXgJ82XOACYDB6VICbjX+1Ja5iVQGDG1x/EXQ31ZUKQUERMnxwpZAwJcbuMAsB
QFTHw2q/SZbuNu/9cu3zyKpwVfbz13yOErYU6GvyrZbGNucdH+/IYeJJAlIicLJoDHOBm2dNv2df
xLblvtZJsTOc2lRxgfOKkKk9BcFmaRFcXcmFNhkbg8Ebb+aEU5r5T9mCc1C+rX9RzxAnOKclTI+P
urRv6SK035JBLixjCrm0Wr5HFSZUL+1fuzaY2cva5wIPvCabfC49PAFLPngVNUpGatOfvUvjCXY8
5NFYVt7lJbcEtAcrQuAIG5IYIyABH3F3ZPp1c+mi4gKARwiI4Eld38BVpZBZYhxVTPYCmabUP1zf
D7NqsajqF6P/ULnNQX7YHRV2pzwtKBe4aPmu9qTTv2XlzFkULiHh7qBaNE2WSxY2MqhEC02T3YWf
pN8kFoEGKdg16kezu3len0AVNnuqlgrlubM/Bd3vVbIdtsIfmfRoO5B6utM6hl4IhvKywLQwgJON
gHqCkEJxrxwaMhJjBCb613V4n8ndRX6o/R/afm0quSUvZ7uiTSd+gNxfRuC5sYpQ29MYIJSUysjl
/xcVeg4XRY4w+GOwGPEk6RXpZ4qy3L1bzdZrWhYKU4mga78xa1bZZVjROGOWyDjnSme2GJHnfnl2
rEW7QczT5r3s3uTe3FijiE1BNH8GBUPgi/58h7KJE6cLGUyqz1BkCNkWIMKI9/z8RalAcGz/E0IM
rBp8MumDjLk9YywtVGQBb2X9GzxWhq+10PVHkh9sXo523Hv+8BIW5wyOGmRwpme4eG7AUrzCoBoP
wplyqtzHFEdVgm7qwW9NOx7N5o4CZMEKvXEjNlA2j6nUOUpqboNmXWFcWetpmwfm+yQT3agpqW50
1ijcMxY0lzeIdBdpRikgvDv4jppxDjlgI0k7BRmJD87b9AVZtkx7k2CfAaStMxTd+WmHeLrs2tXA
kjfBo8oEgr5/W4IIZqnIfM3U2dhtwDd6iWL1ADSAQVfuAfexWJMNFhoMjMX97iznbisULbm1DE5g
VNXBYZyfx+TSusIsbTXoORB+iQchxNls7gd0QA2PcukCNJUFfnUH/tJGPoobVWReBHVZYmgG0pAe
zK1tOZwRkabQVUtkYs3dnYOWmthVG6cG6pgcrMwZ4iRxuBFjHfjcs8ElHI2COhzA7hrzPLbfAvJJ
d518u10Pso71H2ueE7Knb0vCnKiNCl2PAhR32p5DuVNNOB+axBDTFZxOM1B2eLsNpz2ma3u+d9VY
89cpcQJdXBjvl8toJoHMioSM6E1ysbBS7P9QprBESVNGMmemmQaKRwicXAkGZGlbnh5XSX/umaov
TIzqpxdk63IqhVBm4F4KopApw9a1wqYzz+5z2j4PbEV7ngYPLxlQgiSbM3QkOEw16qLmwhazHIUk
e26G6SJEDYx6TRjq0uzzsjg/qJkOjV29P42OSDqNiNrBNvIoMIHd8ArKxdjmjJwnsOzUYtA2QnLc
hVwxdSPzW/ZNBjAUK4Ne2jThP0LTc7+uy6mukb/Sk5u9XGzBeKpryU3VBSaoOYkiRGizaGG20vLW
vKjb1bXW3GqS0xkpSpWDJsIRL0dyDqPdvp90B3A6K1jtRCmv2aUmwewHekxbz/9Jp3PFKiBUq+OT
PmoFjkGPv8vsg+KqqfGHnxzy7g6/VzcWTlObIC8Z5rYgJKVmqUqm2i7oYm/z+CZqH2cH6MdDl7Aa
Xb4y8STLjJhE2o5bp4sse5hO72ffl95yA9uGjG03W7rM9lxK1AxaYraAys5h3ng4SeQmK5bojKQ5
IcJpGCpU+6fSk8pjJo33hdj0rPFeic/04Wh22JfO7AJ7uOdn1whwNUFuXU4ERAVPV8rYhm4s5nka
f807raffFQNJltQv4dxg6lZgmP7brT5UJSqmTh7Wy+wNXNCCU79uAzLUdouGMmpWcYNxMvNJ7HHM
LinuKdYhDfIQ6FZLZlKKtmdvyCVlRsecUflpUm09Ps8MA+wlkgjvsqI/7XaPyXsrWHMnUzbHRuSC
OH93fvFX6MFjIRkEJV5bQ/bVI+JDULjJ29m8HHwQf3/H+jpFqds9vFuEea1HghRHFyI7FUbR0hyC
/K+YbZjIIl1EtJnFe/HJUJScMaqDxKgV9cLJFEx8igilhrOwS8NqTIZqorIwuO7HSltLL3FmOMxP
iVzTfvcREWhje+2okLPQsi2z7ySzwMK4sI+VPRKloyqp7stMWm9KNVAoRwq818pUSN+xMP9/lz2t
v3RmZ7dnFFXrmZVR9OAsHZr6kUoRpN+BytADGRaAWsawF8nneNe7BUZE0gHZm49D6mc9uNS40QSH
cqEACkYoRzV4teFADCtxwc5Gh9XxI4Anmulg+5PAjINV9D8TRHyNsNI3HxQbNmXoQPpOmNPEUuJI
tXogI3iuiI1gGHF9TqxKjBgfaA+eW3uT4qf2KKNe51ET/UAZ/jelWPNrFAr25Tfmo2M+QVuR4mOD
7WXyXaNu6aXwiBLoz0Ejias3986aimIHK6GZJrCu6gDwYT9HCVR+8orcCS/aXwsJjKenutCV2erM
WlzO/jTRn3qQoXWs3obr1uzqBom6PGHUXzatI2+axu3St7OyVor1a9+l/wFYRK2q6d+w9tpG1beJ
2R/HM1tXRdLSvdGHGcLTjTopDP4vcukzYBrROD7x6DlSp4R8zjE3qdqRVpjzkBIoheLB/bivZs/r
wGrtd8ZkG4vqvJUCpJFsrEO5zEMTLzf3j6XZKE+2WWOtkGJdxzYdXX+zc5cgX+LTj3Zb1XK5rb/x
rfX0dH7J7nU1ioFLtCJf6PSZGmkf7tFwaFcHYWoT3l4a3zHtzXsHwrqpt8peDllLfij2LYlkRJ89
ZFD0ad0auCHGmI9L60mW0EFm6JmPoZ9mjl4Ts63/AXSc5w5dO28mSm8S8PSwYcuYZaco5+Tf5J6R
oJoEEz6kjR9+IsnXWAacHPSTezbNc3j+C99TvL/5jwiGi10EJ512DdOWDZv2H0Xf8g04+9MwcdfI
CrHd+NRLFbT+JCLESs3BZPeeYq38loofxbF/LoiIpndionOKwRcefRgJ5kFV9nu4jMOYF5Y/dhCM
BJr/pVRvEzbYanbfhW9D93x64KGwQ4xz19Tzm0HBWpwExvelSa4MHwc4Jr39B1bpk6u47f/w8RbO
GR+WRvIDB4iVxlaly3xGO6m9G9txpNwYI4qivLITU/pkbcKPqM14KwFCRQ/tx9BY3cOyqkB3ECsZ
8e0+qv3l35TilX5AOgEUzPfiWxc5Ffmp+0tis36gF7Bqg2P1VX35L4hZamsvEPhIsGXVejXRr3ae
LABmoQqA2izvwaTFP/eP8I6tfpEbCrCHjubJLEY0e8Ey1aCDswIuJ5/Cv/mqBGpoUTlMLbTqV6Iz
6v5z2T1atCsD+oWfXgRndlG8UdWxjpAlJhLhxJtKeK5YUdGlHAsplvMuQ5+g4RWcFp2DlyX3R5wo
HbfrNc/c0FkJ8+cp5+1pnuTNGB7SbjDCC2I+k4OVLt868IL94CNMbjLCNt1YUx5ob6ui7Bifa6hg
wmsmMUEtazsaGj1gtyHPVOm6PGUmgTJ+6NKTEem+M1kAROm5Hm6dDSSnfEkuByNlHv6wNpKi64Px
w9OZcXDE5yPAz6nYpqm5gGQAVLH/AVR4KxfOLF2oz3fbsPKpCWz9pdJ06djsZ0g1Td23bRorWEFr
cnBaTqw+kMnEaR6xBUtH457PHzyndURmBxDpwO6VSZgk2nvfVCMR70orNZkt+AHtgSp66hVRSQYo
nnzIUZ4lSOYsNO+CTxNfjJ8geIFFyaaeY6bckYvn2oWmiB5Oy6/cVRSY3Cy+SZBsyQAIBTNdZzKk
fFemfV/j5BzhhOOASm2AdpxakAS+bOoR/JrH7bd+GhdcTQxDwcU2QHs8e2FVQMmHcTWPJLvn00rU
EuhiJ+Dnkew5LfBdMyQjkysakdWRuCYArJe5GPqkJf8s6uT0XPHBSMPZS3DjlaXCLLIW1P5At7gO
ohkzCVF1SI+G7IV5NfFTTF/HKs8foHH1PuhVlWvVgagLDBYO0jiymQXDEwC3wZRnNwg16sbrzywo
KMKOIg2Li11paZGZdcWjyukhtI2KhBfySBw/1jvZHeEs6ZPXJFJXRgGnJKkwH9xIab5u2Fvn5wno
UgXnqNbUz0tTtItH2MyDdjBgohg4JJHJWn+p3noNHyNDYcplZCkUoA0carNmoIa5rqvN2GOmLXnE
mALgTdS8zuXLypKt62VeRqPs3Zo4ODR6HdxCgLotHN0nv0IrqSlL9HP2E8oc1AbRI6JV7hNvNuZL
/Tg6A9Mmkd3GZhnu23FFEEDc3Ci5m8TWZP2wve+5yWKwV45Xs1TvDxEw5WbFKyl+Kk8+y7sCB0Ue
/maUTa/vCFQILNsZhm0dB03PZhN269vIh4PQvhzolHNA3kBeiZ44vGiyKTRFt1Eqj+nnff94ZMGe
3+1RtsrU27pc8WpZF34KJo8BZ20ZYmDfWcOPutTn+tDKKRVVrYBnBTtM4cwSw4HqYvHHYvP8WzLT
L68x9/Elaxpkq76Yj7/uWdcwfu7am9CfbqshIJ/Rf+cfoP/bY/UpRd8nnt3+3LCOka7UOC3WhgRN
lgQGPvNuO2DFyJNQjDx9amnWFPAxwWfV27kfc+Ja8ur2EXQqinkcw8hdds+1yemXPvRGEw/9BSHV
T5i9AtJDGzAYGNCXrwXS760fvXZxVbH7jXygH8s2QIFXcailZKpqfOmIbfS/TXX4bM67Q98uPwzh
2wW0OYWfN5RuJhe/SexfScLJ3wBgeLID1DBY43aLmtavt4s0LCeTYrUMF9kb/QUV3dAgzx0/u6wH
PRHt2aknGSZIm5js4GdssRDQzjdbqKqIgWGq8qlg/f47Dy62lQfqWneluuUZMtVLSNGu1ZfL+wkY
FuuN13tePSiVNuU9umTExQ/d7ArRtrLAqHGJVhXHvK7xpYhIZtws8ssYwpqy5kFAKpVPNfR78VGe
GtwSvr2NmbwuJwAbpF9Y3Yq6XS+2C5nJZXcysT7RAMcjZQkapWj6U+QRULbIXV48s53msnBiPdHj
/C9DgzvDlGWxf/xHvYdCGdZ+IIVaSGtCGPyL4OmTc4klaxQ1UyhDk9431nFA4CF0CgSXO1+sVd5b
GulkTf2prBo+khc811QqBiqMnmF0JCNIyLBZDdgXHuL645Qfs39RVn91HB000TI3H2Rww924CGPo
yzECEWzEiTx5pPm44SQjpTlexYJDspxXijcde4lESaQslyBYmxkPv2EFTgCdEYb3GY36W+m1LuKc
UR8GXPc+oOowN60uSXVwUGuybwAXEMdPAvVlK4iQNSrbMlsl0vQeLiQStYfn2mQ6qZdcSB7O2ACr
GPLf4IqteyprZQ6ojSaQJvhBK0konkI9HRiFp4Gvd7YDd0X9m8y2CwX4A7gioV7gwlGbuJfWi7E1
KZZbmXeDTpvfe/9l4dmq7ZGGpoRHqFsxMFEpSB/8tU/014ff41eABERl9THDEHIWmXbE693itH2L
FuN5gBsHRsFEvVCfzGqBB0qOoYypeFqzLy+JehCvI+qv5KqJo31FTLauUqinNIug3s8r6Wnz88fM
Yj2tr36dfnr9t4ElC/qcc7ZsCESwz2NNCB7BIkf5JL4m/+2sg6Hu9xGpkKVbyfpSwfs9dd73sXJq
KeJB6lsN5PuH695mKEQ96jTJyy0iDGhW7V0zMQVEqQ9T5KJMoeJOnv6L7x/W/8ALI7CK0Oa/mGuu
GWSwvvYnfLTYmA8REFmfVm629b/ezjBP8afjBNjiPG0mJfgQdgdLFgvA4RWt+uAs+GqGkz8iVCJC
6s9Zk6N3vWXmgYqqv17VMZXZf2s4HsDHC42pFWNQEPUnSFNb87lE6sdcytvaI9pn5oSrWOo2pbSI
3BEi5XW0qvhQHqd/gmSmPpEVEuT/zxRIAksb0hx4wPTDgrSpiBsLl9U06nu5EKrRTNtbWytQkP2u
ovttLp2AXAr78tLVUf91xewz0m41NnryfYGsREp0VwA2BuUnsR//3XTjGgxwLxHm5kf2oaJ/UH6j
3wuxwJbp0KwkDhqsBlQ6g9Lt4srQ+waUUCSFnWUlOqO3JhLnUJeVCxphQ6hVPszTQzPP9fWr65+H
iaPZibmOeBaNtsjClNNeMZPoKmGcSBKxRJ7R1X52jqGJKrZnhQLAthRMDS0SdXuK9q/T7XGYgzbr
YV2b5hAk9aYLg8k7Id/Fbn8pNgbgaHA7pBecRDodPooeRX7LupGW1ijJNDwxioHE8gP0rDtuQUKk
y4B0IcdPZOH6GdDt1rg+tDaZuJWvBUJzWzF7CV9Xo5HFHPoQWHHiijpaivsioGv/Z41j3USSiHni
BVP3Sy44HA7A9gd6gMFfIBklZMiHPdGBhADUj9DEkSoYjYr0Ep6pqRo8Jy2gkRbaTIVQyLp5+nfr
BsWtR7aKwrwsW/SZtstqC/SzuNfM1f5U2K+9lUv9YEI/rqJGTP3mpQYeReuw94BhphBGZknEafQ7
ivXi2QbHZsAdnAgnCES5qjWSeI+ApDvfP7sDS7IpYc8ynBJ7eSYBHVErS6XnPJ/NaEy1NTWpmpH1
6XB4bOX/CfTcFAlaS0MXsTyZaGRd8Jj9y0fMZuGhUNLy6uJDnH5K2d/zZrMX7l7vgJfYs7INFAFW
npTOEBAeHiqbZwzax4Aah/WsQed3qyHHLaZyw7rh9rLAa8S/yHOKOhBcrwDv6WYHDegBJ7I5TqrN
+KKtmERAa3hNG0gY/Ao1qffid8d5Y6nWaH3HfIM8TP2F0KdB7hfHJ2ayAotDJNCQ2CoVPCr71MGA
xTuIcnOtkwd34mVZ74kIWCYrSdN7fcUCox30T7qh4PhILelSmr4CA2lvsQBQjPB0cMHunaGHD2vx
jdnNBhli8VJAlr1W2AS4/95J5c+GQ/YdThJDuLWr2k9rUzOhvz45Yr/8R7mAlkaUmW1UZSSx6Re+
I3lPur7sekT6k6FzXyLkND63UcDpkrvBMpDSrTFukdgWFQY6O9tQ0f7HFzRU5Ssa80gQv8w44l2B
sMfomcSgN9Q1aMmmokFKq66+SIy6larxVVjiVi2JWXIHdfPHdHwyW9T83KgFB+PIF3X6HTIt2NRl
0GBGA6WPNw73OZbd+rgmS2UB4smx4ZaSmsEqYF7YiWZYmrUqSyw+CROqnoDN6mAVHBf1jQCZGqZW
ExJE3b3VCuIrjyWJVhCjc/ftkwE/X9DEJLGqT9QjInJABniqMVYYNbaaxOkfcT2FqSJB46aSM0O4
VrWbqC3K6/uc9o0acyMuoK+q/l+Ghh3RqKHx9MD/ww69P4vHy0F/S9ot3N0v0a08qLM4TVAmPkVt
iNm2JAvT+xwNWqc6q55QG36LpwC9R9/6IoMpGsbOPiOp2ZDikAdBj4BQTqGswLvTFy1o+U72PJgl
dYas1jznD3fTS1ndwu11hYLMZGNBtbKyNKTtaNszMj+28SQVqh2L2IkOOY0EeSONfThrerUzmPOb
A8nMKGZWZNvv2g0xFr70IWzafXoDPPVOG7dJWBqjma6Tvcvn/GzDo0ZRWC9WxMYVTz75QYWA06w2
D5QrECcnzB8lBPv5Av/JUflpZt7UtjU/OUkX3Kl4ZDOCBJT+K07m5wZEZYdRZgnvlfXHA/LPX7lx
zeu21Zr6Cr3kd4qqpAw53OpgVbabdN/kMau66TqJnN0f0o1m1bc5TygqxJRl4Dx+oabeVgQp8cgN
SZPfa4uRTPJ/coykHLbaAomY8aglAmoVLhjNNpQumCw7qcqnra9qZ5jJiNqNqjRwicawGSOdyxi4
ADpUEyx58zJKZlZOxyERr0Njzgk3kf8HXdQ36gzXljQeauEYEmO6Iq5bS+HYTN5VwR1BprbwWHQ2
xjcXuVjVwIVipe8jKsPDnrJ22p6M0IWYqMwzij4WxZL8HWKxsTX1oUyGCBgCy8qRMFxjqJxZE1OW
/aeimojKChRBydFg2379ykM0Xl1DZkWi8c0IFP0rHHrqHycbuVmzz80KVjzbJGbYq8liMgGD0IlG
+wF9Ec9pFSUB+Igi3KAm13AUYYIefivgstIHHFBdR+aEy2RqarnnyuLhuYrDCSOl5rIeZx9HMBCw
eQci5tNleZlhAyd9XWMdsoepwy7JrcNbv9zQV6YtYLQURFHWagbXYcr70IOjJCdYeIqShyVem3eY
7Naqoa4KKmxH700DOzHyeoLMgc1BlvnE7ayKKlmTdFdxnfhEuBcyvkkpXfd623rOwyJyyQpyDJXY
waP+UZ5EJnVfDcIabNE10OZtb4IGouhzpv6ZqXp8QYS/w1L1QuC8U+EHNDkOdOseDODdwV86ys+A
RwY5bIC6iEjvfPuPYHgMy4qud3jwyEP44t5sa5ytEclNvX1eHz7HNIV9eRLMxqqVTBg1sX2BYp43
oF1WbTMRsF/TJ6i9PQkIOsc+ZcfsuGky3TIMbgeZqrMa32PKfmWS1QO0DtzXF9/rB3qTwhh/I9Jv
s5/dusssNY0qmERQhc4tLx4GkvyQqBR63WAJFbnzT/Pe2egAMXjkrPOaRdxSMw5TKDGt52ScOAxt
+k3VOT8P+AYw92ZNG0zytGOdJWNR4R2CA5TZmOKCLWULRijBlLPhhiqwFOQn4MqQDaVCPdwbMF38
wz4Mf3BzsSsHmMnvAgT9wf1pDHu6xJzdXciSzvO2IQ4v5OUH7WGLFI0sFNnbcru9h9HMvkmPM8Mj
ei9UZeispFj5uQF+c/6dVlA3m6c9xrs6GC3GnccpLoEnI8btY4R27gPQIr0Ob3y6lktF5IHzRouj
M1O5hXqS49KHYe+egiT5GltEFsgVWds/vuakeFayBii89q3zCHKIt3Rqo/s0Dv3P3xojlJiAzKxT
7kzxiwUHylg6sRiutsNZzpKnKOdwh1mgOtQEXk9WG9nW2qrvC+YngGazoYj8IBjREK4gr9RH1LXU
OwVtl3qvySgnpYWtUIjxZ/KzWNKo2bHc5mdviyoJmPrdp6PawXWSzzjdYJl9dm7TuH1vNvsSJ2+v
2YoR1N/X05pL4s0MESAhhSoC/5/cltx0mLPYqBUUsotcXT4Zw/nLO4rH0qifR+M6+ZeoTBMXlWfD
Yw4BVzxTxyLdIlHoFgzERjegUUL9sV368xKR5AuPzJYrtcSX5/z8xB/jllBhNS0KEYyvoccLju3Z
H2EOoD17WwmiWGsO2WSFc9f/MwPPmeOmEBjZYkLwvSanCCM7OSzTztp8j7HqoE/FEa8GT1W1mNHW
hFZyNnjB/t8I2tQ+zgrl/GjlUgrFZ4e9OHHj42hNolUIZtcaOqBCanUoNZFALT+Q9dC56OF1heId
jT/GlY0XB6XrmuXToW7+OZslZTv8FrbfBHOsBfgKI3GCKdYSQhjhHHdz7Cs9zsVuGWrBhsZkP4Uj
+jlwlaU1uYHoN1SkCAa6mnwkjpmANlRXlGafI5WofqYZgYu51CPKOv6O4hU3U+mWtOi/dGrX12+d
1No5E7PIAEvNJ3KtYDJPaxvpPaGhm6xmz6sp7FFI0jbBgYy5/UlCUr3FbcKKIiFnHsbBgcMvsC89
v4/cuXsJMIfkCNv+jAb/HpviW27Ie9vjel1czz6QzzkEfmhUgegC3xB1vMYOcs6J8SeE3p9vV+NS
cBbFf924LWmqCskr56Z2BKa6ikqPykENMPUN/dPJQE3VbRDM+PwscS8Qbs7C3YBrJjDWnk4n3iJX
xL6Z3lhll1K7BVUrD2P6MSysZUKUfyUbBx0Wjzh+Hf2TYNqAYeu3i4a92X3p8WcAgsD68t1uhyGf
yZIp0DDlsUTdFJiwWk3Du83qD9hvJH7VKB4JCqrgZH2cqZ4a95Hpka72tmRhXAuIdLisI/l2E8fF
k6ZXaLHNSuZiWuVfmNgb8tO6iP2q6jGdRnxn9hK2LckplRzpTNhDaQf++xvY86hCiaDpkc7cVBgU
FP37We2QJOA1SXmDXvis0ma6F1dPtcsZ1Uyq8sI/SckX08ogPr1rG2IOAqlAUPhaFifYjxIcruKj
viL2CMUgPBBNrsClUTSkRH+azmnEcDGSgtSobewoGx2STKGk/zvwskBQRnBZhWSp87r/9sW2Eowk
fLwEqyWAORnS9QkENBleJVN9EdmBhGhZUybYjia6gDGq1Wkhg7uEyGHoLWJXTyMQ5HTfnS8dCgE4
aV/z+pM/UfZMbvjgvhIhp7Vx6o04U0guamrEpCeiis1pJO7+yL0HZNhD/4M0TMS443MKSGExFTFb
zKGYB+6yMuF59QushQdqlF8NRqIEqZhT/T/ITrUo+mQqka/dKnnyCONjDBjhgKpXMNf2z6vi1zJv
cS+VCVDkJ+PPtLF532Fn2J62twk443AYLrj0OhV/o67obhpGoCRTG2+XFg26i7p/L4STZommwtWA
G40m9XmeX/mYtAegpB++d5G74Po5VP+0xxYW55mE33zcVZE8BhNTAUHY18O1PXJmlohIk0fyaTLP
R3+emYNpP9hn6gH9ITBMAtMCd8u1FjVjeXAD9maCDbcsU4RnJjaGyEW1qGdqbBJHaZwcbPq0mguR
jNU/PvKeZVim2rxvszIZtLnzXWWbC6dkIhamzonZPmIA+h0QyZ1bD3CITLk/0XSNC1FTsr61AA5c
YyJA9lfiNwSZ94MOFpYrFiIDSIvAnr1tdtUQnLdR4LUtRGZ9KCDZogqfTEKiQ1Zk6xl9ja7AcE6j
smGNVQ4bxobPaxI9y9iE46K+kkoU7TcMDbYNIknkyerUzLCbwaqx0ozme6dlVGhdDlQf8vqijS5A
aKOm2Wfr9BOeVYain7Mhfixhydqjvm+ok8BONXY8O01R3dgAMBrYD3H3wmfmiX5MPX/GiGQSPSDK
+iJ8N1MtUZ+C1hLFzZc/3cpxOfH+kwiuZql+aL9m78P+TJKH+HqjHr7sxe29mXyftndcxZ9RyGTc
qNZxnuUzde9cB2Eof8gnIOp0Cf4MDTPS7Hqyw4CBFlVKb/pYYj2dRDs85JcYzkdaRyPyjK8wRozT
w5JSdrXv63jicVpbmXLoIUd4wYua9WrITlY7TZEoLU8LR2zBxtdrbtDi0DkU77eDFhvSyIUqurGm
rKp9T0TqTP3CdTcKJtxOo/XqE3ZxU/5rgdC1QzPJ26GyBT2hTdouwZ+jv7EEfu2o/DNdtg0YZKNy
a5zjDSLTVlexbogglU9hFlKohgzmwzVFc7scUjiYEOLBe/2Ks15kwKK7tIzmoxVtErMgWQfFi/Gi
z7tGXyAp4ld7CjUx6CmNW+aXkhJvtTpHv3kH5oLlNW8GnrNYIBOz0HO0gftoDkxYwVqGZu+987b7
8fTnwVt9RCUmXjdtTc5UurJ8JbJCKyEO/RPiGCqZnCzohdR32JGtb+e9RVjTC5S5HUp7+hFP3pR7
Pd8/wXkP2XKR/ATHcrtq1WmGLdhbJf9sRxbHm2ibh8kN7mtq/blbvVg5aPxYp5s0KzwVsz6Wv4i9
9d16KLS6/VczkaTwJqwL5NmYlIk52KqLtI040e6iEjEebSeDrMNmuetrBx6EDXO6EX2PB7m3OwvU
7Mx8vRbRLsbx26qIx9RC95NHN6xugViXORBMUICH4pXvPrEkEZxSig36ZhHAQhczoW9knPl3tZ4s
lIHbhignOexvb6hG5f6uwcPxHg8+vK0+g6Y6jU3lvh3CYumYnABqdxN/Eu3nX0xEa/gMInPvbB8h
0jObB9mcl8elRIqQGwBh9zqDK+vo6ZpNtUxsafqfU9ny/g/WbrUriE0sjo7HbASu5gWKHyRcFMGl
knQCHIQ7nFGtM35aLlCdBzlSfMQcUTUQwz2FhV4oNsGSkE4H/75thzWM6r/3Tq0M6i/jVjpg1bcs
ivL4mvWsCu1DdHiC7bzteiQinMuAoJNn21wmE6JtGsTTWg0gbcvomuuuB38caCytD/FQRptfQFtU
pWC/uI+23X66ag9Lkhb0U/vCE+WgSVX488aBcNw3qyHIzIOv8LTWmgwUtG7SiWoSntyttAs2xVwd
4bgl7UquHkouFccsYE/jGy9+HK2EM/uCGwnMzlHNE/k/d/dyfBVTMGBwE4WzH+u/DyRJw6RfgIVP
VUbc2pvNPKFe69IPa7w862cTWb1u1TMS/vwvpqVaGpYl+YzWG5DK1krPSEmEVCxWvhNdLdxZFtIN
LjTYYbvwxYpRdf7IrnVaIACHaDROCqsOBd2w/6kP5wEXDL/fhQTVXYQo3fFXvVtK4vdsKva5dSsz
CnSWROFzv7rFzbrqz+NM8Z06eTexqv+tOX0Ae5BGtNRf7BrVP/y5RO08EXgq0SYjs6J+LKO/FcZw
V3Slimnfqm1gIs29/PvQX/bO0ZFpkQHOm5BlvE9AprK7XR4edIO2w5dw4hJyFBk+Y+KyS1s+1iCT
r1N4Iin3JZ+WHvEKE+L/Fl++8KOOkH50w8M6lXU1xvX7fJ+fA2ktrj/mYUZ/nOh9kVEkxS6Tyoe9
fTrldjtRsVUya4fQL0wkzLE/l39WGxMVBZ/so15RSGLjbOSy1Zzv6s1oN+sI3JiwKwYOkbTP1hZN
1ZECj+k4dT7Ee+qn5sfy/TtSNACTFMaolF5dUTmB0GDOwv/OmClXi/TNPDo2Mbzgzq/lGpXnfhq/
jQZVqj5kov74SBmErOI29hJfyQEqvqgpJRa8KvUyoox50jaMaqSdeAFC84OBOnjD4FG5UlJOiM8a
7katGlF+NLohoE25YON32q4aNdtIf9Dp0dO2+ZRgzUP4k0evQE2LB99EiUP1H33/KoS48HakZS5h
LS8FGzMStJ6t6kS1I1MmgI/T+o3MIx9+LLwVgEC6C+Oradk0GrB4ctGYOto5IsFkCYtvWKmkv91g
sVLSWq/rsysajYbcjgIgoVYQfKb54w3KymsizYkhBmpIc7qEJ3PyVX7MI6xP+jPMvtgOidXMzW77
o98qBkAbdFo9p6EG/RjvHftra0RBX6mUtXXMWh0bDAQlTJ3/BowcRQGFa/s+bG7mTiExpH1zZPY+
f1JdgpgWJBy/AZp7dLlIkvHruTURbLmc522Q8/XwIjep3uo1S8BhQs5V/foVHolHFu5g45berAsN
V2BYwsi3OxSnAEvJdt36d05GdxR6KaH37HdOha7XByum/1GGIhiOw+fH2fpEOrF/tLpxXOWQV0Rn
PVEn6+rTwpuw0g8au1cedwwJAOwBPwwFvPf517h2ENlqwSIUHuCgWCxW0FZUXsmSO6+6BRamLTpO
a8Xx+BVfqqDc5wdTGamIqxZwAGxuxy4m9Ws+lHtVlEX7YT2fk3XXkppt1mWr03sM9z02X493P/+t
nUgUXVMZIpy5+2nLPpji3n3uH3/nNudD4i6J9nQuHoHrC/RYq7qKLCOlCpL+i8fHEjDACKnPYvnn
c/yHiCFs6c/VM/Qt8Z/HJRiovjwxma/CN6sWx+MT1bNoMHJ4mhxVizbbmXp+qdJZgDnZK0i7CTRk
exaNtBq9Gm6FNxrwXgJusRS0aBXVXuZhvAubCO+MYeMU/HXGCKBYdywPgNSBZAkRmgKMZQHfFG1E
4ka2jezoPiInP2QAX7SUpW2VyLkIw1RI+0ElCQeQ08Gz5UfOGibZ7ZxLmFPx19KhTV2j88TXnsmA
JH8fQHwiLspYCjE/kPDQ4tmoJAj2iAEzeB0ho3zP3xpSj0wjc1L6ZASGPu2k8/kLakLLEA/xuZ2u
LDGrMoJFtatB+uiqRiKeMOGBLk00GoDpdO/5CF6kG8oqdOgWjFfTqh4gMlw7cSYICR6XXFlzBv3D
2qtD7o0WnvpnzwvMQ+6/5ixW76iA+ypT+qYZOG59/ZVmsOxdvZLAx50CUkq6K8/gZLs0VkW+Ji3a
ZF1AzeOJlWcn4oSlAux1+FnBB0ykotLJy5ePGCxzd3Odf9VC7F/kjHVcebkxWXWttfdCVTrm77lP
9ZhM7ogFofOtIPnpvxbZY3cTAhwc6AAmJq9ltG1rUxYHiblC01kvpuSfaQm7Or6kuC+5ms0f5A6Q
JejuiKvSPp4qkzmptE0dgNcwqIFbtIAPyLQnHrRfum53q0u4zlf99GrxEcNiv7Flt3IG//Pa+ii+
E+BLMdCFPsoMj7CRv5+iNL8WUxScyVewNxNFA3BFoqC6lDElCynfB6QIBkkOSfefq9FGc04jkcZ1
Brh7kSTLPfa+F0ExANIul6hWU6nSEgrQkmMtZG2jWswVMf73pyDZalbnFJ/p8/Sd093fXAggf959
u0fBQyjZnl9g84Y/nFS0547O5Or7q+lxION4qHmj9A9v5UNgCoFM+8Rj/VO7tekfz7qm2OBmokct
qpNoygOQ94chHaOiXNIP9GvuIrdRSEIdagvbMJM6clCs2ToX8QSgBsJCmAGXQAJA7WktOySrhQkw
1ZiwNM168o8dqms2SHQtrMyPdaaj5jP1luMYSU0enwiClqBVEHErXBw8SXgzSbViEqJEid9gAUPZ
TLrXUi/WjTlDlpCCPhIhlVUAt0QaKAzAH19OaXY803jW9okfD6VLLS83MBOPIwXgV2kR4QbdD7NT
UDLwM5dPmnMZRPJoYJimsBo+22CfovDiF8EgYop2tnp2V2A9fk9+bGaRB98g4Ygir6kUx7W0gB//
bLYYfq0idJoiiPTkGbPa8bjFmVde2FEC9QWPEKrYQ/hHBkj8x9cOuut2Cgh93JXVey5oeaVQxE7Y
G1CJkC43dlTSEHngJkq5tV+XCqJPirPXzCm8iunwA6Z6TYAAoVifLadOAjUKAlotsOISxTW74Rzd
7HXoKSgq54iu+wVcgXlUSqsFHoRAkzJYPMNVkT3c9N1KktxXK8Av3fVL6EDe9R3GgXkyCp94rkDm
8ypMm2sadVoKhfD76spxpStsfldsU74GYa1fxaUlSdq8bawUhWyd7fb4Jnkz9JNIleVraBG+39FJ
ZQ93k2ZdM1B7VYEEVyg2CUbsGDopZYWSFRrWfUj9EVuNj3quF5gZ2dhNMjH/dp9R9YEb7Hicxay3
sKwEEcX6btjrLgTl7VnSHd/su+8LCOmbMbqDwp8LZ6fyNkgXlTisyDgeBq5/ysbZ4Y/bm8V+T5Jf
bGDuoysErRn0oPgN0xc31ozXECuSQoojCmvnzPKtI+C/shJydkyKX4P3cTII/4cY0kSY5K4/uu05
SzVcgQmxdcFjuKsjfwgRTYGEyF1tunIB/pbnLa69t/KqNkaJyp6rh44Av/Pyce3PkFbQqXFuVt4J
7phhio2RX59EOv9nWErpYj1U9iKCRvDNnCiAF7HjjO+kVv/Ds+MRRSycVRFU7MLpmJ4468vIfOVK
tsJ8TYQC1Z4B/jGaVB2Q43c5q6/MBQ7OSJWv+GCEfYW+/2gTzJlJLtYDOJHMxU/SuzkK0s2fajAq
0o0DCDYRLhf79M2+RMpzKg/8WDxG6genGV3Qymx/EXsPudxfSGORgqQWfhMg9tcUF6983IOGp9U2
e79HIATiIPTmv1ClrxxykQgyLCVGrdURNUTAG9bb+qY6hgt7ooKfH9riITTnCHOc3Z2cv2SEPDoD
bFVWbnneisZ37zrCIBGrtEKI1MoDi4kAREkc7WBF9pev629WeFUJwjJNgNMk+zCIBL/vIwcqzqhP
CBtNw1GyMPrt6onMFiW1bMlLmp/DPR+PrPQrru64YDQpiSzNCsxfv4defnf2gUfwdh8HlWuFjjEg
f0bycfflyXYth9kF8jpZUY6xad858CpcKaoJ4tD48OkaFZ2xY6YFtlb5tv7CD2gja7qJOhCRwjXN
bHFc0cuKco2/bZstosds0p2J8xIH4efeN5fq/wTLn01BFbL6caYKbW2iKfY+PdL4PDQE4M0Gfo2l
5Tevk9rg8iAm0N2m47ApoD9NODrCPLZWJpuHDm1oJuwmroVs9tqSg7nEnXyaKYd9WUj3iA67QCqM
rjrIlionOJT+OYcqA45ihZ2wRJxojL6Irsy1hryrEZP8OvtVxhWZX19aYQdSoGZbHhHBlW0pTCCQ
xRt269yXFKNIW17BsM00RYIUDfY9wfYxfNK0VwjOAsURuTZIhrjpVQBVeSu5DWgPMAO3Kl/PmZTF
WPmu4xenR+fC/2lv0xNloG13RPqLCIXALJA4SUJ9bRfAmFAqaJF7I+0KbC4n9+TWjtF/mWLI9htP
FO9Ahh8SZV+SvbqYVACAoACLOOxuLYmjmBT0CEw4SXQCwT/IU3m3VgAC/GTG3lY6DxB5KMywtyeX
qQC3aR3HwW5mjjE4vbWX8tzHbdk/NbzyZitm+rf9oHz+HnsAv00pJh0S+JucxsFegaL+UywHBvCS
7uXDPt318ylRRsTxT2NL6s7q4hLwpp+YHKmRMFT3wGVHbXfwhmW4xEE2FPhL4viHbSQptPTUgqdm
YXmSsrxGWYSA1bLxsn5uiOZ9TKbS5QJpuvb3nQy3J3siKpBOAIkp9c/JclR46+5QDR0cllpcEukC
v0kzEqGugn7f2xXrqF1hnXx6HGyksE+SUVfYRgTIjAo8gjQQ9pvOysM+zYD9zxCqrOT1nZyOqxOg
1RZR3lzGBbDlaJ8SeRTSsoaa1Blv7RgIHbo0Y5VRtgJfJukErUno2r16oSM4Cp60uHMlWHFhkCkm
56/kc0AkFVYgOEOiu4apWtLLuSXycSNA1OsGb4+eNsDpGJAKIGqZaQCuufuD8DaxOh6QtZgC9Vk/
TFW2Kf+Z9fI6uE1xWCSsC9ExGYhCb5HL55FfAxFkxsMqI5+kh7j3RGEr3qg9pVQEGyQ+5CMfy6zJ
Jz4numP/QnMh9QGqTWGfg+J8fjv+dNcQMIqpQFBx2gR1EGoxc8ytd9mrhYm1L6EVez2fck9fhWtm
iwpLPTgpoDVYNZIaw1gjQup7MECeUxNF5hmYCi2jYAfH3qhvcqYlRdXrdHDGfUtohddwcK5CAkLb
E7q6mbZbQeWtJJLk/POkFpewpMhfe6YmgAPsgjgx9yv76fI39KHM5NyH3JT7QqqIZIjamsrFkBhJ
lkqEqFIeLyDjfIGsqlow5sdWugZJb3sQV/tF2cYR6L5UmT7pjeoy/p2yILax2LlSkpM84uio+6AF
yTXTQ+jtt3Gguon2Fuhxvl1MOJHT9QbovYbziAI6Xp5267l9/0nsvX2F49PnlLacFrQG6v1YoomB
14jyUw+0TapGuRVKxlSAMopxNZostd8WethlP11F/XXhVrtXf1wY09Fj8/DqACw5ERP5NvFMy3ZH
DElG67VvYQC6IBdQySAYnMdHvIBEujNTfJ+Kkz6CklEBB4E5HzfYJL2BY3IySTDkvTw9hz7DpgXf
el1oAi+ES7NtV8MwJoFtUt9aB1rUjDqMzIekftpoZn3oAawXXZPKtWnifrC/BDFKOMR288wUfXrL
kbq/xazLPUIgkvzcOhpApLFxuO8ba/6S0a/o2477eYhI5Ea7n8+l/rU2eK0wCEuRM0Blnx6aPg42
H964LYrbKEocMN9ZMmZ5az4cSD7KmypIYeuBkmZ0augA+U0w2GLq77fErQ56uX9JD2N6tuM+k4vs
bAwEgZ5+h8pJjnXsnJVUeaTgbk7/6qVxcudY8ebodElIVMsMmPnl3dZytD6rQUh7HZEaFGKk5LTg
7sYx5fAPcSbRJx8JNXC/f3iSeWqZBaBgascqE64N/NZ/PsiUqwlAo90f4/uJBb/6Z8yJPtR8kDmb
rmoIg+GzNGNZHVXhkpTssp6kbAUILFv7rw1v/JhE+dch6q+bFBGrrhdlB1jeO/i7q965qqfxKW0u
ShLk62bBQg+1xnTsU2xFAE/PLHXBbH2LOn3VPQACTpA1ERXKWISNZUXyYAupkx1r/9QGuja2453/
OveYr9IIyWqm0IVV9djHfmF1oDZdjmdRrNy2Ge282HwCc12pQd+ldGGIv6qcqHfVlRD/jtlivSZj
atrv4no7LMpBXoZ0/9ef/a4qLVLjDLW6oaRLYb7Y6ESH3UaiH3kuOrvJq4Ank4hUyyldoqY8LeoX
TLFXY8zxVnCINmfDeVyXoziCKK5j37w/vxC4iFmRMQkA+mom/1mAfeSJcaGmiq6YPCy32FmnyQrt
3Q/73JHd+jxHiYw687L9oDBR05lh5+DwUtOuv5JYFNE3oBfwgSbeiyCsyuhiyDbLRiN4BNlJNiiw
QIIET+kvxBt/kISWN8MaaqUUxa1xYWPk8Y1X2CQD4+dcUzax2fNfAuawJGUYZEhxH1Iy86Cx7Lmf
QAMmShDDVxZh4MLcVLOG45/K6zpO9UBlTcV+cNLZqxzsohhWPr8UUQPVhOEAdwDTrhHZkB9v8aOu
CO8fuUnZcZ6/lVBnIH0QUzG93SpCn1BH8vBrn5Pe8nPKKyWtzvSym1JEdkwgLZTX0bOBbb46DZmF
1nS/XHBIYsTDPi15jGCFnXBzurASMIc4ZuDeZgNvkU2fFZTm4PzpzwBr0DH7nR30AwSA68Q8YebX
SO9azV5SR6HYKYxjcJtK70XYTyIkFYfvzOmLrqL7YXx1+rlRTiZ7gC/X0kgewCIaNV4xn3nuAxBn
l8b64xo7ee7wrk9FSH4N+rfJlMyuto0w9WSRK39hQOjCvYQBD8jA1qTSdKKcyxYnoGIDoqxew0HW
MwgOeVmiW8uzGffnFcSk+DZy7SWNsTi/E2oCNxm6QcnDo1U70U1XeswA2wTlOGXVn0CbQK4rBXpq
gXZmsPuByRlYE3Qd3bvBS9MQAW9RxI1Jf+cgna/5hYLwXURawSJZNqEjhmeKr3PlD7ENDMyVha8/
MRBHF0pvlbhNpsH28yolmq2Xq8oYsxA1oEwn7z16XIxlHjT034KRARpCR2ooKu3YbRaF0hs7SiwN
FrDdPm/bO8qbFfYFN6bjAEiB6PShhOdFs269pl4DQkdOTgjlpHoylGIIJ6QrJJxvvEzIBA5sLl+l
1yOLkgq3N4DR7s7oWJ4O/YzO/SmaiK5R7lIFsA9oDzB8j6QfZ5//nETkz1N7ypJCdrpLO0Yzem1N
k/TJzOh3BVrKJnjpma19OwgUM/GB5bbV0T9JXjJq1Z+xtZQcplo/v82NhR5pU2eMEaDg1IZY9O+H
Glv8XakwC9vHk6nwKZVNNJyjO2wiiqZlmcaeJCmKCsUlMSy6XA9zYiLMc1IiM2s6+SqbTZevCWqb
9z5KrTxAla7Ziw+gv7wzbF/Fu0i2bP+KXXMlQYjgOhvEjiTtFhhYp+Mctd+8HppbWBTFPILJp+4S
clMtftCMU+xjsALQ1ZC6+a0oGGzlYJ9X0kk4AdAr2p8cfLAymYPG42VydwAxN67lGmYXQ0OWN4j2
zAwoImUc3oQVEpLK5R+ueIiAbHFRvPLJK4mM/jBlN1hCVQ+H0sktbr3s9Copn27c/U+jgIEPyzu5
dHvuzTvwWliFmC9PJHUaAOX1GQats+3pP6GW4f/Y8uTx5ytcN2sdMYZYhbn+x5zaycSzOIgECm2V
cQr/18wKrd+hOTzCLIp9X7G5+IBfxh2e33VRbeGHq6GLv+ZQ0yGyc8pYg4NEkh9fw7rQ4dU53/SE
dOyTHabEbadx2jPcnAM2AWvjCl1mGpFZEct6NwlwB+vfS2lx2xUaoTYhaEEYZzhDnxGeUH863Ir3
MHIWaRYk9Uxl3ICMXLgk9bhaQANcMEzEi65iTdAbiG/PeVmuhLM4jYToyMgqrBUaaduUZc926hwl
dDHa43qL+Ut59c3IDHi6ikxl5k0YqoYVSuPnjhBIPq4aRRTXPIT1cDDgQmpcAywNstolC/WTHc6I
UbEiDGx2knz46lJxvo/DsP2c3mViBJuSUZ+6ml4au/VHFgJYrVA9k8PooaBUqSIo/a/aadaRrZ/h
8ceDEHQ82M6I5K2kmlxRnwupunmDlqKYzJbWJFpOGqg+XcUxjwQWjM1Vra5KU7+K/X6kJF/G2Bwz
UWqVMElKZ1e5fSCO7yNCn9H6q+DY+SzIoFI33DsGPnyHzhHWW4QY7y3GPB1JdLUffBL0rN1L90Wn
T1Q1+UPjEBx7R/HX1qBpl5KDiRWUwrmej4OOY6KwVO6nhpxzm7qlmS2rjNVU5+HhDAPGNZNF0S9W
P3DCmBtjwGT542377CZuyUwvXGCnPOnDzbIcWP/fnEFY7JPKaKpaw7BD5BIF/Mg4V1lRGnZviJJ8
BL73cq9iM/70ec1EmN0Ke29UmU2n9GNl8tAK2bfWHfVBQT+rFkZ3gx6rJTwrZMMyGPRCFtR3tDdN
CaokZyObkytKYGKPKC+BJB5o9lEDnH5lctL6O3Ei+AoQbiB7gNe2nX0aLoKYPPBDYa+tWTU7Dmsf
DsNMSPmW0bknMZmRyOndpwFE6cIsZscoJ9qiuqFNIAwtOWeRy5Kxbb2TR3sseHHrQKL58b31TbCV
eFtiYF9kJZOufzDrdolez6AUNtHr8FK2I5X5vgskIuRSJkxgNbW+QmxDoxRYkq5o5Z252O3dXlXX
Sz20cZroLZzeAWz5Vo+2gvxNbWp0+PU6xsAxmYeNjRFZguqmXAdKJKfe/bt4A2zOU+8x/t6VlUNd
0KBDyo88LCQVAH3IUde3JzyOrthCWt9pWi5pr0kCJigmRX5w9KiJeKGYa8RyDcwCvyWeCjDFpnIm
bijR8qVG6XlsyrJYQW+fB80NqaVnZb8g+/dPodx4gd20XO1yWhk0FcBPFaFfF+aFLpnkzepTALib
PMH2gkMmu1E/khBxvcjj+WNLAt/aJ2GJQ+6fJTc01Fd5Ec8rdwKbhkiD8kBIWP84xrN9IT2/XkiL
dn/ZKiAWWTtSGZj/0rLZQPVQntkfzLwbHMoa5GRoeEwN4y4lo5+hKK5OIDyRAR15Sy8cZhCtZhRn
wDKpzvyN1Dv9bt9RulRMlR3umNunddpbf+oeiLf4kEUBoQRkEhmEC5wpAyPf5ryhd++C04KohsBW
vy0h23MUaRpmc3sLhRyYwnL72kBbbn9ziCOgTD/1/Xtdv2fa4hCxGRJQdUq3d8WgsJ9X6vK6YRvh
1FUx0U7ZKN031Qi1J+inSrf1k9DuJpvIjc3t/zs/j2e3gg+zWrMJpz4RLRpkie/XAm0P0ARxEbz0
lLP8T3QcVJtKfjUI3sjitAnTVdfHHfwJnzzvZ/MvhvzaEnegdewMtNj/HIcaUG2NyXZbedW93XGV
gixni4WwDGs7SSxtAJt3PQAQMdaFd3CtCjF7xOubR47985YPf1r38Trxr0HDn+IbXES63V1PoSPV
dlTagyJu1/uGWrxChcMz8WxIsEtIArLo61ZvCYaUJQSvx4WRHo4EvwrHr3lQbA/pLvZU5WyxID59
zqbE5BmnT8gJz347cHk5kK2CVFJDNeHEsLTveLPYV5pMR6nhqQZVod+iCDRjGDhkDZJbjBDkHJyl
8EpyeyaKXhXWlUWHxNu6msKUkzlWVpoW3CLTTQZhOkIYtpK0Poh+/tbw6CjQ7ypaMwuLRAvxJDXS
T4H1yYWyUudg8TxT4Mxhpt25PrnRVeC+oDQSto5VXprqlJ0cyHbroiXGA8fMkc8UP1GSpwtaDKFY
NrXXRky+62ciZnylMx3ob71thZyFSKE8ZMlvqZoV3JJMq5+PceDlB1fzhIVtwzOqmxFZKa3Yag4L
75Vn59B2qQbR3SukmlRP8lh5ZuW+Z4OlyeXpkFu7T8UDwPiqCK4s5K4UKdsmAoR8Pr3RgHZ+xFRq
3fWJ+qUeRxHkHtl87JsTcS4v5wy2y8oCU2XzdHgla8SQDrLgP1t7sR6lLKZbiFIstBEST4Q+rrdO
rjQNdgjmlP74dhRLwIwUFfFOXwWqGxHViTHlq43sERgBQ6DmIya27kfYyDqeTEAWoyEjKvwgm6ce
TjZuvYHBnm1Nks1Nux8Ip2iaiI0lmm+rJIzGKLSzkCiLWuGHsPvQFyAXT/q6rQTfYMhgzRFDuOEO
tpLP+3TA0pdmUbX58suk1WUl+T+jQOw3LYr3re0Jjn1ogN8G0MZjZYmAYoo1odhru7AdE68GU5LW
Dfk3fZLBblGIb/+mk3wMb6Pqm9+3c7eJ6w3FcrRVDqs/0B1vkCyFdumdqX5JVyWqZvzw0BSlBlKj
mYCPy2V1hnIuVTzUiZYy0i2do1LIDB05jD2iefRDLxNo7fExJ2ozQqH7+iW1sbi8Nl8J3YyWymae
fNuyJnRKJUAHWNmiyZRruE1BnjH/dhSCyMrHX5MartkXyg7Pp9WAI44EKF2rBxMCGaccIE4yFyBd
O8h9Ik/4pYHzj3kyFeR77yHt+bdr4mVPp0xYPpPev2qTWqyFJqqbkKrk23KMQvEQOEYm2pbRyKsQ
5cHERxdr50BLoDA/V6I0yoi28K3bRiKmWeCjM/EqklVA3PXcI8FeloSAhWAupzTbgaRZCyGtmM+J
/zWuMW4cZaFKovoo0qKsWAl3DLFWAhqUHL5xyIcx9AI5Z07tGrUWYk/Wgc8NdFRc/ImOFNbrLPur
uFABOUGpZbs+svYKQrrLehbsSJ3TYGIlkvKEerCB1JzNaOld7LL020Cn1J8pj6EF+2GAi4CIPpVM
twHrtUzolk3IYLb0/1vDqadRv0TzpWYEorsYb4aiB90yMk1iQohPlnB3ryYIQpPYSH3Ntu3JHTLJ
AnPWUdOe/iuQmiXKBNdtsQ+l50ko9UoV0VlKbo2LCWwBHLJA622oFCd+lLXWIkmmxTgdiJQ4c4xt
l2nuaJf4HTBCHELMmpqiu7EZtdxUEUQbg6xvYDGU+aR8QClaf+2Lboyy7U9qumo8Zg5r0ae/uMpI
ILnwBkgOIHLBOYyGMmUDobXp9j0Dc8DPMuR2QNIV+H1zTFpSw5rqq2btSvfMabtsk6z6sI5BciWZ
fdGrKx3P6+HtyEJQq4TuN1HR6vq0NPNwzikxNtoLNUd3/yun03lRNYeVTpmLuGBjcslmYxBcoS8+
hRUhInDZXez7lJKzdKFJ11mw2DNdDOhDJZEe+epalv2YsFE5A1+cWWUrghJyAawIc0VOFoUpLOYy
p9f29+HMZa8CGRppIPFf4zAoj+fNyBqgoV3zBLFdhHmo2waXagF+l4JtIUoonw6/bUc9PbIhLYJq
XwNPo9ysnMvSZPvkx8YFuyH8h2rYBbh9ICc/KTLKHGzKHiPIwHzcocSdZSbRX3CL5EP5SOGsnYSl
VRkBkwbFCjvuXYBmuRIUJvtY4vu6U+VFACAZSA9dBZRR8F2dR4/SzwF2qAKtZmGBOffbn2bSkymI
7vHRDGmzdeZgKWGlcQ0A4abvrBCaONfmTLTgHCFfSX3RR2d4FKOAOq5IuUUKsfEZo10/2kRkGDdf
sQ4B8EN5I7nqqCxVfYeP2rr7ucxZ/us5xYqkpXIAVvCwXjY55jfF+CcgSGYRO1meiCw+ovcV5oYY
lOaODZHjaqjzyCoslzCpGBqDc/FMISXWYcSZbXLzGX8rnXc0yVPG7OWVlzqudAcewCEesEAAea5u
sQ/jOYDPy4FbVVHwEbU51olIBQUHuyTVp661GmM/xQF/9+bsvPmIMeSPhY3vmyxlbQz+WPWoOSqK
AP4DPx3f8cIgP0sPm7lmnr+BZxfBDk4c2MjJz2753LWSz2ZJHpGhaXS/ormL8xwGqepJaDRNTPt0
rjtxfp+raBcaZRUIDaQL17etY+vvhLisloiL2RL/5kpd/BcNT/lOK4V1x4cEFilmHh/Y/T/qG/ti
tSahmZX4rbQjrkp0uz9uc5eZChMWKADBQTtvpF0MHjGY7fQ6xXxX2PsR4O+ym/m+YQNFoKlX32us
YUrkyjllMjTuJtekCNycOD8nGc1qftlsshz03P7jSC5qFcYFr7h9XtfomTLXdO5ztqrOozfPTTPY
npdu+WX36isnIyj6Hscd3CsD4fcXScspqeuFQt65mux2wqEIqxuooWbKnptDfkHih+etczFDpQaK
8+pAXVjp2mw0UhUjUhOZ9hO7nutXVv1T0JJkNNfVzbcRCigRAiDFJvy270OW29v1Xs416eJoXtWg
I+vsvvOVxTBtPdjawXuOtgjuZmOQwcM0KAqvrrMZNCMsZmQMOwToLgtgyR4MBG1u0t3YoKb5eWf+
t2GKCB/eN1oPEgG0GD/V8rPWf36goFAmSoo6KP99mfNC194cDeoWMOBMGzvCm9BbrAITmWQkWGCs
JnVZsR+PtATt8vq0zeirdMaCxOlkKI4o+IJJwTrBllf+DYqosf5A29iobURzfethAEikJGGNWmB4
ZahvZjb76LcTX65HT0O7FMCHv8xjCre2QbNX7gXERuYs5CrFVN4AjUV/BICUhgMNFENTzK/e4xFK
vfAu5MAKjpqbqHzefI6f+9O1EDsgp5qnHa2pEPLiPy1vqtrgDGhxk3PULcD0biGWPJtH9SZPjEii
HKzDq7zsXVLEK4GEOBcRYPoB9WlFAm+MrZTtFszRF6S39KP1RGVnYllcrIxgKiVK2f8zVNXQMY6Q
67CSmWaY+UXRKM8ew71qS8Cj8aGJmdJPPTFdOSWe6KOw6gtQ1f6wCJq8SY5dL+NSn3tK+I2fbebF
j4eeG2igWUILvZA8l1wPqyizLhUbFjdGYM4QtdOIX2jvSD6GeENyhxOmrufgPgKaA9UKWH2Lyhde
X+6sjgHU+3cT+57J1r+LuFYetNpORveL0DIZRTHmkXy/YMvMRIDZYq1mBhrvBh3zxB+No4Hie2Dg
Um/om9juZ9x52xL/WvfuaLNwvqKtl0rjwHJIVu09FxvcB4pYJUFF6B6VnEP1ZKt0XpnWPuSXg2YG
oP0NA8r2XqFnWvMTXij3Lxu2wWjqdi/P96J5wV0xoqoulH42KechkMRa0ehXo1SU++wAIqtZ67Pf
dNyGURT/miIpQ/KCRAo6bgORTlsMWkMXYas24PVDcWBjOMo3THQ2/m85Es8P9aWxGfAcuKnbayQS
wU9wLAVUPFN5heTyvoDdjg8TuLDThkQblyJtzxPptJi5J2TYe8xt+Prc/2Wde3P/bJyFIDRzZ46a
056AO17Ey/cBIcLrqdJwJ1ofbDlG1wOkG9N+lPvAR+6nFhh3Urrb11urogiXzUGNXf7RVILqtStJ
Gxn2TKtcXFzNFJEvhHAQqA3Ohrv7AcrZiofaL2JUchtGph19Xoh0rEu1XNbz/1S7fla4zDjuH+qi
LQH5I/uMEb62vxZWxEiYZvtTmmUjpknurzmHgLg2wt1va6zkl2/mUGN2bau7Q2V5oeVuKC+tGKpN
QS1d4OdJxu4iWq2OSoePUSfvk3EZd7/3EvHzgJTg9PPbJTxbnd/HeheWUOd4g7nqgrcYdZxkFtup
ea4s9tK7F/SOvTBZE3h3e6wJoT98CPTMofWiQGWkelhclahzWQt5beNxrhigUkmVBxQzg+Trgt69
svvvf9LWSRz13V84zMA3f1lIVTohBQN3IPgrvAlcVQZrvN2KeRlKBYTvtQzGAaI22fjZLEcQ+rrD
6PEs1JIoI0yTlaXJxHSRO18nqDfKuvZ9/GtCBwcOm1D7EBIYOzDwmVHN+BMYwm0nllJHjN+hpznq
o0R3lt7r0hWKaF6u0vVGKsr8t+WNz4yjbeRIqO36wyRVyiN6gKBywAmOe5DFFhb0rF+1AtwKGGhT
zpbPbvernM/YYqcBGehqQrEIs7FM4WqZbtSx6JihK+Vn27dp+vgzrznymbz/k7f8RNdxZLu/MZo5
rEPtiBjVSj/raCaxg2fzzzPEDhDCeMg7D7Hmf69gl3WN+r0IIg84emGrf8rsCcos1QB2HxxFLle1
nW6OMMVX8INCKhjOev+t15Q4B3oz3bqOnjBE523CZctBGkkRaQPeM7IyH1vMyIJ+NdXcU9PEisgq
Bm9me6J7HRhUZ31mHfaSwPFMqJ7vbVafJcABby/4mWmj8iyaTW5BzDC6m8XzPY+pnuMjBzZ30OHg
iCx8h6ZSRbV0tIzqwBPJloi+j8fHOJxz7tDXc18hT+5cVkSVuZRO5poGFXtwH4GAgkPs7Jhfvtwt
G1U0ILekrdckpw7W/D5RcbAJ+qx7xINaHdXghc4xzZA9FWzhEQdsJpbrjCLmyRnnwwzMAk1FSI59
KQJ8rtWGWRxRwd+m65XIjN2Y9G4lceyMoIYUGzqC6Tyu+jhAuTDm02FvLolCe2oFDNra2wXS5l7q
LMgduJu/Q8kN9k6BgG7P8rYCw9DRG9i/DLDm0CINPqqiQV8TI5hypmfSgSyLHaVToJZuPRASkXbd
S4ZZRunhSTIpbfY7mqamcYC+jyoEPhZEcsY98DRR62uY8Por6QhCVMZlyX5xdYH82ogDfsvL7MQJ
wyHNdYkd/AmEVf5zIutmnSrR0duSFMwPKlhKDL28JINxI2T8TzDDsR/zzfgmlGGmqRMdWZ6OmhV1
baxI4DaDhFHofAMczov3hU5WrKqzUuZ+pmA6GT6a/LzfM+F5X8yVJKYgIkdbwdV3C3IT8WfWbgxB
hDAt615BAfUDhZc0Atd0SHYBTRAjaWLgLEG65n9V9UtdqFbH6+B7qQJCgHwWsekslfcjN3qE/i52
SMygETT1+G9a+jFl84eugiOom5iA8QbEtPlfq5jSDnjyiBUGhawMEhEiRptnmoQAqKQ/CsC18MbC
LhCSy5awx4CoIZs/vvY5ELBkEr2dT3B5BR/qn9sDKUXPpHV+AV4VXdTXj9vRQUyDzNvQ55cfR5Sn
OsrRTz/fOIZeM37IQcOgpV18Zyz5WnqH4mqxrelbvLwPMsgDt9nh8C27m3rxuMtzHmnO0a+2DBM/
C1jYgz4T38xRnoq8foYax+FkvBtyMdmdhY39WABBBOGDPmPVRX3FdMO+hOmlpAw2k+A5sXaQ0n6Z
N780nrfTsMeEZospSdhYNIsKJ4Q9Hi2rNOOkK/fjolIcg7YAF97/aU6Vh1kPeyP1scB8fQatogOd
++mFPEq5D6LoGC1czARD2Tjb7LGCTVPKMtoKhDRYbV/XgZSCKv6ulv8F+3daY40ZcQ2K5XmHIZI5
OYFc1pVcHJ45yLPmt8BrnA/ktGmV2BZg0NE0pXdhMQYDapZ7njGaM7u8VUW0LsBOJX/+mGuWl6Ir
bFF/qulohORWTWyY0tCcHJ7wlwW+CzaB2vofVA8WSH0XYcpbWSvVMOVrQ3ev21iK+5S3KEIolcSV
3hZ4fxt5Imp3RtMATWMew+qhmEJ0I/UxA9vQ9SOlrMrs54nSYoSbsuk289ZGCKHpV4c6e2I3DtRU
wEUZEoQnklUYHcokNIPClQ5I+yltfSUJT06r+hmBkU9qHVivFYr6AGP9GyrUUdvGvoElUoF09U8Y
z3LJcoJyJcY3T8PFFTWCim+gisDkjJrCCI6muz8WP3EhD6QprCUqlkN9MEp4h23DIDTv07ajiKoR
tDo8To3GdiETYjnhjqakC6VlxwSxErSESf2fOI7euwLDO6qSTYYo1HnMLGy4burCMMpLgMy0DKKl
EOOtl0rM1ykRSB4dM4yzvkO9ypYLDHp8Xm5BfP+iFsqMQHSTV0FWxNiPcMCY5aTHJf9bTks+8zqH
Vy1JKOiYs+OuZkX87UIWtyAojt3r9pZc1MtvJ5b84PNRmOMRpf10oqUxMsRFHq/F8VzU/eJ9rGaE
dMtZHOokWi321DARuj/2PHfXIMFpHgvePuxgNoTM9hSR3WN0lFF4iiF51/WmdRMq2IVXKBauHbuJ
2CQEVlpZ5hG+aUwTYDT9Ynme7/sh0Vm5orUYUbd69a5GDdsYGspryGz8LPDjfxu7zkTDB7Qp5tG9
sg88jOnx5PlfZvjF/2K4cNAcmx+3hDtDSRZ4Rf/GnTGfOhwz0w6LstF79SPE7Ox6ZnJ84QxZqn0W
+6/oSmPOMxLuTUJ9HRnv72nCB615Dy/J1na/EFR7agvm7aAtmlctD0zFUemwQf0cfUDZVeXm7M37
8FEez2+mIpBM3xe74ODDRNPeclf4vOl1tPCo3x89Tjg3Y2iSzAotu5Q3HE3UCKUPHchphPU0JHJV
EjEIqDJ5PtW5yhubALvfuehj9B9WJyI7PtJ59UVvtcFI3I9fmHCCJEsEzI5Xlz0+jnJf/qB83RV5
Mhtj6HoXDVUr4NE7sJqH4qxmn6mPixP5t38zAXGs8aMnwbAV8vcY+A/nBeeqvtfFvo3/uoAFZzYY
yheRzLQps9/3aqkFkU1h85wC0hTn8qlg7BKuwfsmxyq5jKEQeoydn7D6IRrRn4ukrGJ923NKMJ5e
tBinuThv7PvC5fgr7faKoVPbAYp9lIy4eY0kCG4CcutY5X1zZ9k2MhIo96xG28YDvTUaW3ZnrpXG
zJD9MMnQnieiVUprm/DOeeHC+Q58wKzocI4RPPs/CGGi9HnN+AsFnTFUJzUyqmiyq0MDLZ+sWcIQ
sJjiVUe54ewxx7wQnBytUtbA4jjKa+zsEAsVHxdyVJnb1ADSLKhFnuEI+M+M4IWthpg0LqBFOhaS
382CXQy3ajk949/OSSplEWmGMhkRtPgRG+FIo5xrkqd3VmF4QT7SW0PIOSBNG2Ny0qBhKNJL+YCA
JrK76j3uHUJOYe8z8Wt6zKa4m9loEIB3LLbCBTHSrwTEdzbvqNUXEnxxU9GHWR+djKZi6uADTRS5
gYR8r7Md8CML11opn9FkXG5s4PN+CVKZeVY8ysjbw9Q0j0t/CX8W+dcpIQHPIM+2VRCAej3vGubh
OvNndFsbJyCYbh25v+IzZuOtG0hKLZvhzS/6wbggxrVSezQaRZq3qTL7ZV1A49M8hXzx6p3PeMuB
EGDScqnlieT3fikHsSaif/He+XQeldNqtbx5T/oon64i2AAmf0vxI84bJ7VuoszfTSQNijQx4XwR
tQ314zeEESVxgYq5tDENKDXtbc7zq5diU4Y7flmBpiuVJbZ1SV0H5eKs1o2KWiEz0Glu98O4M5d7
mgP6TtSGFer+nw5aMeYVaQi2JH6V4pP2oMYaQ7BTq5qB6KdCE8grmhFfF2HS3dk8K8wYyDuVqOyZ
q75lecxVD9obqczuBMmaA5uBAn/kVBOc2SPGrv9ixMCm2t6owjcjMdbCBh8AKoKq4RCEFKId8UL4
rMrbhuMdkMVyzrF3/RcvnDadPsIDS6MVPKi3X6qwZ+L+PyaVH/muH3S0B8cbXOPMluzAlqDfzoji
YVrtolIgSEeWBZsh8hpWcSIjvSseYryJMEr78Z43mN6VvmvAtYd3LEAyxh0yYoVt9wuAM3WyreyI
n8yqPcrpiPzJPdXxN7XC8Rr+sCIzCt9qkNFU5oCbwxDJFfxqPaCxlBl5lm103NgoxE08Nt2a/cOs
8d2oEhgaGVeDVcdVkrEIUIGCqlzVZaNTdZ71oFcfVmb89aFFR/jDjjcsX3vq0Okv1YNJqFeTC2Vj
rHSeyZYBB7tRkqf+H9ZD3n9tVkh52CJA51wPyhk0+j0mmXQ7n8cpHfhIZtmZg3UmrcjVnqp9GWqS
w3AVsXQDvdSAWFl/5MA7QQ+aBIb0nmDVKbOu5rDA0tsjA9cXZcW6CYohQ0HNUwMJaKdMuz1QPA2V
lePxa81E+TyrNIHPDh2uPzJdCHt6TGLXEJS9e/poeRf7OOZpiHK1U63tYi+XqkesIp+/CZj81Gxc
ChZD8ZsQch+cR+Rq6qFw/jdARJBwn5Gka8O2MDYAMHQSevFvbEAOTho+LWjLiq5o6ETlAnIB8NrA
yf7l0FcMiaJ+91xVFK3fWdVHr8ww4iDRFqxlbNB/PGo4v00Fx55U0eqgIwMYYOLY1cWiRpnlwhxb
CRX9YHX3b8apDo4CClpBaiM0iPzWkQ8zroEvQZttAkt7y9n6SNYfo0ay8b8mM9fbVkNC1v6otTHZ
2HF6FXlRNlXfETfN6jVDZD2hXJ+w6YzaoDvPuLIIY6qnap2RTRVAorEOi5bQwAcSSgR8cMmzOEex
QpYMSx3asLnqauhKTsJEtDXnqwIsnXcXzuC3N1BUvHn/hAiYn/8XCEulVxCVvTIudn/e9iLa4j3/
FNtm1uK+3TN7p4Ej7WByhZg0PTJlsCZWhP9lRAFymPVE2keupVc3t8drHfU31dIUeyb8/X9NSWkb
31Nuaihsjtdtnh3BD78bl9LBaK6CQEJxL1WZjE1AfFTEDWDwwbUYxqYvwRrtMx5m5wx6hoU2ZJNK
N1mm7wPSFaddh5QcKYJA3tduq7kychFp5EkSHoCBWYsgmU699rtVPiiacQ6GLSoL2QrMpm4twbN6
t05e150O3U1xxS2FKb0xJYMLDI0ahJap4qbUFKN2MiTFD8ZGMwVuX4G8xU4ExFgNWdV/WkDCNVZY
PvU4Hv3J2UBlw2oMy4JYVfC2XBUsaVqvq35l2q+8pBxjEtM9zxaQyAYavO/3bT/gd5UD3gpfdeSz
ZBnaWKB5iOKnZ0qSKhFgF1HUHJj/59SjG6lUuDOfa80RStdXtL0ekZ9BRYOtQnxzCiccUg6i0K56
s9bJ8MY0aJN4mv7bd/PYFNAhH51eJDHEwIgv6CCBYeCbPktiWy0o9ndWsCYRHk20HYX7LQmdTqlC
rmuvNNz0u/0OyzqPsUuEocIaFigYxi9wGqTKtMbQj/HOGAbZvyJafGijoM2Z4ClXtyoAJYUUw8mz
uIb2F0hvM2HHOGZKIbKK3YnBwJHwOYBAk6pO+9dYisrvbHvF8zV8sI0EQ7Ao9/ZlWVIwFysbRDEX
oN0ldid6DVxuDfxgxTtrEQFBptWdZGO6fZXIWjC83L/Jj7nSWShW9ak3HTFBzqIYiYtD9onsppzB
5ZClRqEZamfydLgtzWAOKqGOxoGqrFcHUlDl4GPknUwYyhlz4G/dlZAVAq1VeCZOPCdjIQy7q7Oz
FPcmYvf4KK3dRSQ3oJplsZMvvyv8tQwTM5FwskkCDpNIIsdD2k3CMLAqs/MNIPW/q0MxZyQ4c8fC
Z5rBXL+5fHUdHHr7aEovrzFW8F1Tm1ybg7woX3OePrK5yPuylV9rbWcvb1Kcb2W5GhW2yO7PuoXE
qgx8XjpWWCQIqtMNgjMC9OwVImuAbb1+HMaCQ/mBCNkeuxH0wFmQsmvJoFl811A49oQ6clnvvF5H
3wAhpGCUtFvccomz+XxF1YKJrkkY1U5HDMb2wUluSnyiYt6+0ABg8OzuJb7wFxHRv1I9EceywuNw
IMklrmM9JJfPsBA5QwRFuhQJ3/+dMwL32Ozo/xJyC93F7nemuGxW0s3YwnXdZb2ILP7Knqh4eRsZ
Tz51LIgVLIGLOeLrr+J70PzVsTwLnq8qi2ruUlapbRNtjgHYPYPKXnGnOxxGv3xoDksllmiZMsMT
kH0BnMUVjXLh7xU6B9iXTZ+NWrxzFrFW3dNjgMX82qC3TsvnjneoukL9s+gZ3LHy7D83LRYVakfS
XZG5Px3ckjls56F2dp9Z6kHUlpUjoWrESqv6kKTzD4ewFrwgawiYsgwtrjEx1i8TsYYhK0zlNXXc
YBGT9dN9tcLNx1wj9bt/7wbxISaVQEifRNW1LvPpXDbRioptCAKFF+CLl7XU0dhtJ1lPEJXQenkj
UUav3VbIoj+IKPn4eFMwjrajO/fDNkNKv1lvYaKpx3eeWX/I++iZpyasmElR0eKN4rq562bf/+PT
fu2XW23Vj8IWmRW7LBY93vgRtVYjV5sSO4AfD67xrcVRVFnS5tOb0OImEsKr5/FYw7h/SxNBB0aM
aLnB6bMXRmQhIyXSE4l6dBPf8FTRg39DuYFrKX7GjgnrS0i0oN65OW5zPLdiXZlRvUgyW9TgbBZu
gF4Ni66rnE3WzDnXJxdR10yRfhAHCDXA4Wo6xeVCMaxvxLZV5t1CQlLZqmgon1TxuYy19DY/llEp
8Ns6P/TfjBS5ytuKQOLdFXOTkpvIkmiosl/7lpLFvpw+O7OQDcXtgF/7kW2jruaRL6tCRvgIymik
zYQeETpw+Rp8kqMo5Womw8hg+b2U2Os3pHLhsfiG05IvNHJeAUK65ul7lSiCFdT2qfQpzOnzcfbm
C9cadzB50920bdInbt18tp6caS1hb/8NSHeupgh+DxOF5czEkKqMdM8Btv+wf3asw9g0v+NHoqmB
QpoeGcB3+FzRYzlpD7v8G2hw3n1g0vAGKU54iT05LBsb9UafgLnM2IRCX6DUh4egnDkoQ6Q1iDeN
FC+vL2HgI9J5TTS6+bhFXTbj7hjv9Ez7glYWHJgHdN8yOi68UdqDoiWGCn8cjQ9NoSZrz/FfWlI8
QtS2MPXURmNreDC+lypDN42Xi38k6fo445qt4C6q5wM1c87UVmFa6SLgDjNov70qwmdIf6JXQNc/
W5K1R6B6g27te/fkEzbO9NK40nL3zcUtNwGkgCuIyW16POeaNzDWnNV2NXIge/IA9tkgXLa473SY
xv37Y91UCTbOPhs5VXKyKeUGa9Ek16wJcSfaGx6MttrchHM01eKdQTuvfCHrrt9TioeDyXubyw6C
dMiNvhF1lSTz/7hgP61dZMzE+4wCe1g1EDcMNrxH7Me0tqxhJDtCL9OYCC0sk+XrJ+LuleAMx5FT
bvk/0BVWqyIWz7+j0abHOiSElLozilhtNBmt9eOAumtqU/lUh+UjsDVsIE/JBPVy197h2AoxPh8Q
CB8H4uxiCvEq4ahCUcgLvMWgqPwFilByUBVM6hwV1PnGHzUjqPuV4/H503vc2Vuj1V+rSlST7GXj
b1sXHYMpcfFWRaql70luaHj/fmnfHcp+C+i1mbaA6AwxpBzzU2QwFYRSIIK9koJ3VlvhylvQSi4m
htnIlSOuXcE5srz8pESkePwpS+2ThNsRR1QttJPjCOBceAhaM3GXpp4ZIn3PGDKZdxh2BrdTuFl9
dO4jpw085Xdy4QSE8BM0+L6aotvOS2SjBkDr3ay3uanhgemlKc2Y3t6UU5VjPtCPZF6qQDz116D5
rxxGf8twpujTb/QlZIWl+WD01b//37yJY9GJ1h5HUUvBDpV2dlOQQ3eBEeEBXeHaM/GocOdrwMGg
6x3Bmwo0CtDeb685C7QurMIInz/YrbG+4d4AlgdRdpFtBGyA/U0hnjisBOMX6iQuPl3Fr/ZqvtYu
K8OjMdmsbFyNId5bU0MKR+1okfP1Fcya/gtFez9LoIWpEgUY5scHrOE5sSZ2eTLbfWS9UB4+uWYB
fR115KOpz2KTkG3fO/lwdO6n8GWV7WucGYLyLdOWRG/MkxCdAgTo+15y3eoukj13QKw+Ai91FJNC
w5+AdtZYYmV6XSm22OcugRFtQLv2iQkkU2HpPNO1Bq8VrMLuR3G4qqYeCUuDLD4N8vV8/7ywX1ko
bcdz98Rq9LZdh5hOthK5cQQ98Pn+ye68oZ4U0WVVZUye7HRbNh7J8gM330fxHgb8vi/H2Ped7Bvi
Rm15I8ULEAxCzwzMK10kqcPoFZYz+tjPIqzpRR6S8Cx9VHNldoJrZPvRERbeSlL2JP7wG0EkVP+g
wpYJToh8JtWjT3uCgwrTsAqBFWvaoMzgq6CwHVnj3OtkiOrFA6YRDYPsmwNwGfHhUsWiJVH5wsoJ
BRw1FEUUPx8SjTTnyXmom2LYQ48g8Emek9KJoVBmg52sPC4NHIdr5Ao0n4F4kQoWrtc/hoi5kwOd
H5T1fETZWFh+0UT5RV5UsEaFQufiHk+PDuIt2KCPd9APsodiVo/N9pnBR+EJAck5PO/lX3F/zNi6
0vURaPd14jE4kh6z4J5p6BtOw4C2pfubhOmWMksXJFkWpmRA9JSJ4biJsajvBEGQ2DrSFxwDHy4y
7tsIjcN+3HzmcgRU+SO5y+hRqkAvoPxcHScCKLhVn1nI+ITKpLlsCeKo4X8Jlt87nQtLron3I2IK
2W12hKteK5dSSYj/z3WgWV2ncYCj7Ioo6b2BBp0CkIsmZY9HtFSZG4h3RjMazDmsz5dyuW+6tLqI
X2lLHIaGcvxyFFZ2YgpGALfgTD8bNEE1m1DzGBjArgmnu+2E4ExDBamw8haEzTRnTGviM1pA5R68
gRRg+f36PrnNzTwseTBXD6TSX0Z+8lJQ5X0vFgZE52wXbbUaIsx+4VWbO9tfYCUgrnctoxuZtR2w
DyfelWCb4A/J3JudfDdWZri5HY4aZ5WDJQDqbaj5Z5VKDhUdDEoOR//NqRF6/Ec/SqXNHYbTvFoo
k3CWZICksY/JeAIwr68jg1gjDt1yFE8ouPCT3Gs1zq/cZApHBAuC2XbYn11+fZ1RvBgemGeTaF/O
CLoWg7HBscOy8hS5YHiSB7ELrTh7/dVKcMTZiG7jySzsG1Na1Q79EJ8MRbp/tq68g4AoHNKvt9Gg
uez+dbQHGiUY8kTyOEPjzj+nSV/ERB/m3nGNSWPB9nvyllmmICfxN81/4RLlWB4yRrdHwnsOTW9R
P+W11KEpPb4/eRZTr9AIE0PxgwHTkWX6XTsAsg1D4cHbz+J46e4/SyIkYw+vubLq+hU8tp7pMdz3
dozTCAtKjwfousH8cQJtjFJNPrmI6I2Sh3mpBb/otp//Ey+9J4mP7bKP9RWAFzPfKgjPLsPXsyDF
nxBNeRS5+YQ3CIdMt2XV37LBRhVe6DwcTxfoQCtAQ8J705MRhJNvd6iyvKfG1YPP0pYpBrDMHRLQ
frX4qpn+F75waZB1tpH6Rt56YbQKe72gRf1m4kPKT2nxbPNFLjg+xQXnmr81CJW3jSh38HTIDiU9
Q5t23qgA1ti4n27X7NOuavsr6Y21t2EWlSM47TutsqOcBfkZryAhtg551Tn0eJymrPz3EPL8J69M
YZfEUr4lHZNKftOsgiyw3/zGl3rYy55EAG6RWKe8mwUyceRsxVJGqjmMN1uH/lKgSCHqf+X630ob
F5AheFcMGYMLIHc5+5b6aQOSE0yxYaQeD/dtFit2Nwe7ORI9fr1cauMBT9sYstdIzPMNgHExzpkg
CzdvW8TN7NNUIAbCcgHul/PZMYJtvuEt8XUX8qN85YrJQSh9LmgGdYGfdL8J4CBNA1kuel9N8C0a
f7EKQ9I0Sq9yCX5rISrdWUuvfoG8qwYBF2Z5NS3Bts1ECZwOiPW4xWzo1mv+sac9qpcJHE3kkEHc
FHqpBMWhh5Hzm0OueyJw+ZnYT5aIddzv2O7TSIpn1/PPoMbo+rDMUV2l4RlMrwThcGwC+5cxhbO3
yMU8u1gTgVCdPeGTlo3dLGRe2r9sSuLuHacce46WemOh1sh5uzcHrLB0FuzjXfYhDlzphg5/MPYz
MoB3e/eq7oumEucy/83Q5rg0RbSJGDjIpWyPhfqPy9Cp4djhcIRXS8eg1rlTTkv8Piyi/8GUZXgP
hMetr5vmK7d27aJQrsRd2zEURjq2h73MEwBliL0NG/6oTNq+JlorFl52z4Cyba1Hle6DazOmOZd5
JEnGcI57KBZhB28rJGmkTARXZg2SWvTVHvckGVgKkq0RJwbdvvhuXEFRlfENZew+ro5oFcTUoxnl
AHBdeVQ1r8G1YskZmF5nJl7t7LP5ACWkF+SAquMFq8VGbOKevLg03RiUhEvcYKmHqQQee0uVJYix
nI8ps12EfuX0uXRNgQWan5JRIbxTbx1I1Y9AHCR9PZo3LjKe0GT11yQvRUjtW/h22ITG0Mr8tA6b
W1c3EjuOQpCLd82suzLrwv0m4qb4tUfCKzF2n2EnmivZhgUX//Zy3dTKP2RN93CKntG0z/raMvkv
q8F+L7pftY9YzEM3xd4UlKlNCTnLxOXG8uu1xCHaKVOYnuM1Hpm460LMVebg50Hw6L5/N4CKSN2b
aMI46meUeyvvEXoxwP792Wbf1lGHax/VxMins7govXq2A+V0l2GSA+q8hg/Ob7FG3w+hj3BYaKKC
/49vGdpTbDpCytYfCGlR6zDRhVrd0I8kQdJhpO+iCnacHmHVJUg2KQ4F5WhFAjhPQQpRRND7ZnWK
wwVcsJ8tG3zI9pv3nKk62fnpPSEHSY4TEmwMyQQGu6f1ll8Kfb+5eBWJNMgelS5wZLtslOLlvAQ5
5qSqnFT6i3LtOkpYL+HOnp2Ib/btnF3nnhrGIwAgw2jVmRJEI/hHuVr0JgHEctYKdFZNO0FL1oKG
/RiCMwMNA2z4Ic2l1ArSTxX2MWp5NZ9udZUHFWBS5siZJhMAKZ/Zig3zdSM/XRrkoitSztsI3p6w
lcQZLEd879NUbZ6bzht/LyCBLKqtMe8zKcXNB01+FzUKQvOhcoj1tbb3cAaCWDowd1n8Ft8ffHEq
w4hv9i3p0nDqNFrwkEpEvJbuOsBLPIW8Ozyz1P92grpMSyE+Zgo6XwWfD4a0Z+7uhWwGYp9Zw9g6
bqtZqvydB9SE3eIExV8dKOWoI6OxE13ZOX71BnefasK39LaLrFjWYj6m1f2NGDvymDNax/5xUNFb
xktvQHTHcu1llr58UWE3PGnTheTxi6TOrkfgIe4+I8ohrjL40Qv/9GICx1QIK2ZdBtyMn0efCrhX
hBJX4NCHS7wg4jHohMOFXxjBNeDDTNuAUd+YFZ1Dwd36syYgxxX/mvxqTbMdC7CPHL4SYHba4fGE
SCgj1/h2nj5A7kiMElOkVNwFWm2yJU+5tIpGbz65RcR6cGAAXfYfFF1klNS5wlyvoYaG2n/BixFw
5/TEuWKpj6dSIxMEb6K/MwKkEINHE3E59RjH5uyBo00SJw4n1K2Ryrz3FZEd6rgWAABxFNglh5bZ
pQlF/AQIINRnh8ebcM2KjDAU2wd0ZgdadPCZYiruX8qivjkK8APQUo5H0xWRdGRHO6GnJyIglD3w
ueduexdqvBzygFaUTF3VCroyxcOdrTs8wXKN2j9iA1BmKePrwcRXbBDfX63z3/yDxs/vmC8Bjytp
np5LETt83EAOl4K7P8M3qsiQGmzmUTo7usnDpPouNbpzTlDd7jX26mUI+3qzUPAlRuZpGlCb3JXT
6T1HZY1vaNSxZ37BjiaHmSw+hWMDeeNrOyT174VsYvX3u4SX5juQMrsnUZ95FBAwnU6Vq/LMomcC
F6sp4ADCA4mSKWlV1xbDyoY8PY1jOWZLvnH042PcizO5foPB6wBMZs1Dg5NQsemopxAkS+ybYrJ8
kAN/j2xIrlQRbV9F+o97suKmmD8lCoggfzAzkD/jSQ1LUv+iVFfkZuqbieM34QHMS8JzP85rB08S
wv3mmLCGkHvsyLVRyKqoNBiPmnvvxrL/2EbGnsPXHcj0oBHo4fVspBwFinZcYwXUedSmoadlpZpp
R9ObilO/H54=
`protect end_protected
